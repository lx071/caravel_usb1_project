// This is the unpowered netlist.
module usb_top (app_clk,
    reg_ack,
    reg_cs,
    reg_wr,
    usb_clk,
    usb_in_dn,
    usb_in_dp,
    usb_intr_o,
    usb_out_dn,
    usb_out_dp,
    usb_out_tx_oen,
    usb_rstn,
    wbd_clk_int,
    wbd_clk_usb,
    cfg_cska_usb,
    reg_addr,
    reg_be,
    reg_rdata,
    reg_wdata);
 input app_clk;
 output reg_ack;
 input reg_cs;
 input reg_wr;
 input usb_clk;
 input usb_in_dn;
 input usb_in_dp;
 output usb_intr_o;
 output usb_out_dn;
 output usb_out_dp;
 output usb_out_tx_oen;
 input usb_rstn;
 input wbd_clk_int;
 output wbd_clk_usb;
 input [3:0] cfg_cska_usb;
 input [8:0] reg_addr;
 input [3:0] reg_be;
 output [31:0] reg_rdata;
 input [31:0] reg_wdata;

 wire clknet_0_app_clk;
 wire \clknet_0_u_usb_host.u_async_wb.u_cmd_if._033_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_cmd_if._034_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_cmd_if._035_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_cmd_if._036_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_cmd_if._037_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_cmd_if._038_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_cmd_if._039_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_cmd_if._040_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_resp_if._014_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_resp_if._015_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_resp_if._016_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_resp_if._017_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_resp_if._018_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_resp_if._019_ ;
 wire \clknet_0_u_usb_host.u_core._171_ ;
 wire \clknet_0_u_usb_host.u_core._172_ ;
 wire \clknet_0_u_usb_host.u_core._178_ ;
 wire \clknet_0_u_usb_host.u_core._183_ ;
 wire \clknet_0_u_usb_host.u_core._184_ ;
 wire \clknet_0_u_usb_host.u_core._185_ ;
 wire \clknet_0_u_usb_host.u_core._193_ ;
 wire \clknet_0_u_usb_host.u_core._200_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0717_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0718_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0719_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0720_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0721_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0722_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0723_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0724_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0725_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0726_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0727_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0728_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0729_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0730_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0731_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0732_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0733_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0734_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0735_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0736_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0737_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0738_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0739_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0740_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0741_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0742_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0743_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0744_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0745_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0746_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0747_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0748_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0749_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0750_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0751_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0752_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0753_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0754_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0755_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0756_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0757_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0758_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0759_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0760_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0761_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0762_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0763_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0764_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0765_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0766_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0767_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0768_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0769_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0770_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0771_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0772_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0773_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0774_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0775_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0776_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0777_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0778_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0779_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0780_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0781_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0782_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0783_ ;
 wire \clknet_0_u_usb_host.u_core.u_sie._00_ ;
 wire \clknet_0_u_usb_host.u_phy._175_ ;
 wire \clknet_0_u_usb_host.u_phy._178_ ;
 wire \clknet_0_u_usb_host.u_phy._180_ ;
 wire \clknet_0_u_usb_host.u_phy._187_ ;
 wire \clknet_0_u_usb_host.u_phy._188_ ;
 wire clknet_0_usb_clk;
 wire clknet_1_0__leaf_app_clk;
 wire \clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._033_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._034_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._035_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._036_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._014_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._015_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._016_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._017_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core._171_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core._172_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core._178_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core._183_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core._184_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core._185_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core._193_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0717_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0718_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0719_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0720_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_phy._175_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_phy._178_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_phy._180_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_phy._187_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_phy._188_ ;
 wire clknet_1_1__leaf_app_clk;
 wire \clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._033_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._034_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._035_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._036_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._014_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._015_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._016_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._017_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core._171_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core._172_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core._178_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core._183_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core._184_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core._185_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core._193_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0717_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0718_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0719_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0720_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_phy._175_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_phy._178_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_phy._180_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_phy._187_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_phy._188_ ;
 wire \clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ;
 wire \clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ;
 wire \clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ;
 wire \clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ;
 wire \clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ;
 wire \clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ;
 wire \clknet_2_0__leaf_u_usb_host.u_core._200_ ;
 wire \clknet_2_0__leaf_u_usb_host.u_core.u_sie._00_ ;
 wire \clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ;
 wire \clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ;
 wire \clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ;
 wire \clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ;
 wire \clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ;
 wire \clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ;
 wire \clknet_2_1__leaf_u_usb_host.u_core._200_ ;
 wire \clknet_2_1__leaf_u_usb_host.u_core.u_sie._00_ ;
 wire \clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ;
 wire \clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ;
 wire \clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ;
 wire \clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ;
 wire \clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ;
 wire \clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ;
 wire \clknet_2_2__leaf_u_usb_host.u_core._200_ ;
 wire \clknet_2_2__leaf_u_usb_host.u_core.u_sie._00_ ;
 wire \clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ;
 wire \clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ;
 wire \clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ;
 wire \clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ;
 wire \clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ;
 wire \clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ;
 wire \clknet_2_3__leaf_u_usb_host.u_core._200_ ;
 wire \clknet_2_3__leaf_u_usb_host.u_core.u_sie._00_ ;
 wire clknet_4_0_0_usb_clk;
 wire clknet_4_10_0_usb_clk;
 wire clknet_4_11_0_usb_clk;
 wire clknet_4_12_0_usb_clk;
 wire clknet_4_13_0_usb_clk;
 wire clknet_4_14_0_usb_clk;
 wire clknet_4_15_0_usb_clk;
 wire clknet_4_1_0_usb_clk;
 wire clknet_4_2_0_usb_clk;
 wire clknet_4_3_0_usb_clk;
 wire clknet_4_4_0_usb_clk;
 wire clknet_4_5_0_usb_clk;
 wire clknet_4_6_0_usb_clk;
 wire clknet_4_7_0_usb_clk;
 wire clknet_4_8_0_usb_clk;
 wire clknet_4_9_0_usb_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \u_skew_usb.clk_d1 ;
 wire \u_skew_usb.clk_d10 ;
 wire \u_skew_usb.clk_d11 ;
 wire \u_skew_usb.clk_d12 ;
 wire \u_skew_usb.clk_d13 ;
 wire \u_skew_usb.clk_d14 ;
 wire \u_skew_usb.clk_d15 ;
 wire \u_skew_usb.clk_d2 ;
 wire \u_skew_usb.clk_d3 ;
 wire \u_skew_usb.clk_d4 ;
 wire \u_skew_usb.clk_d5 ;
 wire \u_skew_usb.clk_d6 ;
 wire \u_skew_usb.clk_d7 ;
 wire \u_skew_usb.clk_d8 ;
 wire \u_skew_usb.clk_d9 ;
 wire \u_skew_usb.clk_inbuf ;
 wire \u_skew_usb.clkbuf_1.X1 ;
 wire \u_skew_usb.clkbuf_1.X2 ;
 wire \u_skew_usb.clkbuf_1.X3 ;
 wire \u_skew_usb.clkbuf_10.X1 ;
 wire \u_skew_usb.clkbuf_10.X2 ;
 wire \u_skew_usb.clkbuf_10.X3 ;
 wire \u_skew_usb.clkbuf_11.X1 ;
 wire \u_skew_usb.clkbuf_11.X2 ;
 wire \u_skew_usb.clkbuf_11.X3 ;
 wire \u_skew_usb.clkbuf_12.X1 ;
 wire \u_skew_usb.clkbuf_12.X2 ;
 wire \u_skew_usb.clkbuf_12.X3 ;
 wire \u_skew_usb.clkbuf_13.X1 ;
 wire \u_skew_usb.clkbuf_13.X2 ;
 wire \u_skew_usb.clkbuf_13.X3 ;
 wire \u_skew_usb.clkbuf_14.X1 ;
 wire \u_skew_usb.clkbuf_14.X2 ;
 wire \u_skew_usb.clkbuf_14.X3 ;
 wire \u_skew_usb.clkbuf_15.X1 ;
 wire \u_skew_usb.clkbuf_15.X2 ;
 wire \u_skew_usb.clkbuf_15.X3 ;
 wire \u_skew_usb.clkbuf_2.X1 ;
 wire \u_skew_usb.clkbuf_2.X2 ;
 wire \u_skew_usb.clkbuf_2.X3 ;
 wire \u_skew_usb.clkbuf_3.X1 ;
 wire \u_skew_usb.clkbuf_3.X2 ;
 wire \u_skew_usb.clkbuf_3.X3 ;
 wire \u_skew_usb.clkbuf_4.X1 ;
 wire \u_skew_usb.clkbuf_4.X2 ;
 wire \u_skew_usb.clkbuf_4.X3 ;
 wire \u_skew_usb.clkbuf_5.X1 ;
 wire \u_skew_usb.clkbuf_5.X2 ;
 wire \u_skew_usb.clkbuf_5.X3 ;
 wire \u_skew_usb.clkbuf_6.X1 ;
 wire \u_skew_usb.clkbuf_6.X2 ;
 wire \u_skew_usb.clkbuf_6.X3 ;
 wire \u_skew_usb.clkbuf_7.X1 ;
 wire \u_skew_usb.clkbuf_7.X2 ;
 wire \u_skew_usb.clkbuf_7.X3 ;
 wire \u_skew_usb.clkbuf_8.X1 ;
 wire \u_skew_usb.clkbuf_8.X2 ;
 wire \u_skew_usb.clkbuf_8.X3 ;
 wire \u_skew_usb.clkbuf_9.X1 ;
 wire \u_skew_usb.clkbuf_9.X2 ;
 wire \u_skew_usb.clkbuf_9.X3 ;
 wire \u_skew_usb.d00 ;
 wire \u_skew_usb.d01 ;
 wire \u_skew_usb.d02 ;
 wire \u_skew_usb.d03 ;
 wire \u_skew_usb.d04 ;
 wire \u_skew_usb.d05 ;
 wire \u_skew_usb.d06 ;
 wire \u_skew_usb.d07 ;
 wire \u_skew_usb.d10 ;
 wire \u_skew_usb.d11 ;
 wire \u_skew_usb.d12 ;
 wire \u_skew_usb.d13 ;
 wire \u_skew_usb.d20 ;
 wire \u_skew_usb.d21 ;
 wire \u_skew_usb.d30 ;
 wire \u_skew_usb.in0 ;
 wire \u_skew_usb.in1 ;
 wire \u_skew_usb.in10 ;
 wire \u_skew_usb.in11 ;
 wire \u_skew_usb.in12 ;
 wire \u_skew_usb.in13 ;
 wire \u_skew_usb.in14 ;
 wire \u_skew_usb.in15 ;
 wire \u_skew_usb.in2 ;
 wire \u_skew_usb.in3 ;
 wire \u_skew_usb.in4 ;
 wire \u_skew_usb.in5 ;
 wire \u_skew_usb.in6 ;
 wire \u_skew_usb.in7 ;
 wire \u_skew_usb.in8 ;
 wire \u_skew_usb.in9 ;
 wire \u_usb_host.reg_ack ;
 wire \u_usb_host.reg_addr[0] ;
 wire \u_usb_host.reg_addr[1] ;
 wire \u_usb_host.reg_addr[2] ;
 wire \u_usb_host.reg_addr[3] ;
 wire \u_usb_host.reg_addr[4] ;
 wire \u_usb_host.reg_addr[5] ;
 wire \u_usb_host.reg_cs ;
 wire \u_usb_host.reg_rdata[0] ;
 wire \u_usb_host.reg_rdata[10] ;
 wire \u_usb_host.reg_rdata[11] ;
 wire \u_usb_host.reg_rdata[12] ;
 wire \u_usb_host.reg_rdata[13] ;
 wire \u_usb_host.reg_rdata[14] ;
 wire \u_usb_host.reg_rdata[15] ;
 wire \u_usb_host.reg_rdata[16] ;
 wire \u_usb_host.reg_rdata[17] ;
 wire \u_usb_host.reg_rdata[18] ;
 wire \u_usb_host.reg_rdata[19] ;
 wire \u_usb_host.reg_rdata[1] ;
 wire \u_usb_host.reg_rdata[20] ;
 wire \u_usb_host.reg_rdata[21] ;
 wire \u_usb_host.reg_rdata[22] ;
 wire \u_usb_host.reg_rdata[23] ;
 wire \u_usb_host.reg_rdata[24] ;
 wire \u_usb_host.reg_rdata[25] ;
 wire \u_usb_host.reg_rdata[26] ;
 wire \u_usb_host.reg_rdata[27] ;
 wire \u_usb_host.reg_rdata[28] ;
 wire \u_usb_host.reg_rdata[29] ;
 wire \u_usb_host.reg_rdata[2] ;
 wire \u_usb_host.reg_rdata[30] ;
 wire \u_usb_host.reg_rdata[31] ;
 wire \u_usb_host.reg_rdata[3] ;
 wire \u_usb_host.reg_rdata[4] ;
 wire \u_usb_host.reg_rdata[5] ;
 wire \u_usb_host.reg_rdata[6] ;
 wire \u_usb_host.reg_rdata[7] ;
 wire \u_usb_host.reg_rdata[8] ;
 wire \u_usb_host.reg_rdata[9] ;
 wire \u_usb_host.reg_wdata[0] ;
 wire \u_usb_host.reg_wdata[10] ;
 wire \u_usb_host.reg_wdata[11] ;
 wire \u_usb_host.reg_wdata[12] ;
 wire \u_usb_host.reg_wdata[13] ;
 wire \u_usb_host.reg_wdata[14] ;
 wire \u_usb_host.reg_wdata[15] ;
 wire \u_usb_host.reg_wdata[16] ;
 wire \u_usb_host.reg_wdata[17] ;
 wire \u_usb_host.reg_wdata[18] ;
 wire \u_usb_host.reg_wdata[19] ;
 wire \u_usb_host.reg_wdata[1] ;
 wire \u_usb_host.reg_wdata[20] ;
 wire \u_usb_host.reg_wdata[21] ;
 wire \u_usb_host.reg_wdata[22] ;
 wire \u_usb_host.reg_wdata[23] ;
 wire \u_usb_host.reg_wdata[28] ;
 wire \u_usb_host.reg_wdata[29] ;
 wire \u_usb_host.reg_wdata[2] ;
 wire \u_usb_host.reg_wdata[30] ;
 wire \u_usb_host.reg_wdata[31] ;
 wire \u_usb_host.reg_wdata[3] ;
 wire \u_usb_host.reg_wdata[4] ;
 wire \u_usb_host.reg_wdata[5] ;
 wire \u_usb_host.reg_wdata[6] ;
 wire \u_usb_host.reg_wdata[7] ;
 wire \u_usb_host.reg_wdata[8] ;
 wire \u_usb_host.reg_wdata[9] ;
 wire \u_usb_host.reg_wr ;
 wire \u_usb_host.u_async_wb.PendingRd ;
 wire \u_usb_host.u_async_wb._00_ ;
 wire \u_usb_host.u_async_wb._01_ ;
 wire \u_usb_host.u_async_wb._02_ ;
 wire \u_usb_host.u_async_wb._03_ ;
 wire \u_usb_host.u_async_wb._04_ ;
 wire \u_usb_host.u_async_wb._05_ ;
 wire \u_usb_host.u_async_wb.m_cmd_wr_afull ;
 wire \u_usb_host.u_async_wb.m_cmd_wr_en ;
 wire \u_usb_host.u_async_wb.m_cmd_wr_full ;
 wire \u_usb_host.u_async_wb.m_resp_rd_empty ;
 wire \u_usb_host.u_async_wb.m_resp_rd_en ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[10] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[11] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[12] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[13] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[14] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[15] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[16] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[17] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[18] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[19] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[20] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[21] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[22] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[23] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[24] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[25] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[26] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[27] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[32] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[33] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[34] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[35] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[36] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[37] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[38] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[39] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[40] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[41] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[42] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[4] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[5] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[6] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[7] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[8] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[9] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_empty ;
 wire \u_usb_host.u_async_wb.s_resp_wr_en ;
 wire \u_usb_host.u_async_wb.s_resp_wr_full ;
 wire \u_usb_host.u_async_wb.u_cmd_if._000_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._001_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._002_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._003_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._004_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._005_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._006_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._007_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._008_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._009_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._010_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._011_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._012_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._013_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._014_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._015_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._016_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._017_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._018_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._019_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._020_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._021_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._022_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._023_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._024_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._025_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._026_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._027_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._028_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._029_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._031_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._032_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._033_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._034_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._035_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._036_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._037_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._038_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._039_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._040_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if.grey_rd_ptr[0] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.grey_rd_ptr[1] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.grey_rd_ptr[2] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.grey_wr_ptr[0] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.grey_wr_ptr[1] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.grey_wr_ptr[2] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][10] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][11] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][12] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][13] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][14] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][15] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][16] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][17] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][18] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][19] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][20] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][21] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][22] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][23] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][24] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][25] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][26] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][27] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][32] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][33] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][34] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][35] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][36] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][37] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][38] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][39] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][40] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][41] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][42] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][4] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][5] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][6] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][7] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][8] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][9] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][10] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][11] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][12] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][13] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][14] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][15] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][16] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][17] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][18] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][19] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][20] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][21] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][22] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][23] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][24] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][25] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][26] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][27] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][32] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][33] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][34] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][35] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][36] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][37] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][38] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][39] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][40] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][41] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][42] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][4] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][5] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][6] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][7] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][8] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][9] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][10] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][11] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][12] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][13] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][14] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][15] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][16] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][17] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][18] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][19] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][20] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][21] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][22] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][23] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][24] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][25] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][26] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][27] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][32] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][33] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][34] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][35] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][36] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][37] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][38] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][39] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][40] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][41] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][42] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][4] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][5] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][6] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][7] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][8] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][9] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][10] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][11] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][12] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][13] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][14] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][15] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][16] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][17] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][18] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][19] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][20] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][21] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][22] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][23] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][24] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][25] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][26] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][27] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][32] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][33] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][34] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][35] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][36] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][37] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][38] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][39] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][40] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][41] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][42] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][4] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][5] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][6] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][7] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][8] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][9] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.rd_ptr[0] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.rd_ptr[1] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.rd_ptr[2] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[0] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[1] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[2] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.rd_reset_n ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr[2] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_0[0] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_0[1] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_0[2] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_1[0] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_1[1] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr[2] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_0[0] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_0[1] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_0[2] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_1[0] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_1[1] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.wr_ptr[0] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.wr_ptr[1] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.wr_ptr[2] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[0] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[1] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[2] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.wr_reset_n ;
 wire \u_usb_host.u_async_wb.u_resp_if._000_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._001_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._002_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._003_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._004_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._005_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._006_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._007_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._008_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._009_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._010_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._011_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._012_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._013_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._014_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._015_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._016_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._017_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._018_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._019_ ;
 wire \u_usb_host.u_async_wb.u_resp_if.grey_rd_ptr[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.grey_rd_ptr[1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.grey_wr_ptr[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.grey_wr_ptr[1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][10] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][11] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][12] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][13] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][14] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][15] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][16] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][17] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][18] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][19] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][20] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][21] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][22] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][23] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][24] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][25] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][26] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][27] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][28] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][29] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][2] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][30] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][31] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][3] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][4] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][5] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][6] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][7] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][8] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][9] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][10] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][11] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][12] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][13] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][14] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][15] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][16] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][17] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][18] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][19] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][20] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][21] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][22] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][23] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][24] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][25] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][26] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][27] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][28] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][29] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][2] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][30] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][31] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][3] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][4] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][5] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][6] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][7] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][8] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][9] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[10] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[11] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[12] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[13] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[14] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[15] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[16] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[17] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[18] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[19] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[20] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[21] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[22] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[23] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[24] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[25] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[26] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[27] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[28] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[29] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[2] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[30] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[31] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[3] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[4] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[5] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[6] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[7] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[8] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[9] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_ptr[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_ptr[1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_ptr_inc[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_ptr_inc[1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_0[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_0[1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_1[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_1[1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_0[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_0[1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_1[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_1[1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.wr_ptr[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.wr_ptr[1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.wr_ptr_inc[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.wr_ptr_inc[1] ;
 wire \u_usb_host.u_async_wb.wbm_cyc_i ;
 wire \u_usb_host.u_async_wb.wbs_ack_f ;
 wire \u_usb_host.u_async_wb.wbs_cyc_o ;
 wire \u_usb_host.u_core._000_ ;
 wire \u_usb_host.u_core._001_ ;
 wire \u_usb_host.u_core._002_ ;
 wire \u_usb_host.u_core._003_ ;
 wire \u_usb_host.u_core._004_ ;
 wire \u_usb_host.u_core._005_ ;
 wire \u_usb_host.u_core._006_ ;
 wire \u_usb_host.u_core._007_ ;
 wire \u_usb_host.u_core._008_ ;
 wire \u_usb_host.u_core._009_ ;
 wire \u_usb_host.u_core._010_ ;
 wire \u_usb_host.u_core._011_ ;
 wire \u_usb_host.u_core._012_ ;
 wire \u_usb_host.u_core._013_ ;
 wire \u_usb_host.u_core._014_ ;
 wire \u_usb_host.u_core._015_ ;
 wire \u_usb_host.u_core._016_ ;
 wire \u_usb_host.u_core._017_ ;
 wire \u_usb_host.u_core._018_ ;
 wire \u_usb_host.u_core._019_ ;
 wire \u_usb_host.u_core._020_ ;
 wire \u_usb_host.u_core._021_ ;
 wire \u_usb_host.u_core._022_ ;
 wire \u_usb_host.u_core._023_ ;
 wire \u_usb_host.u_core._025_ ;
 wire \u_usb_host.u_core._026_ ;
 wire \u_usb_host.u_core._027_ ;
 wire \u_usb_host.u_core._028_ ;
 wire \u_usb_host.u_core._029_ ;
 wire \u_usb_host.u_core._030_ ;
 wire \u_usb_host.u_core._032_ ;
 wire \u_usb_host.u_core._033_ ;
 wire \u_usb_host.u_core._034_ ;
 wire \u_usb_host.u_core._035_ ;
 wire \u_usb_host.u_core._036_ ;
 wire \u_usb_host.u_core._037_ ;
 wire \u_usb_host.u_core._038_ ;
 wire \u_usb_host.u_core._040_ ;
 wire \u_usb_host.u_core._041_ ;
 wire \u_usb_host.u_core._042_ ;
 wire \u_usb_host.u_core._043_ ;
 wire \u_usb_host.u_core._044_ ;
 wire \u_usb_host.u_core._045_ ;
 wire \u_usb_host.u_core._046_ ;
 wire \u_usb_host.u_core._047_ ;
 wire \u_usb_host.u_core._061_ ;
 wire \u_usb_host.u_core._062_ ;
 wire \u_usb_host.u_core._063_ ;
 wire \u_usb_host.u_core._064_ ;
 wire \u_usb_host.u_core._065_ ;
 wire \u_usb_host.u_core._066_ ;
 wire \u_usb_host.u_core._067_ ;
 wire \u_usb_host.u_core._068_ ;
 wire \u_usb_host.u_core._069_ ;
 wire \u_usb_host.u_core._070_ ;
 wire \u_usb_host.u_core._071_ ;
 wire \u_usb_host.u_core._072_ ;
 wire \u_usb_host.u_core._073_ ;
 wire \u_usb_host.u_core._074_ ;
 wire \u_usb_host.u_core._075_ ;
 wire \u_usb_host.u_core._076_ ;
 wire \u_usb_host.u_core._077_ ;
 wire \u_usb_host.u_core._078_ ;
 wire \u_usb_host.u_core._079_ ;
 wire \u_usb_host.u_core._080_ ;
 wire \u_usb_host.u_core._081_ ;
 wire \u_usb_host.u_core._082_ ;
 wire \u_usb_host.u_core._083_ ;
 wire \u_usb_host.u_core._084_ ;
 wire \u_usb_host.u_core._085_ ;
 wire \u_usb_host.u_core._086_ ;
 wire \u_usb_host.u_core._087_ ;
 wire \u_usb_host.u_core._088_ ;
 wire \u_usb_host.u_core._089_ ;
 wire \u_usb_host.u_core._090_ ;
 wire \u_usb_host.u_core._091_ ;
 wire \u_usb_host.u_core._092_ ;
 wire \u_usb_host.u_core._093_ ;
 wire \u_usb_host.u_core._094_ ;
 wire \u_usb_host.u_core._095_ ;
 wire \u_usb_host.u_core._096_ ;
 wire \u_usb_host.u_core._097_ ;
 wire \u_usb_host.u_core._098_ ;
 wire \u_usb_host.u_core._099_ ;
 wire \u_usb_host.u_core._100_ ;
 wire \u_usb_host.u_core._101_ ;
 wire \u_usb_host.u_core._102_ ;
 wire \u_usb_host.u_core._103_ ;
 wire \u_usb_host.u_core._104_ ;
 wire \u_usb_host.u_core._105_ ;
 wire \u_usb_host.u_core._106_ ;
 wire \u_usb_host.u_core._107_ ;
 wire \u_usb_host.u_core._108_ ;
 wire \u_usb_host.u_core._109_ ;
 wire \u_usb_host.u_core._110_ ;
 wire \u_usb_host.u_core._111_ ;
 wire \u_usb_host.u_core._112_ ;
 wire \u_usb_host.u_core._113_ ;
 wire \u_usb_host.u_core._114_ ;
 wire \u_usb_host.u_core._115_ ;
 wire \u_usb_host.u_core._116_ ;
 wire \u_usb_host.u_core._117_ ;
 wire \u_usb_host.u_core._118_ ;
 wire \u_usb_host.u_core._119_ ;
 wire \u_usb_host.u_core._120_ ;
 wire \u_usb_host.u_core._121_ ;
 wire \u_usb_host.u_core._122_ ;
 wire \u_usb_host.u_core._123_ ;
 wire \u_usb_host.u_core._124_ ;
 wire \u_usb_host.u_core._125_ ;
 wire \u_usb_host.u_core._126_ ;
 wire \u_usb_host.u_core._127_ ;
 wire \u_usb_host.u_core._128_ ;
 wire \u_usb_host.u_core._129_ ;
 wire \u_usb_host.u_core._130_ ;
 wire \u_usb_host.u_core._131_ ;
 wire \u_usb_host.u_core._132_ ;
 wire \u_usb_host.u_core._133_ ;
 wire \u_usb_host.u_core._134_ ;
 wire \u_usb_host.u_core._135_ ;
 wire \u_usb_host.u_core._136_ ;
 wire \u_usb_host.u_core._137_ ;
 wire \u_usb_host.u_core._138_ ;
 wire \u_usb_host.u_core._139_ ;
 wire \u_usb_host.u_core._140_ ;
 wire \u_usb_host.u_core._141_ ;
 wire \u_usb_host.u_core._142_ ;
 wire \u_usb_host.u_core._143_ ;
 wire \u_usb_host.u_core._144_ ;
 wire \u_usb_host.u_core._145_ ;
 wire \u_usb_host.u_core._146_ ;
 wire \u_usb_host.u_core._147_ ;
 wire \u_usb_host.u_core._148_ ;
 wire \u_usb_host.u_core._149_ ;
 wire \u_usb_host.u_core._150_ ;
 wire \u_usb_host.u_core._151_ ;
 wire \u_usb_host.u_core._152_ ;
 wire \u_usb_host.u_core._153_ ;
 wire \u_usb_host.u_core._154_ ;
 wire \u_usb_host.u_core._155_ ;
 wire \u_usb_host.u_core._156_ ;
 wire \u_usb_host.u_core._157_ ;
 wire \u_usb_host.u_core._158_ ;
 wire \u_usb_host.u_core._171_ ;
 wire \u_usb_host.u_core._172_ ;
 wire \u_usb_host.u_core._173_ ;
 wire \u_usb_host.u_core._174_ ;
 wire \u_usb_host.u_core._175_ ;
 wire \u_usb_host.u_core._176_ ;
 wire \u_usb_host.u_core._177_ ;
 wire \u_usb_host.u_core._178_ ;
 wire \u_usb_host.u_core._179_ ;
 wire \u_usb_host.u_core._180_ ;
 wire \u_usb_host.u_core._181_ ;
 wire \u_usb_host.u_core._182_ ;
 wire \u_usb_host.u_core._183_ ;
 wire \u_usb_host.u_core._184_ ;
 wire \u_usb_host.u_core._185_ ;
 wire \u_usb_host.u_core._187_ ;
 wire \u_usb_host.u_core._188_ ;
 wire \u_usb_host.u_core._193_ ;
 wire \u_usb_host.u_core._194_ ;
 wire \u_usb_host.u_core._195_ ;
 wire \u_usb_host.u_core._196_ ;
 wire \u_usb_host.u_core._197_ ;
 wire \u_usb_host.u_core._198_ ;
 wire \u_usb_host.u_core._199_ ;
 wire \u_usb_host.u_core._200_ ;
 wire \u_usb_host.u_core._201_ ;
 wire \u_usb_host.u_core._202_ ;
 wire \u_usb_host.u_core.cfg_wr ;
 wire \u_usb_host.u_core.device_det_q ;
 wire \u_usb_host.u_core.err_cond_q ;
 wire \u_usb_host.u_core.fifo_flush_q ;
 wire \u_usb_host.u_core.fifo_rx_data_w[0] ;
 wire \u_usb_host.u_core.fifo_rx_data_w[1] ;
 wire \u_usb_host.u_core.fifo_rx_data_w[2] ;
 wire \u_usb_host.u_core.fifo_rx_data_w[3] ;
 wire \u_usb_host.u_core.fifo_rx_data_w[4] ;
 wire \u_usb_host.u_core.fifo_rx_data_w[5] ;
 wire \u_usb_host.u_core.fifo_rx_data_w[6] ;
 wire \u_usb_host.u_core.fifo_rx_data_w[7] ;
 wire \u_usb_host.u_core.intr_done_q ;
 wire \u_usb_host.u_core.intr_err_q ;
 wire \u_usb_host.u_core.intr_sof_q ;
 wire \u_usb_host.u_core.reg_rdata_r[0] ;
 wire \u_usb_host.u_core.reg_rdata_r[10] ;
 wire \u_usb_host.u_core.reg_rdata_r[11] ;
 wire \u_usb_host.u_core.reg_rdata_r[12] ;
 wire \u_usb_host.u_core.reg_rdata_r[13] ;
 wire \u_usb_host.u_core.reg_rdata_r[14] ;
 wire \u_usb_host.u_core.reg_rdata_r[15] ;
 wire \u_usb_host.u_core.reg_rdata_r[16] ;
 wire \u_usb_host.u_core.reg_rdata_r[17] ;
 wire \u_usb_host.u_core.reg_rdata_r[18] ;
 wire \u_usb_host.u_core.reg_rdata_r[19] ;
 wire \u_usb_host.u_core.reg_rdata_r[1] ;
 wire \u_usb_host.u_core.reg_rdata_r[20] ;
 wire \u_usb_host.u_core.reg_rdata_r[21] ;
 wire \u_usb_host.u_core.reg_rdata_r[22] ;
 wire \u_usb_host.u_core.reg_rdata_r[23] ;
 wire \u_usb_host.u_core.reg_rdata_r[24] ;
 wire \u_usb_host.u_core.reg_rdata_r[25] ;
 wire \u_usb_host.u_core.reg_rdata_r[26] ;
 wire \u_usb_host.u_core.reg_rdata_r[27] ;
 wire \u_usb_host.u_core.reg_rdata_r[28] ;
 wire \u_usb_host.u_core.reg_rdata_r[29] ;
 wire \u_usb_host.u_core.reg_rdata_r[2] ;
 wire \u_usb_host.u_core.reg_rdata_r[30] ;
 wire \u_usb_host.u_core.reg_rdata_r[31] ;
 wire \u_usb_host.u_core.reg_rdata_r[3] ;
 wire \u_usb_host.u_core.reg_rdata_r[4] ;
 wire \u_usb_host.u_core.reg_rdata_r[5] ;
 wire \u_usb_host.u_core.reg_rdata_r[6] ;
 wire \u_usb_host.u_core.reg_rdata_r[7] ;
 wire \u_usb_host.u_core.reg_rdata_r[8] ;
 wire \u_usb_host.u_core.reg_rdata_r[9] ;
 wire \u_usb_host.u_core.send_sof_w ;
 wire \u_usb_host.u_core.sof_irq_q ;
 wire \u_usb_host.u_core.sof_time_q[0] ;
 wire \u_usb_host.u_core.sof_time_q[10] ;
 wire \u_usb_host.u_core.sof_time_q[11] ;
 wire \u_usb_host.u_core.sof_time_q[12] ;
 wire \u_usb_host.u_core.sof_time_q[13] ;
 wire \u_usb_host.u_core.sof_time_q[14] ;
 wire \u_usb_host.u_core.sof_time_q[15] ;
 wire \u_usb_host.u_core.sof_time_q[1] ;
 wire \u_usb_host.u_core.sof_time_q[2] ;
 wire \u_usb_host.u_core.sof_time_q[3] ;
 wire \u_usb_host.u_core.sof_time_q[4] ;
 wire \u_usb_host.u_core.sof_time_q[5] ;
 wire \u_usb_host.u_core.sof_time_q[6] ;
 wire \u_usb_host.u_core.sof_time_q[7] ;
 wire \u_usb_host.u_core.sof_time_q[8] ;
 wire \u_usb_host.u_core.sof_time_q[9] ;
 wire \u_usb_host.u_core.transfer_start_q ;
 wire \u_usb_host.u_core.u_fifo_rx._0000_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0001_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0002_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0003_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0004_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0005_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0006_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0007_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0008_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0009_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0010_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0011_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0012_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0013_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0014_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0015_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0016_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0017_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0018_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0019_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0020_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0021_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0022_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0023_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0024_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0025_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0026_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0027_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0028_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0029_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0030_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0031_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0032_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0033_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0034_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0035_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0036_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0037_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0038_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0039_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0040_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0041_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0042_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0043_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0044_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0045_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0046_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0047_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0048_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0049_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0050_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0051_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0052_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0053_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0054_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0055_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0056_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0057_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0058_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0059_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0060_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0061_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0062_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0063_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0064_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0065_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0066_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0067_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0068_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0069_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0070_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0071_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0072_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0073_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0074_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0075_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0076_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0077_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0078_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0079_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0080_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0081_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0082_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0083_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0084_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0085_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0086_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0087_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0088_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0089_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0090_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0091_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0092_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0093_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0094_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0095_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0096_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0097_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0098_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0099_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0100_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0101_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0102_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0103_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0104_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0105_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0106_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0107_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0108_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0109_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0110_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0111_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0112_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0113_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0114_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0115_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0116_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0117_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0118_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0119_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0120_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0121_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0122_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0123_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0124_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0125_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0126_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0127_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0128_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0129_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0130_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0131_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0132_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0133_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0134_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0135_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0136_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0137_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0138_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0139_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0140_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0141_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0142_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0143_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0144_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0145_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0146_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0147_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0148_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0149_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0150_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0151_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0152_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0153_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0154_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0155_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0156_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0157_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0158_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0159_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0160_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0161_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0162_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0163_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0164_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0165_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0166_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0167_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0168_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0169_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0170_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0171_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0172_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0173_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0174_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0175_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0176_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0177_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0178_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0179_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0180_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0181_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0182_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0183_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0184_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0185_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0186_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0187_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0188_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0189_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0190_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0191_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0192_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0193_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0194_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0195_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0196_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0197_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0198_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0199_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0200_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0201_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0202_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0203_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0204_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0205_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0206_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0207_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0208_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0209_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0210_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0211_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0212_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0213_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0214_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0215_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0216_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0217_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0218_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0219_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0220_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0221_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0222_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0223_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0224_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0225_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0226_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0227_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0228_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0229_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0230_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0231_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0232_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0233_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0234_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0235_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0236_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0237_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0238_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0239_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0240_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0241_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0242_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0243_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0244_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0245_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0246_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0247_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0248_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0249_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0250_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0251_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0252_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0253_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0254_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0255_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0256_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0257_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0258_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0259_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0260_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0261_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0262_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0263_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0264_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0265_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0266_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0267_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0268_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0269_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0270_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0271_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0272_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0273_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0274_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0275_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0276_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0277_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0278_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0279_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0280_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0281_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0282_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0283_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0284_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0285_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0286_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0287_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0288_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0289_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0290_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0291_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0292_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0293_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0294_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0295_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0296_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0297_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0298_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0299_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0300_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0301_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0302_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0303_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0304_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0305_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0306_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0307_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0308_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0309_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0310_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0311_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0312_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0313_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0314_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0315_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0316_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0317_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0318_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0319_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0320_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0321_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0322_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0323_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0324_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0325_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0326_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0327_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0328_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0329_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0330_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0331_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0332_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0333_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0334_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0335_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0336_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0337_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0338_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0339_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0340_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0341_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0342_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0343_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0344_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0345_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0346_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0347_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0348_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0349_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0350_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0351_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0352_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0353_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0354_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0355_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0356_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0357_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0358_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0359_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0360_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0361_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0362_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0363_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0364_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0365_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0366_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0367_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0368_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0369_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0370_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0371_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0372_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0373_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0374_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0375_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0376_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0377_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0378_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0379_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0380_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0381_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0382_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0383_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0384_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0385_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0386_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0387_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0388_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0389_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0390_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0391_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0392_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0393_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0394_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0395_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0396_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0397_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0398_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0399_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0400_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0401_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0402_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0403_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0404_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0405_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0406_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0407_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0408_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0409_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0410_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0411_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0412_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0413_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0414_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0415_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0416_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0417_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0418_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0419_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0420_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0421_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0422_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0423_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0424_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0425_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0426_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0427_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0428_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0429_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0430_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0431_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0432_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0433_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0434_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0435_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0436_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0437_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0438_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0439_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0440_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0441_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0442_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0443_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0444_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0445_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0446_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0447_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0448_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0449_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0450_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0451_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0452_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0453_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0454_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0455_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0456_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0457_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0458_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0459_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0460_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0461_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0462_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0463_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0464_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0465_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0466_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0467_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0468_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0469_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0470_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0471_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0472_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0473_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0474_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0475_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0476_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0477_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0478_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0479_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0480_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0481_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0482_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0483_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0484_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0485_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0486_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0487_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0488_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0489_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0490_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0491_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0492_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0493_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0494_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0495_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0496_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0497_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0498_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0499_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0500_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0501_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0502_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0503_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0504_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0505_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0506_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0507_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0508_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0509_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0510_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0511_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0512_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0513_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0514_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0515_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0516_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0517_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0518_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0519_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0520_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0521_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0522_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0523_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0524_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0525_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0526_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0527_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0528_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0529_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0530_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0531_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0532_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0533_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0534_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0535_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0536_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0537_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0538_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0539_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0540_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0541_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0542_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0543_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0544_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0545_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0546_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0547_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0548_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0549_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0550_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0551_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0552_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0553_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0554_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0555_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0556_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0557_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0558_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0559_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0560_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0561_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0562_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0563_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0564_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0565_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0566_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0567_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0568_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0569_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0570_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0571_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0572_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0573_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0574_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0575_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0576_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0577_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0578_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0579_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0580_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0581_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0582_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0583_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0584_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0585_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0586_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0587_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0588_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0589_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0590_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0591_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0592_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0593_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0594_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0595_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0596_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0597_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0598_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0599_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0600_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0601_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0602_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0603_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0604_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0605_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0606_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0607_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0608_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0609_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0610_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0611_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0612_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0613_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0614_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0615_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0616_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0617_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0618_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0619_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0620_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0621_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0622_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0623_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0624_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0625_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0626_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0627_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0628_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0629_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0630_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0631_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0632_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0633_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0634_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0635_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0636_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0637_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0638_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0639_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0640_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0641_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0642_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0643_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0644_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0645_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0646_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0647_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0648_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0649_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0650_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0651_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0652_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0653_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0654_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0655_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0656_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0657_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0658_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0659_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0660_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0661_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0662_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0663_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0664_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0665_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0666_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0667_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0668_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0669_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0670_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0671_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0672_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0673_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0674_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0675_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0676_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0677_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0678_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0679_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0680_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0681_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0682_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0683_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0684_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0685_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0686_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0687_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0688_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0689_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0690_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0691_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0692_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0693_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0694_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0695_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0696_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0697_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0698_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0699_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0700_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0701_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0702_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0703_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0704_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0705_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0706_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0707_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0708_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0709_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0710_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0711_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0712_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0713_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0714_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0715_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0716_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0717_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0718_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0719_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0720_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0721_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0722_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0723_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0724_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0725_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0726_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0727_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0728_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0729_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0730_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0731_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0732_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0733_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0734_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0735_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0736_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0737_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0738_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0739_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0740_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0741_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0742_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0743_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0744_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0745_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0746_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0747_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0748_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0749_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0750_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0751_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0752_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0753_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0754_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0755_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0756_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0757_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0758_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0759_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0760_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0761_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0762_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0763_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0764_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0765_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0766_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0767_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0768_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0769_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0770_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0771_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0772_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0773_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0774_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0775_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0776_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0777_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0778_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0779_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0780_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0781_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0782_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0783_ ;
 wire \u_usb_host.u_core.u_fifo_rx.count[0] ;
 wire \u_usb_host.u_core.u_fifo_rx.count[1] ;
 wire \u_usb_host.u_core.u_fifo_rx.count[2] ;
 wire \u_usb_host.u_core.u_fifo_rx.count[3] ;
 wire \u_usb_host.u_core.u_fifo_rx.count[4] ;
 wire \u_usb_host.u_core.u_fifo_rx.count[5] ;
 wire \u_usb_host.u_core.u_fifo_rx.count[6] ;
 wire \u_usb_host.u_core.u_fifo_rx.data_o[0] ;
 wire \u_usb_host.u_core.u_fifo_rx.data_o[1] ;
 wire \u_usb_host.u_core.u_fifo_rx.data_o[2] ;
 wire \u_usb_host.u_core.u_fifo_rx.data_o[3] ;
 wire \u_usb_host.u_core.u_fifo_rx.data_o[4] ;
 wire \u_usb_host.u_core.u_fifo_rx.data_o[5] ;
 wire \u_usb_host.u_core.u_fifo_rx.data_o[6] ;
 wire \u_usb_host.u_core.u_fifo_rx.data_o[7] ;
 wire \u_usb_host.u_core.u_fifo_rx.pop_i ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[0][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[0][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[0][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[0][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[0][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[0][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[0][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[0][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[10][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[10][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[10][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[10][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[10][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[10][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[10][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[10][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[11][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[11][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[11][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[11][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[11][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[11][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[11][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[11][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[12][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[12][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[12][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[12][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[12][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[12][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[12][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[12][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[13][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[13][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[13][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[13][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[13][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[13][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[13][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[13][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[14][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[14][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[14][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[14][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[14][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[14][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[14][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[14][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[15][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[15][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[15][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[15][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[15][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[15][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[15][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[15][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[16][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[16][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[16][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[16][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[16][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[16][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[16][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[16][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[17][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[17][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[17][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[17][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[17][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[17][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[17][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[17][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[18][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[18][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[18][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[18][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[18][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[18][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[18][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[18][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[19][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[19][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[19][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[19][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[19][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[19][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[19][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[19][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[1][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[1][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[1][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[1][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[1][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[1][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[1][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[1][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[20][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[20][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[20][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[20][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[20][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[20][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[20][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[20][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[21][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[21][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[21][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[21][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[21][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[21][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[21][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[21][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[22][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[22][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[22][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[22][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[22][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[22][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[22][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[22][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[23][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[23][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[23][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[23][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[23][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[23][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[23][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[23][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[24][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[24][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[24][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[24][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[24][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[24][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[24][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[24][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[25][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[25][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[25][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[25][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[25][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[25][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[25][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[25][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[26][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[26][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[26][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[26][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[26][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[26][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[26][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[26][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[27][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[27][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[27][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[27][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[27][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[27][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[27][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[27][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[28][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[28][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[28][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[28][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[28][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[28][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[28][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[28][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[29][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[29][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[29][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[29][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[29][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[29][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[29][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[29][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[2][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[2][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[2][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[2][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[2][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[2][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[2][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[2][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[30][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[30][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[30][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[30][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[30][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[30][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[30][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[30][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[31][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[31][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[31][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[31][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[31][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[31][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[31][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[31][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[32][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[32][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[32][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[32][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[32][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[32][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[32][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[32][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[33][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[33][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[33][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[33][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[33][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[33][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[33][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[33][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[34][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[34][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[34][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[34][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[34][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[34][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[34][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[34][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[35][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[35][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[35][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[35][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[35][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[35][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[35][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[35][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[36][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[36][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[36][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[36][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[36][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[36][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[36][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[36][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[37][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[37][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[37][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[37][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[37][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[37][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[37][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[37][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[38][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[38][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[38][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[38][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[38][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[38][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[38][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[38][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[39][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[39][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[39][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[39][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[39][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[39][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[39][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[39][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[3][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[3][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[3][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[3][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[3][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[3][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[3][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[3][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[40][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[40][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[40][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[40][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[40][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[40][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[40][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[40][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[41][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[41][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[41][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[41][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[41][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[41][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[41][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[41][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[42][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[42][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[42][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[42][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[42][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[42][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[42][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[42][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[43][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[43][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[43][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[43][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[43][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[43][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[43][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[43][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[44][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[44][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[44][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[44][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[44][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[44][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[44][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[45][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[45][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[45][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[45][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[45][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[45][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[45][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[45][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[46][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[46][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[46][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[46][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[46][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[46][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[46][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[46][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[47][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[47][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[47][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[47][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[47][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[47][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[47][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[47][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[48][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[48][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[48][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[48][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[48][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[48][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[48][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[48][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[49][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[49][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[49][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[49][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[49][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[49][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[49][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[49][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[4][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[4][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[4][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[4][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[4][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[4][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[4][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[4][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[50][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[50][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[50][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[50][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[50][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[50][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[50][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[50][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[51][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[51][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[51][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[51][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[51][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[51][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[51][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[51][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[52][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[52][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[52][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[52][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[52][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[52][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[52][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[52][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[53][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[53][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[53][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[53][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[53][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[53][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[53][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[53][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[54][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[54][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[54][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[54][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[54][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[54][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[54][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[54][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[55][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[55][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[55][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[55][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[55][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[55][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[55][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[55][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[56][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[56][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[56][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[56][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[56][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[56][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[56][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[56][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[57][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[57][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[57][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[57][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[57][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[57][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[57][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[57][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[58][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[58][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[58][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[58][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[58][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[58][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[58][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[58][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[59][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[59][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[59][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[59][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[59][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[59][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[59][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[59][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[5][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[5][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[5][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[5][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[5][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[5][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[5][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[5][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[60][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[60][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[60][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[60][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[60][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[60][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[60][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[60][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[61][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[61][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[61][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[61][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[61][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[61][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[61][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[61][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[62][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[62][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[62][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[62][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[62][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[62][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[62][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[62][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[63][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[63][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[63][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[63][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[63][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[63][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[63][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[63][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[6][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[6][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[6][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[6][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[6][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[6][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[6][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[6][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[7][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[7][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[7][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[7][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[7][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[7][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[7][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[7][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[8][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[8][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[8][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[8][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[8][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[8][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[8][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[8][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[9][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[9][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[9][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[9][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[9][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[9][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[9][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[9][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.rd_ptr[0] ;
 wire \u_usb_host.u_core.u_fifo_rx.rd_ptr[1] ;
 wire \u_usb_host.u_core.u_fifo_rx.rd_ptr[2] ;
 wire \u_usb_host.u_core.u_fifo_rx.rd_ptr[3] ;
 wire \u_usb_host.u_core.u_fifo_rx.rd_ptr[4] ;
 wire \u_usb_host.u_core.u_fifo_rx.rd_ptr[5] ;
 wire \u_usb_host.u_core.u_fifo_rx.wr_ptr[0] ;
 wire \u_usb_host.u_core.u_fifo_rx.wr_ptr[1] ;
 wire \u_usb_host.u_core.u_fifo_rx.wr_ptr[2] ;
 wire \u_usb_host.u_core.u_fifo_rx.wr_ptr[3] ;
 wire \u_usb_host.u_core.u_fifo_rx.wr_ptr[4] ;
 wire \u_usb_host.u_core.u_fifo_rx.wr_ptr[5] ;
 wire \u_usb_host.u_core.u_sie._00_ ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[0] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[10] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[11] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[12] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[13] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[14] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[15] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[16] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[17] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[18] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[19] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[1] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[20] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[21] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[22] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[23] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[24] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[25] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[26] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[27] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[28] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[29] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[2] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[30] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[31] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[3] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[4] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[5] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[6] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[7] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[8] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[9] ;
 wire \u_usb_host.u_core.u_sie.data_idx_i ;
 wire \u_usb_host.u_core.u_sie.data_len_i[0] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[10] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[11] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[12] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[13] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[14] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[15] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[1] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[2] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[3] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[4] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[5] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[6] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[7] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[8] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[9] ;
 wire \u_usb_host.u_core.u_sie.shift_en_w ;
 wire \u_usb_host.u_core.u_sie.utmi_data_i[0] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_i[1] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_i[2] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_i[3] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_i[4] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_i[5] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_i[6] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_i[7] ;
 wire \u_usb_host.u_core.u_sie.utmi_linestate_i[0] ;
 wire \u_usb_host.u_core.u_sie.utmi_linestate_i[1] ;
 wire \u_usb_host.u_core.u_sie.utmi_rxactive_i ;
 wire \u_usb_host.u_core.u_sie.utmi_rxvalid_i ;
 wire \u_usb_host.u_core.usb_ctrl_enable_sof_out_w ;
 wire \u_usb_host.u_core.usb_ctrl_wr_q ;
 wire \u_usb_host.u_core.usb_err_q ;
 wire \u_usb_host.u_core.usb_irq_ack_device_detect_out_w ;
 wire \u_usb_host.u_core.usb_irq_ack_done_out_w ;
 wire \u_usb_host.u_core.usb_irq_ack_err_out_w ;
 wire \u_usb_host.u_core.usb_irq_ack_sof_out_w ;
 wire \u_usb_host.u_core.usb_irq_mask_device_detect_out_w ;
 wire \u_usb_host.u_core.usb_irq_mask_done_out_w ;
 wire \u_usb_host.u_core.usb_irq_mask_err_out_w ;
 wire \u_usb_host.u_core.usb_irq_mask_sof_out_w ;
 wire \u_usb_host.u_core.usb_rx_stat_start_pend_in_w ;
 wire \u_usb_host.u_core.usb_xfer_token_ack_out_w ;
 wire \u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[0] ;
 wire \u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[1] ;
 wire \u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[2] ;
 wire \u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[3] ;
 wire \u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[4] ;
 wire \u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[5] ;
 wire \u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[6] ;
 wire \u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[0] ;
 wire \u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[1] ;
 wire \u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[2] ;
 wire \u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[3] ;
 wire \u_usb_host.u_core.usb_xfer_token_in_out_w ;
 wire \u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[0] ;
 wire \u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[1] ;
 wire \u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[2] ;
 wire \u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[3] ;
 wire \u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[4] ;
 wire \u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[5] ;
 wire \u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[6] ;
 wire \u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[7] ;
 wire \u_usb_host.u_core.utmi_dmpulldown_o ;
 wire \u_usb_host.u_core.utmi_dppulldown_o ;
 wire \u_usb_host.u_core.utmi_op_mode_o[0] ;
 wire \u_usb_host.u_core.utmi_op_mode_o[1] ;
 wire \u_usb_host.u_core.utmi_rxerror_i ;
 wire \u_usb_host.u_core.utmi_termselect_o ;
 wire \u_usb_host.u_core.utmi_xcvrselect_o[0] ;
 wire \u_usb_host.u_core.utmi_xcvrselect_o[1] ;
 wire \u_usb_host.u_phy._000_ ;
 wire \u_usb_host.u_phy._001_ ;
 wire \u_usb_host.u_phy._002_ ;
 wire \u_usb_host.u_phy._003_ ;
 wire \u_usb_host.u_phy._004_ ;
 wire \u_usb_host.u_phy._005_ ;
 wire \u_usb_host.u_phy._006_ ;
 wire \u_usb_host.u_phy._007_ ;
 wire \u_usb_host.u_phy._008_ ;
 wire \u_usb_host.u_phy._009_ ;
 wire \u_usb_host.u_phy._010_ ;
 wire \u_usb_host.u_phy._011_ ;
 wire \u_usb_host.u_phy._012_ ;
 wire \u_usb_host.u_phy._021_ ;
 wire \u_usb_host.u_phy._023_ ;
 wire \u_usb_host.u_phy._024_ ;
 wire \u_usb_host.u_phy._025_ ;
 wire \u_usb_host.u_phy._026_ ;
 wire \u_usb_host.u_phy._027_ ;
 wire \u_usb_host.u_phy._028_ ;
 wire \u_usb_host.u_phy._029_ ;
 wire \u_usb_host.u_phy._030_ ;
 wire \u_usb_host.u_phy._031_ ;
 wire \u_usb_host.u_phy._032_ ;
 wire \u_usb_host.u_phy._033_ ;
 wire \u_usb_host.u_phy._034_ ;
 wire \u_usb_host.u_phy._035_ ;
 wire \u_usb_host.u_phy._036_ ;
 wire \u_usb_host.u_phy._037_ ;
 wire \u_usb_host.u_phy._038_ ;
 wire \u_usb_host.u_phy._039_ ;
 wire \u_usb_host.u_phy._040_ ;
 wire \u_usb_host.u_phy._041_ ;
 wire \u_usb_host.u_phy._042_ ;
 wire \u_usb_host.u_phy._043_ ;
 wire \u_usb_host.u_phy._044_ ;
 wire \u_usb_host.u_phy._045_ ;
 wire \u_usb_host.u_phy._046_ ;
 wire \u_usb_host.u_phy._047_ ;
 wire \u_usb_host.u_phy._048_ ;
 wire \u_usb_host.u_phy._049_ ;
 wire \u_usb_host.u_phy._050_ ;
 wire \u_usb_host.u_phy._051_ ;
 wire \u_usb_host.u_phy._052_ ;
 wire \u_usb_host.u_phy._053_ ;
 wire \u_usb_host.u_phy._054_ ;
 wire \u_usb_host.u_phy._055_ ;
 wire \u_usb_host.u_phy._056_ ;
 wire \u_usb_host.u_phy._057_ ;
 wire \u_usb_host.u_phy._058_ ;
 wire \u_usb_host.u_phy._059_ ;
 wire \u_usb_host.u_phy._060_ ;
 wire \u_usb_host.u_phy._061_ ;
 wire \u_usb_host.u_phy._062_ ;
 wire \u_usb_host.u_phy._063_ ;
 wire \u_usb_host.u_phy._064_ ;
 wire \u_usb_host.u_phy._065_ ;
 wire \u_usb_host.u_phy._066_ ;
 wire \u_usb_host.u_phy._067_ ;
 wire \u_usb_host.u_phy._068_ ;
 wire \u_usb_host.u_phy._069_ ;
 wire \u_usb_host.u_phy._070_ ;
 wire \u_usb_host.u_phy._071_ ;
 wire \u_usb_host.u_phy._072_ ;
 wire \u_usb_host.u_phy._073_ ;
 wire \u_usb_host.u_phy._074_ ;
 wire \u_usb_host.u_phy._075_ ;
 wire \u_usb_host.u_phy._076_ ;
 wire \u_usb_host.u_phy._077_ ;
 wire \u_usb_host.u_phy._078_ ;
 wire \u_usb_host.u_phy._079_ ;
 wire \u_usb_host.u_phy._080_ ;
 wire \u_usb_host.u_phy._081_ ;
 wire \u_usb_host.u_phy._082_ ;
 wire \u_usb_host.u_phy._083_ ;
 wire \u_usb_host.u_phy._084_ ;
 wire \u_usb_host.u_phy._085_ ;
 wire \u_usb_host.u_phy._086_ ;
 wire \u_usb_host.u_phy._087_ ;
 wire \u_usb_host.u_phy._088_ ;
 wire \u_usb_host.u_phy._089_ ;
 wire \u_usb_host.u_phy._090_ ;
 wire \u_usb_host.u_phy._091_ ;
 wire \u_usb_host.u_phy._092_ ;
 wire \u_usb_host.u_phy._093_ ;
 wire \u_usb_host.u_phy._094_ ;
 wire \u_usb_host.u_phy._095_ ;
 wire \u_usb_host.u_phy._096_ ;
 wire \u_usb_host.u_phy._097_ ;
 wire \u_usb_host.u_phy._098_ ;
 wire \u_usb_host.u_phy._099_ ;
 wire \u_usb_host.u_phy._100_ ;
 wire \u_usb_host.u_phy._101_ ;
 wire \u_usb_host.u_phy._102_ ;
 wire \u_usb_host.u_phy._103_ ;
 wire \u_usb_host.u_phy._104_ ;
 wire \u_usb_host.u_phy._107_ ;
 wire \u_usb_host.u_phy._108_ ;
 wire \u_usb_host.u_phy._116_ ;
 wire \u_usb_host.u_phy._117_ ;
 wire \u_usb_host.u_phy._118_ ;
 wire \u_usb_host.u_phy._119_ ;
 wire \u_usb_host.u_phy._120_ ;
 wire \u_usb_host.u_phy._121_ ;
 wire \u_usb_host.u_phy._122_ ;
 wire \u_usb_host.u_phy._123_ ;
 wire \u_usb_host.u_phy._124_ ;
 wire \u_usb_host.u_phy._125_ ;
 wire \u_usb_host.u_phy._126_ ;
 wire \u_usb_host.u_phy._127_ ;
 wire \u_usb_host.u_phy._128_ ;
 wire \u_usb_host.u_phy._129_ ;
 wire \u_usb_host.u_phy._130_ ;
 wire \u_usb_host.u_phy._131_ ;
 wire \u_usb_host.u_phy._132_ ;
 wire \u_usb_host.u_phy._133_ ;
 wire \u_usb_host.u_phy._134_ ;
 wire \u_usb_host.u_phy._135_ ;
 wire \u_usb_host.u_phy._136_ ;
 wire \u_usb_host.u_phy._137_ ;
 wire \u_usb_host.u_phy._138_ ;
 wire \u_usb_host.u_phy._139_ ;
 wire \u_usb_host.u_phy._140_ ;
 wire \u_usb_host.u_phy._141_ ;
 wire \u_usb_host.u_phy._142_ ;
 wire \u_usb_host.u_phy._143_ ;
 wire \u_usb_host.u_phy._144_ ;
 wire \u_usb_host.u_phy._145_ ;
 wire \u_usb_host.u_phy._146_ ;
 wire \u_usb_host.u_phy._147_ ;
 wire \u_usb_host.u_phy._148_ ;
 wire \u_usb_host.u_phy._150_ ;
 wire \u_usb_host.u_phy._151_ ;
 wire \u_usb_host.u_phy._152_ ;
 wire \u_usb_host.u_phy._153_ ;
 wire \u_usb_host.u_phy._154_ ;
 wire \u_usb_host.u_phy._155_ ;
 wire \u_usb_host.u_phy._156_ ;
 wire \u_usb_host.u_phy._157_ ;
 wire \u_usb_host.u_phy._158_ ;
 wire \u_usb_host.u_phy._159_ ;
 wire \u_usb_host.u_phy._160_ ;
 wire \u_usb_host.u_phy._161_ ;
 wire \u_usb_host.u_phy._162_ ;
 wire \u_usb_host.u_phy._163_ ;
 wire \u_usb_host.u_phy._164_ ;
 wire \u_usb_host.u_phy._165_ ;
 wire \u_usb_host.u_phy._166_ ;
 wire \u_usb_host.u_phy._167_ ;
 wire \u_usb_host.u_phy._168_ ;
 wire \u_usb_host.u_phy._169_ ;
 wire \u_usb_host.u_phy._170_ ;
 wire \u_usb_host.u_phy._171_ ;
 wire \u_usb_host.u_phy._173_ ;
 wire \u_usb_host.u_phy._175_ ;
 wire \u_usb_host.u_phy._176_ ;
 wire \u_usb_host.u_phy._177_ ;
 wire \u_usb_host.u_phy._178_ ;
 wire \u_usb_host.u_phy._179_ ;
 wire \u_usb_host.u_phy._180_ ;
 wire \u_usb_host.u_phy._181_ ;
 wire \u_usb_host.u_phy._182_ ;
 wire \u_usb_host.u_phy._183_ ;
 wire \u_usb_host.u_phy._184_ ;
 wire \u_usb_host.u_phy._185_ ;
 wire \u_usb_host.u_phy._186_ ;
 wire \u_usb_host.u_phy._187_ ;
 wire \u_usb_host.u_phy._188_ ;
 wire \u_usb_host.u_phy._189_ ;
 wire \u_usb_host.u_phy._190_ ;
 wire \u_usb_host.u_phy._192_ ;
 wire \u_usb_host.u_phy._193_ ;
 wire \u_usb_host.u_phy.adjust_delayed_q ;
 wire \u_usb_host.u_phy.bit_count_q[0] ;
 wire \u_usb_host.u_phy.bit_count_q[1] ;
 wire \u_usb_host.u_phy.bit_count_q[2] ;
 wire \u_usb_host.u_phy.in_j_w ;
 wire \u_usb_host.u_phy.next_state_r[0] ;
 wire \u_usb_host.u_phy.next_state_r[1] ;
 wire \u_usb_host.u_phy.next_state_r[2] ;
 wire \u_usb_host.u_phy.next_state_r[3] ;
 wire \u_usb_host.u_phy.ones_count_q[0] ;
 wire \u_usb_host.u_phy.ones_count_q[1] ;
 wire \u_usb_host.u_phy.ones_count_q[2] ;
 wire \u_usb_host.u_phy.rx_dn0_q ;
 wire \u_usb_host.u_phy.rx_dn1_q ;
 wire \u_usb_host.u_phy.rx_dn_ms ;
 wire \u_usb_host.u_phy.rx_dn_q ;
 wire \u_usb_host.u_phy.rx_dp0_q ;
 wire \u_usb_host.u_phy.rx_dp1_q ;
 wire \u_usb_host.u_phy.rx_dp_ms ;
 wire \u_usb_host.u_phy.rx_dp_q ;
 wire \u_usb_host.u_phy.rxd0_q ;
 wire \u_usb_host.u_phy.rxd1_q ;
 wire \u_usb_host.u_phy.rxd_last_j_q ;
 wire \u_usb_host.u_phy.rxd_last_q ;
 wire \u_usb_host.u_phy.rxd_ms ;
 wire \u_usb_host.u_phy.rxd_q ;
 wire \u_usb_host.u_phy.sample_cnt_q[0] ;
 wire \u_usb_host.u_phy.sample_cnt_q[1] ;
 wire \u_usb_host.u_phy.sample_cnt_q[2] ;
 wire \u_usb_host.u_phy.send_eop_q ;
 wire \u_usb_host.u_phy.state_q[0] ;
 wire \u_usb_host.u_phy.state_q[1] ;
 wire \u_usb_host.u_phy.state_q[2] ;
 wire \u_usb_host.u_phy.state_q[3] ;
 wire \u_usb_host.u_phy.sync_j_detected_q ;
 wire \u_usb_host.u_phy.usb_rx_dn_i ;
 wire \u_usb_host.u_phy.usb_rx_dp_i ;
 wire \u_usb_host.u_phy.usb_rx_rcv_i ;
 wire \u_usb_host.u_phy.usb_tx_dn_o ;
 wire \u_usb_host.u_phy.usb_tx_dp_o ;
 wire \u_usb_host.u_phy.usb_tx_oen_o ;
 wire \u_usb_host.u_usb_rst.in_data_2s ;
 wire \u_usb_host.u_usb_rst.in_data_s ;
 wire \u_usb_host.u_usb_xcvr._0_ ;
 wire \u_usb_host.u_usb_xcvr._1_ ;
 wire \u_usb_host.u_wb_rst.in_data_2s ;
 wire \u_usb_host.u_wb_rst.in_data_s ;

 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_app_clk_A (.DIODE(app_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_0_u_usb_host.u_core._200__A  (.DIODE(\u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_usb_clk_A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_usb_clk_A (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_usb_clk_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_usb_clk_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_usb_clk_A (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_usb_clk_A (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_usb_clk_A (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_usb_clk_A (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_usb_clk_A (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_usb_clk_A (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_usb_clk_A (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_usb_clk_A (.DIODE(clknet_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_usb_clk_A (.DIODE(clknet_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_usb_clk_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_usb_clk_A (.DIODE(clknet_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_usb_clk_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_usb_clk_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_A (.DIODE(\u_usb_host.u_async_wb.s_cmd_rd_empty ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0563_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0563_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0560_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0559_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0559_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0559_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0556_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0554_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0554_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0554_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0526_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0526_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0524_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0524_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0522_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0520_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0520_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0518_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0515_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0515_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0514_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0514_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0512_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0512_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0509_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0509_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0497_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout261_A (.DIODE(\u_usb_host.u_async_wb.u_cmd_if.wr_reset_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout262_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout264_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout266_A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout268_A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout270_A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout272_A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout273_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout278_A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout282_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout285_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout288_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout290_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout291_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout292_A (.DIODE(\u_usb_host.u_async_wb.u_cmd_if.rd_reset_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout307_A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout308_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout309_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout310_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout312_A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout313_A (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout314_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout315_A (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout317_A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout318_A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout319_A (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout320_A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_A (.DIODE(\u_usb_host.u_core._117_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(\u_usb_host.u_core._117_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout93_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_A (.DIODE(\u_usb_host.u_core._095_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(\u_usb_host.u_core._095_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_A (.DIODE(\u_usb_host.u_async_wb.s_cmd_rd_empty ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2_A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold6_A (.DIODE(\u_usb_host.u_async_wb.u_cmd_if.wr_reset_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(reg_addr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(reg_addr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(reg_addr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(reg_addr[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(reg_cs));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(reg_wdata[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(reg_wdata[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(reg_wdata[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(reg_wdata[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(reg_wdata[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(cfg_cska_usb[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(reg_wdata[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(reg_wdata[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(reg_wdata[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(reg_wdata[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(reg_wdata[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(reg_wdata[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(reg_wdata[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(reg_wdata[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(reg_wdata[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(reg_wdata[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(cfg_cska_usb[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(reg_wdata[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(reg_wdata[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(reg_wdata[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(reg_wdata[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(reg_wdata[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(reg_wdata[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(reg_wdata[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(reg_wdata[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(reg_wdata[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(reg_wdata[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(cfg_cska_usb[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(reg_wdata[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(reg_wdata[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(reg_wdata[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(reg_wr));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(usb_in_dn));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(usb_in_dp));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(usb_rstn));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(wbd_clk_int));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(cfg_cska_usb[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(reg_addr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(reg_addr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(reg_addr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(reg_addr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(reg_addr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length3_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length4_A (.DIODE(clknet_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length5_A (.DIODE(clknet_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_output48_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._19__A_N  (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._20__A_N  (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._21__A_N  (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._22__A_N  (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._22__B  (.DIODE(\u_usb_host.u_async_wb.s_cmd_rd_data[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._23__A_N  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._24__A_N  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._25__A_N  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._26__A_N  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._27__A_N  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._28__A_N  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._29__A_N  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._30__A_N  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._31__A_N  (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._31__B  (.DIODE(\u_usb_host.u_async_wb.s_cmd_rd_data[16] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._32__A_N  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._32__B  (.DIODE(\u_usb_host.u_async_wb.s_cmd_rd_data[17] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._33__A_N  (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._33__B  (.DIODE(\u_usb_host.u_async_wb.s_cmd_rd_data[18] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._34__A_N  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._34__B  (.DIODE(\u_usb_host.u_async_wb.s_cmd_rd_data[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._58__D  (.DIODE(\u_usb_host.reg_ack ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._60__D  (.DIODE(\u_usb_host.reg_ack ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._60__RESET_B  (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._043__A  (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._044__A  (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._045__A  (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._045__B  (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._046__A  (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._046__B  (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._064__A  (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._069__A1  (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._070__A1  (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._084__S0  (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._084__S1  (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._085__S0  (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._085__S1  (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._086__S0  (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._086__S1  (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._087__S0  (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._087__S1  (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._088__S0  (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._088__S1  (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._089__S0  (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._089__S1  (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._090__S0  (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._090__S1  (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._091__S0  (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._091__S1  (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._092__S0  (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._092__S1  (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._093__S0  (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._093__S1  (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._094__S0  (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._094__S1  (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._095__S0  (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._095__S1  (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._096__S0  (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._096__S1  (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._097__S0  (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._097__S1  (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._098__S0  (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._098__S1  (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._099__S0  (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._099__S1  (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._100__S0  (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._100__S1  (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._101__S0  (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._101__S1  (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._102__S0  (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._102__S1  (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._103__S0  (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._103__S1  (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._104__S0  (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._104__S1  (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._105__S0  (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._105__S1  (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._106__S0  (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._106__S1  (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._107__S0  (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._107__S1  (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._112__S0  (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._112__S1  (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._113__S0  (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._113__S1  (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._114__S0  (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._114__S1  (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._115__S0  (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._115__S1  (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._116__S0  (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._116__S1  (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._117__S0  (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._117__S1  (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._118__S0  (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._118__S1  (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._119__S0  (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._119__S1  (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._120__S0  (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._120__S1  (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._121__S0  (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._121__S1  (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._122__S0  (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._122__S1  (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._131__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._132__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._133__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._134__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._135__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._136__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._136__D  (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._137__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._138__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._139__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._140__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._141__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._142__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._143__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._144__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._145__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._146__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._150__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._151__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._152__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._153__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._154__D  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._161__D  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._163__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._164__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._165__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._166__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._167__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._169__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._174__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._175__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._176__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._177__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._178__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._179__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._179__D  (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._180__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._181__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._182__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._183__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._184__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._185__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._186__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._187__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._188__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._189__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._191__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._194__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._195__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._197__D  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._204__D  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._206__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._207__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._208__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._209__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._210__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._212__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._217__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._218__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._219__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._220__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._221__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._222__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._222__D  (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._223__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._224__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._232__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._234__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._236__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._237__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._238__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._239__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._240__D  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._247__D  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._249__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._250__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._251__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._252__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._253__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._255__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._260__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._261__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._262__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._263__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._264__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._265__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._265__D  (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._266__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._267__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._268__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._269__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._270__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._271__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._272__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._273__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._274__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._275__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._276__CLK  (.DIODE(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._277__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._278__CLK  (.DIODE(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._279__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._280__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._281__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._282__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._283__CLK  (.DIODE(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._283__D  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._288__CLK  (.DIODE(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._289__CLK  (.DIODE(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._290__CLK  (.DIODE(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._290__D  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._291__CLK  (.DIODE(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._292__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._293__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._294__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._295__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._296__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._297__CLK  (.DIODE(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._298__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._317__CLK  (.DIODE(clknet_4_0_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._318__CLK  (.DIODE(clknet_4_0_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._319__CLK  (.DIODE(clknet_4_0_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._320__CLK  (.DIODE(clknet_4_0_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._321__CLK  (.DIODE(clknet_4_0_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._322__CLK  (.DIODE(clknet_4_0_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._323__CLK  (.DIODE(clknet_4_0_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._323__GATE  (.DIODE(\u_usb_host.reg_ack ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._326__CLK  (.DIODE(clknet_4_0_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._326__GATE  (.DIODE(\u_usb_host.reg_ack ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._021__A  (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._025__B  (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._033__A  (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._035__A1  (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._044__S  (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._056__S  (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._057__S  (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._058__S  (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._060__S  (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._063__S  (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._065__S  (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._074__B  (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._083__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._096__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._097__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._099__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._102__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._104__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._107__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._143__RESET_B  (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._144__RESET_B  (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._147__RESET_B  (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._148__RESET_B  (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._153__RESET_B  (.DIODE(\u_usb_host.u_async_wb.u_cmd_if.wr_reset_n ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._161__CLK  (.DIODE(clknet_4_2_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._161__GATE  (.DIODE(\u_usb_host.u_async_wb.u_resp_if._000_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._162__CLK  (.DIODE(clknet_4_2_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._162__GATE  (.DIODE(\u_usb_host.u_async_wb.u_resp_if._001_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._235__A  (.DIODE(\u_usb_host.u_core.cfg_wr ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._236__A  (.DIODE(\u_usb_host.u_core.fifo_flush_q ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._236__B  (.DIODE(\u_usb_host.u_core._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._237__A  (.DIODE(\u_usb_host.u_core.u_sie.utmi_linestate_i[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._237__B  (.DIODE(\u_usb_host.u_core.u_sie.utmi_linestate_i[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._250__A_N  (.DIODE(\u_usb_host.reg_ack ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._256__A  (.DIODE(\u_usb_host.u_core.cfg_wr ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._256__B  (.DIODE(\u_usb_host.u_core._092_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._258__A  (.DIODE(\u_usb_host.u_core.cfg_wr ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._258__B  (.DIODE(\u_usb_host.u_core._093_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._261__A  (.DIODE(\u_usb_host.u_core.cfg_wr ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._261__B  (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._327__A2  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._329__A2  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._331__A2  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._333__B1  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._335__B1  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._337__A2  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._339__A2  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._341__A2  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._342__A2  (.DIODE(\u_usb_host.u_core._092_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._342__B1  (.DIODE(\u_usb_host.u_core._096_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._342__B2  (.DIODE(\u_usb_host.u_core.u_fifo_rx.data_o[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._343__B1  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._345__B1  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._346__A2  (.DIODE(\u_usb_host.u_core._092_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._346__B1  (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._346__B2  (.DIODE(\u_usb_host.u_core.u_sie.utmi_linestate_i[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._348__A2  (.DIODE(\u_usb_host.u_core._093_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._348__B1  (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._349__A2  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._349__B1  (.DIODE(\u_usb_host.u_core._129_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._350__A2  (.DIODE(\u_usb_host.u_core._096_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._351__A2  (.DIODE(\u_usb_host.u_core._092_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._351__B1  (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._352__A2  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._352__B1  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._353__A2  (.DIODE(\u_usb_host.u_core._096_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._354__A2  (.DIODE(\u_usb_host.u_core._092_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._354__B1  (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._355__A2  (.DIODE(\u_usb_host.u_core._093_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._355__B1  (.DIODE(\u_usb_host.u_core._096_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._356__A2  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._357__A2  (.DIODE(\u_usb_host.u_core._092_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._357__B1  (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._358__A2  (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._358__B1  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._359__A2  (.DIODE(\u_usb_host.u_core._096_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._360__A2  (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._360__B1  (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._361__A2  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._361__B1  (.DIODE(\u_usb_host.u_core._129_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._362__A2  (.DIODE(\u_usb_host.u_core._092_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._362__B1  (.DIODE(\u_usb_host.u_core._093_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._363__A2  (.DIODE(\u_usb_host.u_core._096_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._364__A2  (.DIODE(\u_usb_host.u_core._092_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._364__B1  (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._365__A2  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._365__B1  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._366__A2  (.DIODE(\u_usb_host.u_core._096_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._367__A2  (.DIODE(\u_usb_host.u_core._093_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._368__A2  (.DIODE(\u_usb_host.u_core._092_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._368__B1  (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._368__B2  (.DIODE(\u_usb_host.u_core.u_sie.utmi_linestate_i[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._369__A2  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._369__B1  (.DIODE(\u_usb_host.u_core._129_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._370__A2  (.DIODE(\u_usb_host.u_core._096_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._372__A2  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._373__A2  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._373__B1  (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._374__A2  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._375__A2  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._376__A2  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._377__A2  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._378__A2  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._379__A2  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._380__A2  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._381__A2  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._382__A2  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._383__A2  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._384__A2  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._385__A2  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._385__B1  (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._386__A2  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._387__A2  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._387__B1  (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._388__A2  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._389__A2  (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._390__A2  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._391__A2  (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._392__A2  (.DIODE(\u_usb_host.u_core._117_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._393__A  (.DIODE(\u_usb_host.reg_ack ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._395__A  (.DIODE(\u_usb_host.u_core.cfg_wr ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._396__A  (.DIODE(\u_usb_host.u_core.cfg_wr ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._397__B  (.DIODE(\u_usb_host.u_core._157_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._398__B  (.DIODE(\u_usb_host.u_core._157_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._399__B  (.DIODE(\u_usb_host.u_core._157_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._400__B  (.DIODE(\u_usb_host.u_core._157_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._402__A  (.DIODE(\u_usb_host.u_core._096_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._428__RESET_B  (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._429__RESET_B  (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._430__CLK  (.DIODE(\clknet_1_1__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._432__CLK  (.DIODE(\clknet_1_1__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._433__CLK  (.DIODE(\clknet_1_1__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._438__CLK  (.DIODE(\clknet_1_1__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._439__CLK  (.DIODE(\clknet_1_1__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._440__CLK  (.DIODE(\clknet_1_1__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._441__CLK  (.DIODE(\clknet_1_1__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._442__CLK  (.DIODE(\clknet_1_1__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._443__CLK  (.DIODE(\clknet_1_1__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._445__RESET_B  (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._446__RESET_B  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._447__RESET_B  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._449__RESET_B  (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._454__RESET_B  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._466__RESET_B  (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._467__RESET_B  (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._468__RESET_B  (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._469__RESET_B  (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._470__RESET_B  (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._471__RESET_B  (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._486__RESET_B  (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._498__RESET_B  (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._506__RESET_B  (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._507__RESET_B  (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._508__RESET_B  (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._509__RESET_B  (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._510__RESET_B  (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._511__RESET_B  (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._512__RESET_B  (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._513__RESET_B  (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._514__RESET_B  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._519__RESET_B  (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._522__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._523__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._524__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._526__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._526__RESET_B  (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._527__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._528__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._529__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._530__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._531__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._532__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._533__CLK  (.DIODE(\clknet_2_2__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._534__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._535__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._538__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._542__RESET_B  (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._543__RESET_B  (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._547__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._548__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._549__CLK  (.DIODE(\clknet_2_0__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._552__RESET_B  (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._555__RESET_B  (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._556__CLK  (.DIODE(clknet_4_11_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._556__D  (.DIODE(\u_usb_host.u_core._025_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._558__CLK  (.DIODE(clknet_4_8_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._559__CLK  (.DIODE(clknet_4_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._560__RESET_B  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._563__CLK  (.DIODE(clknet_4_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._565__CLK  (.DIODE(clknet_4_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._566__RESET_B  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._567__CLK  (.DIODE(clknet_4_10_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._567__GATE  (.DIODE(\u_usb_host.u_core._025_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._568__CLK  (.DIODE(clknet_4_8_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._568__GATE  (.DIODE(\u_usb_host.u_core._025_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._569__CLK  (.DIODE(clknet_4_8_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._569__GATE  (.DIODE(\u_usb_host.u_core._025_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._570__CLK  (.DIODE(clknet_4_8_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._572__CLK  (.DIODE(clknet_4_8_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._574__CLK  (.DIODE(clknet_4_8_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._575__CLK  (.DIODE(clknet_4_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._576__GATE  (.DIODE(\u_usb_host.u_core._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._577__GATE  (.DIODE(\u_usb_host.u_core._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._578__GATE  (.DIODE(\u_usb_host.u_core._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._579__CLK  (.DIODE(clknet_4_2_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._579__GATE  (.DIODE(\u_usb_host.u_core._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._580__CLK  (.DIODE(clknet_4_8_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._580__GATE  (.DIODE(\u_usb_host.u_core._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._581__CLK  (.DIODE(clknet_4_8_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._581__GATE  (.DIODE(\u_usb_host.u_core._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._583__CLK  (.DIODE(clknet_4_8_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._583__GATE  (.DIODE(\u_usb_host.u_core._025_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._584__CLK  (.DIODE(clknet_4_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._589__CLK  (.DIODE(clknet_4_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._590__CLK  (.DIODE(clknet_4_11_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._592__CLK  (.DIODE(clknet_4_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._593__CLK  (.DIODE(clknet_4_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._595__CLK  (.DIODE(clknet_4_8_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._595__GATE  (.DIODE(\u_usb_host.u_core._025_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._596__CLK  (.DIODE(clknet_4_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._597__CLK  (.DIODE(clknet_4_2_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._598__CLK  (.DIODE(clknet_4_8_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._598__GATE  (.DIODE(\u_usb_host.u_core._025_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0797__A  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0798__A  (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0801__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0801__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0452_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0802__A  (.DIODE(\u_usb_host.u_core.fifo_flush_q ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0806__A  (.DIODE(\u_usb_host.u_core.fifo_flush_q ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0809__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0455_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0809__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0812__A  (.DIODE(\u_usb_host.u_core.fifo_flush_q ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0815__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0815__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0460_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0817__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0817__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0818__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0452_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0818__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0820__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0455_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0820__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0822__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0822__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0463_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0823__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0448_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0823__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0825__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0825__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0464_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0827__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0827__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0465_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0829__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0829__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0466_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0830__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0830__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0832__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0832__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0467_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0833__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0833__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0463_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0835__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0835__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0468_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0837__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0837__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0469_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0839__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0839__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0470_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0841__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0841__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0471_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0843__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0843__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0472_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0845__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0845__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0846__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0846__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0460_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0847__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0847__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0848__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0848__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0469_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0849__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0849__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0470_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0850__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0850__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0471_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0851__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0851__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0853__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0472_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0853__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0854__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0466_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0854__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0855__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0464_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0855__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0856__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0465_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0856__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0857__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0455_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0857__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0858__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0448_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0858__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0859__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0460_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0859__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0860__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0452_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0860__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0861__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0861__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0467_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0862__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0862__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0468_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0863__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0863__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0472_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0864__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0864__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0466_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0865__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0865__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0464_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0866__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0866__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0465_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0867__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0867__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0464_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0868__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0868__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0465_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0869__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0869__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0455_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0870__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0448_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0870__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0871__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0460_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0871__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0872__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0452_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0872__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0873__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0873__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0874__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0463_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0874__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0875__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0469_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0875__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0876__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0470_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0876__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0877__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0471_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0877__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0878__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0467_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0878__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0879__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0879__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0880__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0468_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0880__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0881__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0881__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0882__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0882__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0472_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0883__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0883__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0467_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0884__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0884__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0468_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0885__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0885__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0466_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0886__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0886__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0469_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0887__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0887__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0463_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0888__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0888__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0471_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0889__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0889__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0470_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0924__A1  (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0926__A2  (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0927__A2  (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0930__A2  (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0931__A1  (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0931__A2  (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0937__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0448_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0944__A  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0944__B  (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0945__A  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0945__B  (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0947__A  (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0947__B  (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0951__A  (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0951__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0514_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0953__C  (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0955__B  (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0955__C  (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0957__C  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0959__C  (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0961__B  (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0961__C  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0962__B  (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0963__B  (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0964__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0514_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0965__C  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0966__C  (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0968__B  (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0968__C  (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0969__C  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0970__A  (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0970__B  (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0971__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0522_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0972__A  (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0972__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0526_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0973__B  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0973__C  (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0976__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0518_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0977__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0526_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0978__C  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0979__B  (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0979__C  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0980__B  (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0981__B  (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0982__B  (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0983__C  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0984__A  (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0985__C  (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0986__A  (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0987__B  (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0991__C  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0992__C  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0995__C  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0996__A  (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0998__A  (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0998__B  (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0999__C  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1000__B  (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1001__A  (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1001__B  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1002__A  (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1002__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0556_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1003__A  (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1004__C  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1005__B  (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1006__B  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1007__B  (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1008__C  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1009__C  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1011__B  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1012__B  (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1013__C  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1014__B  (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1014__C  (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1015__C  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1016__C  (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1017__A  (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1017__B  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1026__A3  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1027__A3  (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1028__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0590_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1045__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0599_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1045__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0604_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1045__D  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0610_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1048__C  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1049__B  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1049__C  (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1050__C  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1052__B  (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1052__C  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1053__C  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1054__C  (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1056__B  (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1056__C  (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1057__C  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1058__B  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1058__C  (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1060__C  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1061__B  (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1061__C  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1063__B  (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1064__C  (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1065__C  (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1066__B  (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1066__C  (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1068__C  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1069__C  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1070__C  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1071__C  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1072__B  (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1073__C  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1074__B  (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1075__B  (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1076__B  (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1077__C  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1078__C  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1080__C  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1081__B  (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1081__C  (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1082__C  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1083__C  (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1092__A3  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1093__A3  (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1111__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0664_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1111__D  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0675_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1114__C  (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1117__B  (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1119__B  (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1121__C  (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1122__C  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1123__B  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1123__C  (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1124__B  (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1124__C  (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1126__C  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1127__B  (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1127__C  (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1129__C  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1130__C  (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1131__B  (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1131__C  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1132__B  (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1132__C  (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1134__C  (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1135__B  (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1135__C  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1136__C  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1137__C  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1138__B  (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1139__B  (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1139__C  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1141__B  (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1142__B  (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1145__C  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1147__B  (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1147__C  (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1149__C  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1150__B  (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1158__A2  (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1158__A3  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1159__A2  (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1159__A3  (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1160__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0090_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1177__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0099_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1177__D  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0110_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1180__C  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1181__C  (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1184__B  (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1188__C  (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1189__C  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1190__B  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1190__C  (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1192__C  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1193__B  (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1193__C  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1195__B  (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1196__B  (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1196__C  (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1197__C  (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1198__B  (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1200__B  (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1201__C  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1202__C  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1203__C  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1204__B  (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1206__B  (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1207__B  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1208__B  (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1210__C  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1212__C  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1213__B  (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1213__C  (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1214__B  (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1214__C  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1215__C  (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1224__A2  (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1224__A3  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1225__A2  (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1225__A3  (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1243__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0164_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1243__D  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0175_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1246__C  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1247__B  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1247__C  (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1250__B  (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1254__C  (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1255__C  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1256__B  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1256__C  (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1258__C  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1259__B  (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1259__C  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1261__B  (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1261__C  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1262__B  (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1262__C  (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1263__C  (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1264__B  (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1266__B  (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1267__C  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1268__B  (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1268__C  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1269__C  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1270__B  (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1272__B  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1273__B  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1274__B  (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1276__C  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1278__C  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1279__B  (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1279__C  (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1280__B  (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1280__C  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1281__C  (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1290__A2  (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1290__A3  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1291__A2  (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1291__A3  (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1292__D  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0223_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1309__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0229_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1309__D  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0240_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1311__C  (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1313__B  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1313__C  (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1320__C  (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1321__C  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1322__B  (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1322__C  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1323__B  (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1326__C  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1327__C  (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1328__C  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1329__B  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1329__C  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1330__B  (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1330__C  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1332__B  (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1333__C  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1334__B  (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1336__C  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1337__B  (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1340__B  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1341__B  (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1342__C  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1344__C  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1345__C  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1346__C  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1347__C  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1348__B  (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1348__C  (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1356__A3  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1357__A3  (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1375__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0294_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1375__D  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0305_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1378__C  (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1379__B  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1379__C  (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1382__B  (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1386__C  (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1387__C  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1388__C  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1390__C  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1391__B  (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1391__C  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1393__B  (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1394__C  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1395__C  (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1396__B  (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1396__C  (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1398__C  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1399__C  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1400__C  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1401__C  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1402__B  (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1403__C  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1405__B  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1406__B  (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1409__C  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1411__B  (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1411__C  (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1413__C  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1414__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0497_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1414__C  (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1422__A3  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1423__A3  (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1434__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0361_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1441__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0359_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1441__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0364_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1441__D  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0370_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1443__C  (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1445__C  (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1446__B  (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1446__C  (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1447__B  (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1452__C  (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1453__C  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1455__B  (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1458__C  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1459__B  (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1459__C  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1460__B  (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1460__C  (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1461__C  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1462__C  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1464__B  (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1464__C  (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1465__C  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1467__B  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1469__C  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1470__B  (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1473__B  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1474__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0497_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1475__C  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1477__C  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0560_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1478__C  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1479__C  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1480__C  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1481__B  (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1481__C  (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1489__A3  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1490__A3  (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1491__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0416_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1506__A2  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0509_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1508__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0425_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1508__D  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0436_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1510__D  (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1511__D  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1512__D  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1513__D  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1514__D  (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1515__D  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1516__D  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1517__D  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1518__D  (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1519__D  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1520__D  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1521__D  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1522__D  (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1523__D  (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1524__D  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1525__D  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1526__D  (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1527__D  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1528__D  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1529__D  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1530__D  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1531__D  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1532__D  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1533__D  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1534__D  (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1535__D  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1536__D  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1537__D  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1538__D  (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1539__D  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1540__D  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1541__D  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1542__D  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1543__D  (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1544__D  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1545__D  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1546__D  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1547__D  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1548__D  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1549__D  (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1550__D  (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1551__D  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1552__D  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1553__D  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1554__D  (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1555__D  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1556__D  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1557__D  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1558__D  (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1559__D  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1560__D  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1561__D  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1562__D  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1563__D  (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1564__D  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1565__D  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1566__D  (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1567__D  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1568__D  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1569__D  (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1570__D  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1571__D  (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1572__D  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1573__D  (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1574__D  (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1575__D  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1576__D  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1577__D  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1578__D  (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1579__D  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1580__D  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1581__D  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1582__D  (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1583__D  (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1584__D  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1585__D  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1586__D  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1587__D  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1588__D  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1589__D  (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1590__D  (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1591__D  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1592__D  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1593__D  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1594__D  (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1595__D  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1596__D  (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1597__D  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1598__D  (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1599__D  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1600__D  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1601__D  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1602__D  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1603__D  (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1604__D  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1605__D  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1606__D  (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1607__D  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1608__D  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1609__D  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1610__D  (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1611__D  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1612__D  (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1613__D  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1614__D  (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1615__D  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1616__D  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1617__D  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1618__D  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1619__D  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1620__D  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1621__D  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1622__D  (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1623__D  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1624__D  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1625__D  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1626__D  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1627__D  (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1628__D  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1629__D  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1630__D  (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1631__D  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1632__D  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1633__D  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1634__D  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1635__D  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1636__D  (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1637__D  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1638__D  (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1639__D  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1640__D  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1641__D  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1642__D  (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1643__D  (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1644__D  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1645__D  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1646__D  (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1647__D  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1648__D  (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1649__D  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1650__D  (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1651__D  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1652__D  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1653__D  (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1654__D  (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1655__D  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1656__D  (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1657__D  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1658__D  (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1659__D  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1660__D  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1661__D  (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1662__D  (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1663__D  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1664__D  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1665__D  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1666__D  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1667__D  (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1668__D  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1669__D  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1670__D  (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1671__D  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1672__D  (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1673__D  (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1674__D  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1675__D  (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1676__D  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1677__D  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1678__D  (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1679__D  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1680__D  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1681__D  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1682__D  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1683__D  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1684__D  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1685__D  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1686__D  (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1687__D  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1688__D  (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1689__D  (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1690__D  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1691__D  (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1692__D  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1693__D  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1694__D  (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1695__D  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1696__D  (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1697__D  (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1698__D  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1699__D  (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1700__D  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1701__D  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1702__D  (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1703__D  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1704__D  (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1705__D  (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1706__D  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1707__D  (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1708__D  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1709__D  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1710__D  (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1711__D  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1712__D  (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1713__D  (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1714__D  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1715__D  (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1716__D  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1717__D  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1718__D  (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1719__D  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1720__D  (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1721__D  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1722__D  (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1723__D  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1724__D  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1725__D  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1726__D  (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1727__D  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1728__D  (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1729__D  (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1730__D  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1731__D  (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1732__D  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1733__D  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1734__D  (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1735__D  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1736__D  (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1737__D  (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1738__D  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1739__D  (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1740__D  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1741__D  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1742__D  (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1743__D  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1744__D  (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1745__D  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1746__D  (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1747__D  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1748__D  (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1749__D  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1750__D  (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1751__D  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1752__D  (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1753__D  (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1754__D  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1755__D  (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1756__D  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1757__D  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1758__D  (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1759__D  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1760__D  (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1761__D  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1762__D  (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1763__D  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1764__D  (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1765__D  (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1766__D  (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1767__D  (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1768__D  (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1769__D  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1770__D  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1771__D  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1772__D  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1773__D  (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1774__D  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1775__D  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1776__D  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1777__D  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1778__D  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1779__D  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1780__D  (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1781__D  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1782__D  (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1783__D  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1784__D  (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1785__D  (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1786__D  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1787__D  (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1788__D  (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1789__D  (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1790__D  (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1791__D  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1792__D  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1793__D  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1794__D  (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1795__D  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1796__D  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1797__D  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1798__D  (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1799__D  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1800__D  (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1801__D  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1802__D  (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1803__D  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1804__D  (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1805__D  (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1806__D  (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1807__D  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1808__D  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1809__D  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1810__D  (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1811__D  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1812__D  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1813__D  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1814__D  (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1815__D  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1816__D  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1817__D  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1818__D  (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1819__D  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1820__D  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1821__D  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1822__D  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1823__D  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1824__D  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1825__D  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1826__D  (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1827__D  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1828__D  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1829__D  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1830__D  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1831__D  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1832__D  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1833__D  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1834__D  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1835__D  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1836__D  (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1837__D  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1838__D  (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1839__D  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1840__D  (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1841__D  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1842__D  (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1843__D  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1844__D  (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1845__D  (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1846__D  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1847__D  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1848__D  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1849__D  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1850__D  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1851__D  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1852__D  (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1853__D  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1854__D  (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1855__D  (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1856__D  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1857__D  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1858__D  (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1859__D  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1860__D  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1861__D  (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1862__D  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1863__D  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1864__D  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1865__D  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1866__D  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1867__D  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1868__D  (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1869__D  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1870__D  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1871__D  (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1872__D  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1873__D  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1874__D  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1875__D  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1876__D  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1877__D  (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1878__D  (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1879__D  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1880__D  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1881__D  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1882__D  (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1883__D  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1884__D  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1885__D  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1886__D  (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1887__D  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1888__D  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1889__D  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1890__D  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1891__D  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1892__D  (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1893__D  (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1898__RESET_B  (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1899__RESET_B  (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1900__RESET_B  (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1901__D  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1902__D  (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1903__D  (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1904__D  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1905__D  (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1906__D  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1907__D  (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1908__D  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1915__D  (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1916__D  (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1917__D  (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1918__D  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1919__D  (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1920__D  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1921__D  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1922__D  (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1923__CLK  (.DIODE(clknet_4_15_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1924__CLK  (.DIODE(clknet_4_12_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1925__CLK  (.DIODE(clknet_4_14_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1926__CLK  (.DIODE(clknet_4_12_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1930__CLK  (.DIODE(clknet_4_12_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1931__CLK  (.DIODE(clknet_4_14_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1932__CLK  (.DIODE(clknet_4_14_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1933__CLK  (.DIODE(clknet_4_14_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1934__CLK  (.DIODE(clknet_4_12_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1937__CLK  (.DIODE(clknet_4_14_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1938__CLK  (.DIODE(clknet_4_14_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1940__CLK  (.DIODE(clknet_4_4_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1942__CLK  (.DIODE(clknet_4_5_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1943__CLK  (.DIODE(clknet_4_4_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1944__CLK  (.DIODE(clknet_4_4_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1945__CLK  (.DIODE(clknet_4_4_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1946__CLK  (.DIODE(clknet_4_5_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1947__CLK  (.DIODE(clknet_4_5_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1948__CLK  (.DIODE(clknet_4_5_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1949__CLK  (.DIODE(clknet_4_14_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1950__CLK  (.DIODE(clknet_4_13_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1951__CLK  (.DIODE(clknet_4_13_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1952__CLK  (.DIODE(clknet_4_13_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1953__CLK  (.DIODE(clknet_4_5_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1954__CLK  (.DIODE(clknet_4_14_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1955__CLK  (.DIODE(clknet_4_14_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1957__CLK  (.DIODE(clknet_4_12_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1958__CLK  (.DIODE(clknet_4_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1959__CLK  (.DIODE(clknet_4_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1961__CLK  (.DIODE(clknet_4_5_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1962__CLK  (.DIODE(clknet_4_12_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1963__CLK  (.DIODE(clknet_4_15_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1964__CLK  (.DIODE(clknet_4_15_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1965__CLK  (.DIODE(clknet_4_15_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1966__CLK  (.DIODE(clknet_4_15_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1967__CLK  (.DIODE(clknet_4_15_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1968__CLK  (.DIODE(clknet_4_15_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1969__CLK  (.DIODE(clknet_4_14_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1970__CLK  (.DIODE(clknet_4_15_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1971__CLK  (.DIODE(clknet_4_5_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1972__CLK  (.DIODE(clknet_4_5_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1973__CLK  (.DIODE(clknet_4_5_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1974__CLK  (.DIODE(clknet_4_5_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1975__CLK  (.DIODE(clknet_4_4_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1976__CLK  (.DIODE(clknet_4_4_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1977__CLK  (.DIODE(clknet_4_4_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1978__CLK  (.DIODE(clknet_4_5_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1979__CLK  (.DIODE(clknet_4_4_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1980__CLK  (.DIODE(clknet_4_13_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1981__CLK  (.DIODE(clknet_4_13_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1982__CLK  (.DIODE(clknet_4_15_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1983__CLK  (.DIODE(clknet_4_13_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1984__CLK  (.DIODE(clknet_4_13_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1985__CLK  (.DIODE(clknet_4_15_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1986__CLK  (.DIODE(clknet_4_13_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1987__CLK  (.DIODE(clknet_4_15_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1988__CLK  (.DIODE(clknet_4_12_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1989__CLK  (.DIODE(clknet_4_12_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1990__D  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1991__D  (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1992__D  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1993__D  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1994__D  (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1995__D  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1996__D  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1997__D  (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1999__RESET_B  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2002__RESET_B  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2003__RESET_B  (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2004__D  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2005__D  (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2006__D  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2007__D  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2008__D  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2009__D  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2010__D  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2011__D  (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2012__D  (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2013__D  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2014__D  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2015__D  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2016__D  (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2017__D  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2018__D  (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2019__D  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2020__D  (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2021__D  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2022__D  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2023__D  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2024__D  (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2025__D  (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2026__D  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2027__D  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2028__D  (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2029__D  (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2030__D  (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2031__D  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2032__D  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2033__D  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2034__D  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2035__D  (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2036__D  (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2037__D  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2038__D  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2039__D  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2040__D  (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2041__D  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2042__D  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2043__D  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2044__D  (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2045__D  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2046__D  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2047__D  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2048__D  (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2049__D  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2050__D  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2051__D  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2052__D  (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2053__D  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2054__D  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2055__D  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2056__D  (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2057__D  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2058__D  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2059__D  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2060__D  (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2061__D  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2062__D  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2063__D  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2064__D  (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2065__D  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2066__D  (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2067__D  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2068__D  (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2069__D  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2070__D  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2071__D  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2072__D  (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2073__D  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2074__D  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2075__D  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2076__D  (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2077__D  (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2078__D  (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2079__D  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2080__D  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2081__D  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2082__D  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2083__D  (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2084__D  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2085__D  (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2086__D  (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2087__D  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2088__D  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2089__D  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2090__D  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2091__D  (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2092__D  (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2093__D  (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2094__D  (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2095__D  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2096__D  (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2097__D  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2098__D  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2099__D  (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2100__D  (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2101__D  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2102__D  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2103__D  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2104__D  (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2105__D  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2106__D  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2107__D  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._34__CLK  (.DIODE(clknet_4_11_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._226__B  (.DIODE(\u_usb_host.u_phy._049_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._235__A1  (.DIODE(\u_usb_host.u_phy._049_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._238__A1_N  (.DIODE(\u_usb_host.u_phy._049_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._253__B  (.DIODE(\u_usb_host.u_phy._086_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._256__A  (.DIODE(\u_usb_host.u_phy._049_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._257__A  (.DIODE(\u_usb_host.u_phy._049_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._263__C_N  (.DIODE(\u_usb_host.u_phy._086_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._320__B2  (.DIODE(\u_usb_host.u_phy._049_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._321__A0  (.DIODE(\u_usb_host.u_phy.usb_tx_dp_o ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._329__A2  (.DIODE(\u_usb_host.u_phy._049_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._336__A  (.DIODE(\u_usb_host.u_phy._049_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._366__A  (.DIODE(\u_usb_host.u_phy.usb_tx_dp_o ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._372__B  (.DIODE(\u_usb_host.u_phy._049_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._380__RESET_B  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._383__RESET_B  (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._384__RESET_B  (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._385__RESET_B  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._386__RESET_B  (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._395__RESET_B  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._397__RESET_B  (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._409__RESET_B  (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._419__CLK  (.DIODE(clknet_4_10_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._419__RESET_B  (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._420__CLK  (.DIODE(clknet_4_10_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._420__RESET_B  (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._421__CLK  (.DIODE(clknet_4_10_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._421__RESET_B  (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._422__CLK  (.DIODE(clknet_4_10_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._423__CLK  (.DIODE(clknet_4_10_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._424__CLK  (.DIODE(clknet_4_10_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._425__CLK  (.DIODE(clknet_4_10_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._426__CLK  (.DIODE(clknet_4_10_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._426__RESET_B  (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._427__CLK  (.DIODE(clknet_4_10_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._428__CLK  (.DIODE(clknet_4_10_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._430__CLK  (.DIODE(clknet_4_10_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._432__CLK  (.DIODE(clknet_4_11_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._433__CLK  (.DIODE(clknet_4_10_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._434__CLK  (.DIODE(clknet_4_10_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._435__CLK  (.DIODE(clknet_4_10_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._436__CLK  (.DIODE(clknet_4_10_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._437__CLK  (.DIODE(clknet_4_11_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._438__CLK  (.DIODE(clknet_4_11_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._439__CLK  (.DIODE(clknet_4_10_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._440__CLK  (.DIODE(clknet_4_11_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._441__CLK  (.DIODE(clknet_4_11_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._442__CLK  (.DIODE(clknet_4_11_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._443__CLK  (.DIODE(clknet_4_11_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._444__CLK  (.DIODE(clknet_4_11_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._445__CLK  (.DIODE(clknet_4_11_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._446__CLK  (.DIODE(clknet_4_10_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._447__CLK  (.DIODE(clknet_4_10_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_usb_rst._1__CLK  (.DIODE(clknet_4_0_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_usb_rst._1__RESET_B  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_usb_rst._2__CLK  (.DIODE(clknet_4_0_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_usb_rst._2__RESET_B  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_usb_rst.u_buf.genblk1.u_mux_A1  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_usb_xcvr._4__A  (.DIODE(\u_usb_host.u_phy.usb_tx_dp_o ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_usb_xcvr._6__B1  (.DIODE(\u_usb_host.u_phy.usb_tx_dp_o ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_wb_rst._1__RESET_B  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_wb_rst._2__RESET_B  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_wb_rst.u_buf.genblk1.u_mux_A1  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1_A (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2_A (.DIODE(usb_clk));
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_989 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__clkbuf_1 _01_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[0] ),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 _02_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[1] ),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 _03_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[2] ),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 _04_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[3] ),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 _05_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[4] ),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _06_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[5] ),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _07_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[6] ),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 _08_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[7] ),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 _09_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[8] ),
    .X(net79));
 sky130_fd_sc_hd__and4bb_1 _0_ (.A_N(net11),
    .B_N(net13),
    .C(net14),
    .D(net12),
    .X(\u_usb_host.u_async_wb.wbm_cyc_i ));
 sky130_fd_sc_hd__clkbuf_1 _10_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[9] ),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _11_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[10] ),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 _12_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[11] ),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 _13_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[12] ),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 _14_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[13] ),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 _15_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[14] ),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 _16_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[15] ),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 _17_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[16] ),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 _18_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[17] ),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 _19_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[18] ),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 _20_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[19] ),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 _21_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[20] ),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 _22_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[21] ),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 _23_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[22] ),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 _24_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[23] ),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 _25_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[24] ),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 _26_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[25] ),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 _27_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[26] ),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 _28_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[27] ),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 _29_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[28] ),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 _30_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[29] ),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 _31_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[30] ),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 _32_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[31] ),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_app_clk (.A(app_clk),
    .X(clknet_0_app_clk));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_cmd_if._033_  (.A(\u_usb_host.u_async_wb.u_cmd_if._033_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._033_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_cmd_if._034_  (.A(\u_usb_host.u_async_wb.u_cmd_if._034_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._034_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_cmd_if._035_  (.A(\u_usb_host.u_async_wb.u_cmd_if._035_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._035_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_cmd_if._036_  (.A(\u_usb_host.u_async_wb.u_cmd_if._036_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._036_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_cmd_if._037_  (.A(\u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_cmd_if._038_  (.A(\u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_cmd_if._039_  (.A(\u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_cmd_if._040_  (.A(\u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_resp_if._014_  (.A(\u_usb_host.u_async_wb.u_resp_if._014_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_resp_if._014_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_resp_if._015_  (.A(\u_usb_host.u_async_wb.u_resp_if._015_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_resp_if._015_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_resp_if._016_  (.A(\u_usb_host.u_async_wb.u_resp_if._016_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_resp_if._016_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_resp_if._017_  (.A(\u_usb_host.u_async_wb.u_resp_if._017_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_resp_if._017_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_resp_if._018_  (.A(\u_usb_host.u_async_wb.u_resp_if._018_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_resp_if._018_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_resp_if._019_  (.A(\u_usb_host.u_async_wb.u_resp_if._019_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_resp_if._019_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core._171_  (.A(\u_usb_host.u_core._171_ ),
    .X(\clknet_0_u_usb_host.u_core._171_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core._172_  (.A(\u_usb_host.u_core._172_ ),
    .X(\clknet_0_u_usb_host.u_core._172_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core._178_  (.A(\u_usb_host.u_core._178_ ),
    .X(\clknet_0_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core._183_  (.A(\u_usb_host.u_core._183_ ),
    .X(\clknet_0_u_usb_host.u_core._183_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core._184_  (.A(\u_usb_host.u_core._184_ ),
    .X(\clknet_0_u_usb_host.u_core._184_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core._185_  (.A(\u_usb_host.u_core._185_ ),
    .X(\clknet_0_u_usb_host.u_core._185_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core._193_  (.A(\u_usb_host.u_core._193_ ),
    .X(\clknet_0_u_usb_host.u_core._193_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core._200_  (.A(\u_usb_host.u_core._200_ ),
    .X(\clknet_0_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0717_  (.A(\u_usb_host.u_core.u_fifo_rx._0717_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0717_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0718_  (.A(\u_usb_host.u_core.u_fifo_rx._0718_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0718_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0719_  (.A(\u_usb_host.u_core.u_fifo_rx._0719_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0719_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0720_  (.A(\u_usb_host.u_core.u_fifo_rx._0720_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0720_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0721_  (.A(\u_usb_host.u_core.u_fifo_rx._0721_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0721_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0722_  (.A(\u_usb_host.u_core.u_fifo_rx._0722_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0722_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0723_  (.A(\u_usb_host.u_core.u_fifo_rx._0723_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0723_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0724_  (.A(\u_usb_host.u_core.u_fifo_rx._0724_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0724_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0725_  (.A(\u_usb_host.u_core.u_fifo_rx._0725_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0725_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0726_  (.A(\u_usb_host.u_core.u_fifo_rx._0726_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0726_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0727_  (.A(\u_usb_host.u_core.u_fifo_rx._0727_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0727_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0728_  (.A(\u_usb_host.u_core.u_fifo_rx._0728_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0728_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0729_  (.A(\u_usb_host.u_core.u_fifo_rx._0729_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0729_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0730_  (.A(\u_usb_host.u_core.u_fifo_rx._0730_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0730_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0731_  (.A(\u_usb_host.u_core.u_fifo_rx._0731_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0731_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0732_  (.A(\u_usb_host.u_core.u_fifo_rx._0732_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0732_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0733_  (.A(\u_usb_host.u_core.u_fifo_rx._0733_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0733_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0734_  (.A(\u_usb_host.u_core.u_fifo_rx._0734_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0734_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0735_  (.A(\u_usb_host.u_core.u_fifo_rx._0735_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0735_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0736_  (.A(\u_usb_host.u_core.u_fifo_rx._0736_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0736_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0737_  (.A(\u_usb_host.u_core.u_fifo_rx._0737_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0737_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0738_  (.A(\u_usb_host.u_core.u_fifo_rx._0738_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0738_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0739_  (.A(\u_usb_host.u_core.u_fifo_rx._0739_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0739_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0740_  (.A(\u_usb_host.u_core.u_fifo_rx._0740_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0740_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0741_  (.A(\u_usb_host.u_core.u_fifo_rx._0741_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0741_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0742_  (.A(\u_usb_host.u_core.u_fifo_rx._0742_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0742_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0743_  (.A(\u_usb_host.u_core.u_fifo_rx._0743_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0743_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0744_  (.A(\u_usb_host.u_core.u_fifo_rx._0744_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0744_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0745_  (.A(\u_usb_host.u_core.u_fifo_rx._0745_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0745_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0746_  (.A(\u_usb_host.u_core.u_fifo_rx._0746_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0746_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0747_  (.A(\u_usb_host.u_core.u_fifo_rx._0747_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0747_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0748_  (.A(\u_usb_host.u_core.u_fifo_rx._0748_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0748_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0749_  (.A(\u_usb_host.u_core.u_fifo_rx._0749_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0749_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0750_  (.A(\u_usb_host.u_core.u_fifo_rx._0750_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0750_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0751_  (.A(\u_usb_host.u_core.u_fifo_rx._0751_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0751_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0752_  (.A(\u_usb_host.u_core.u_fifo_rx._0752_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0752_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0753_  (.A(\u_usb_host.u_core.u_fifo_rx._0753_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0753_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0754_  (.A(\u_usb_host.u_core.u_fifo_rx._0754_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0754_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0755_  (.A(\u_usb_host.u_core.u_fifo_rx._0755_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0755_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0756_  (.A(\u_usb_host.u_core.u_fifo_rx._0756_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0756_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0757_  (.A(\u_usb_host.u_core.u_fifo_rx._0757_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0757_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0758_  (.A(\u_usb_host.u_core.u_fifo_rx._0758_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0758_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0759_  (.A(\u_usb_host.u_core.u_fifo_rx._0759_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0759_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0760_  (.A(\u_usb_host.u_core.u_fifo_rx._0760_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0760_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0761_  (.A(\u_usb_host.u_core.u_fifo_rx._0761_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0761_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0762_  (.A(\u_usb_host.u_core.u_fifo_rx._0762_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0762_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0763_  (.A(\u_usb_host.u_core.u_fifo_rx._0763_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0763_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0764_  (.A(\u_usb_host.u_core.u_fifo_rx._0764_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0764_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0765_  (.A(\u_usb_host.u_core.u_fifo_rx._0765_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0765_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0766_  (.A(\u_usb_host.u_core.u_fifo_rx._0766_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0766_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0767_  (.A(\u_usb_host.u_core.u_fifo_rx._0767_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0767_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0768_  (.A(\u_usb_host.u_core.u_fifo_rx._0768_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0768_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0769_  (.A(\u_usb_host.u_core.u_fifo_rx._0769_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0769_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0770_  (.A(\u_usb_host.u_core.u_fifo_rx._0770_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0770_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0771_  (.A(\u_usb_host.u_core.u_fifo_rx._0771_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0771_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0772_  (.A(\u_usb_host.u_core.u_fifo_rx._0772_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0772_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0773_  (.A(\u_usb_host.u_core.u_fifo_rx._0773_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0773_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0774_  (.A(\u_usb_host.u_core.u_fifo_rx._0774_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0774_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0775_  (.A(\u_usb_host.u_core.u_fifo_rx._0775_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0775_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0776_  (.A(\u_usb_host.u_core.u_fifo_rx._0776_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0776_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0777_  (.A(\u_usb_host.u_core.u_fifo_rx._0777_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0777_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0778_  (.A(\u_usb_host.u_core.u_fifo_rx._0778_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0778_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0779_  (.A(\u_usb_host.u_core.u_fifo_rx._0779_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0779_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0780_  (.A(\u_usb_host.u_core.u_fifo_rx._0780_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0780_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0781_  (.A(\u_usb_host.u_core.u_fifo_rx._0781_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0781_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0782_  (.A(\u_usb_host.u_core.u_fifo_rx._0782_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0782_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0783_  (.A(\u_usb_host.u_core.u_fifo_rx._0783_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0783_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_sie._00_  (.A(\u_usb_host.u_core.u_sie._00_ ),
    .X(\clknet_0_u_usb_host.u_core.u_sie._00_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_phy._175_  (.A(\u_usb_host.u_phy._175_ ),
    .X(\clknet_0_u_usb_host.u_phy._175_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_phy._178_  (.A(\u_usb_host.u_phy._178_ ),
    .X(\clknet_0_u_usb_host.u_phy._178_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_phy._180_  (.A(\u_usb_host.u_phy._180_ ),
    .X(\clknet_0_u_usb_host.u_phy._180_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_phy._187_  (.A(\u_usb_host.u_phy._187_ ),
    .X(\clknet_0_u_usb_host.u_phy._187_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_phy._188_  (.A(\u_usb_host.u_phy._188_ ),
    .X(\clknet_0_u_usb_host.u_phy._188_ ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_usb_clk (.A(net380),
    .X(clknet_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_app_clk (.A(clknet_0_app_clk),
    .X(clknet_1_0__leaf_app_clk));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_async_wb.u_cmd_if._033_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._033_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._033_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_async_wb.u_cmd_if._034_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._034_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._034_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_async_wb.u_cmd_if._035_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._035_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._035_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_async_wb.u_cmd_if._036_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._036_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._036_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_async_wb.u_resp_if._014_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._014_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._014_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_async_wb.u_resp_if._015_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._015_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._015_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_async_wb.u_resp_if._016_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._016_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._016_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_async_wb.u_resp_if._017_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._017_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._017_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core._171_  (.A(\clknet_0_u_usb_host.u_core._171_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core._171_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core._172_  (.A(\clknet_0_u_usb_host.u_core._172_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core._172_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core._178_  (.A(\clknet_0_u_usb_host.u_core._178_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core._183_  (.A(\clknet_0_u_usb_host.u_core._183_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core._183_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core._184_  (.A(\clknet_0_u_usb_host.u_core._184_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core._184_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core._185_  (.A(\clknet_0_u_usb_host.u_core._185_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core._185_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core._193_  (.A(\clknet_0_u_usb_host.u_core._193_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core._193_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0717_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0717_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0717_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0718_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0718_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0718_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0719_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0719_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0719_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0720_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0720_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0720_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0721_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0721_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0722_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0722_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0723_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0723_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0724_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0724_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0725_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0725_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0726_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0726_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0727_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0727_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0728_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0728_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0729_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0729_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0730_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0730_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0731_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0731_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0732_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0732_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0733_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0733_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0734_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0734_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0735_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0735_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0736_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0736_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0737_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0737_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0738_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0738_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0739_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0739_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0740_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0740_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0741_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0741_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0742_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0742_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0743_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0743_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0744_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0744_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0745_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0745_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0746_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0746_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0747_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0747_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0748_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0748_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0749_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0749_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0750_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0750_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0751_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0751_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0752_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0752_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0753_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0753_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0754_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0754_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0755_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0755_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0756_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0756_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0757_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0757_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0758_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0758_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0759_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0759_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0760_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0760_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0761_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0761_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0762_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0762_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0763_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0763_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0764_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0764_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0765_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0765_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0766_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0766_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0767_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0767_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0768_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0768_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0769_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0769_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0770_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0770_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0771_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0771_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0772_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0772_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0773_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0773_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0774_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0774_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0775_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0775_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0776_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0776_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0777_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0777_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0778_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0778_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0779_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0779_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0780_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0780_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0781_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0781_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0782_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0782_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0783_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0783_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_phy._175_  (.A(\clknet_0_u_usb_host.u_phy._175_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_phy._175_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_phy._178_  (.A(\clknet_0_u_usb_host.u_phy._178_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_phy._178_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_phy._180_  (.A(\clknet_0_u_usb_host.u_phy._180_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_phy._180_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_phy._187_  (.A(\clknet_0_u_usb_host.u_phy._187_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_phy._187_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_phy._188_  (.A(\clknet_0_u_usb_host.u_phy._188_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_phy._188_ ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_app_clk (.A(clknet_0_app_clk),
    .X(clknet_1_1__leaf_app_clk));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_async_wb.u_cmd_if._033_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._033_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._033_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_async_wb.u_cmd_if._034_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._034_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._034_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_async_wb.u_cmd_if._035_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._035_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._035_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_async_wb.u_cmd_if._036_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._036_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._036_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_async_wb.u_resp_if._014_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._014_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._014_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_async_wb.u_resp_if._015_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._015_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._015_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_async_wb.u_resp_if._016_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._016_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._016_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_async_wb.u_resp_if._017_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._017_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._017_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core._171_  (.A(\clknet_0_u_usb_host.u_core._171_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core._171_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core._172_  (.A(\clknet_0_u_usb_host.u_core._172_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core._172_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core._178_  (.A(\clknet_0_u_usb_host.u_core._178_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core._183_  (.A(\clknet_0_u_usb_host.u_core._183_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core._183_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core._184_  (.A(\clknet_0_u_usb_host.u_core._184_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core._184_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core._185_  (.A(\clknet_0_u_usb_host.u_core._185_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core._185_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core._193_  (.A(\clknet_0_u_usb_host.u_core._193_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core._193_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0717_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0717_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0717_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0718_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0718_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0718_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0719_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0719_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0719_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0720_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0720_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0720_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0721_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0721_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0722_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0722_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0723_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0723_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0724_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0724_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0725_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0725_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0726_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0726_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0727_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0727_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0728_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0728_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0729_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0729_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0730_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0730_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0731_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0731_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0732_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0732_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0733_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0733_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0734_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0734_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0735_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0735_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0736_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0736_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0737_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0737_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0738_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0738_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0739_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0739_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0740_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0740_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0741_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0741_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0742_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0742_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0743_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0743_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0744_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0744_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0745_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0745_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0746_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0746_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0747_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0747_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0748_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0748_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0749_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0749_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0750_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0750_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0751_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0751_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0752_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0752_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0753_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0753_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0754_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0754_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0755_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0755_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0756_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0756_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0757_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0757_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0758_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0758_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0759_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0759_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0760_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0760_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0761_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0761_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0762_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0762_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0763_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0763_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0764_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0764_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0765_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0765_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0766_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0766_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0767_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0767_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0768_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0768_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0769_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0769_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0770_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0770_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0771_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0771_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0772_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0772_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0773_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0773_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0774_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0774_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0775_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0775_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0776_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0776_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0777_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0777_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0778_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0778_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0779_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0779_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0780_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0780_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0781_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0781_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0782_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0782_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0783_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0783_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_phy._175_  (.A(\clknet_0_u_usb_host.u_phy._175_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_phy._175_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_phy._178_  (.A(\clknet_0_u_usb_host.u_phy._178_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_phy._178_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_phy._180_  (.A(\clknet_0_u_usb_host.u_phy._180_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_phy._180_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_phy._187_  (.A(\clknet_0_u_usb_host.u_phy._187_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_phy._187_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_phy._188_  (.A(\clknet_0_u_usb_host.u_phy._188_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_phy._188_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_u_usb_host.u_async_wb.u_cmd_if._037_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .X(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_u_usb_host.u_async_wb.u_cmd_if._038_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .X(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_u_usb_host.u_async_wb.u_cmd_if._039_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .X(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_u_usb_host.u_async_wb.u_cmd_if._040_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .X(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_u_usb_host.u_async_wb.u_resp_if._018_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .X(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_u_usb_host.u_async_wb.u_resp_if._019_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .X(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_u_usb_host.u_core._200_  (.A(\clknet_0_u_usb_host.u_core._200_ ),
    .X(\clknet_2_0__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_u_usb_host.u_core.u_sie._00_  (.A(\clknet_0_u_usb_host.u_core.u_sie._00_ ),
    .X(\clknet_2_0__leaf_u_usb_host.u_core.u_sie._00_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_u_usb_host.u_async_wb.u_cmd_if._037_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .X(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_u_usb_host.u_async_wb.u_cmd_if._038_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .X(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_u_usb_host.u_async_wb.u_cmd_if._039_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .X(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_u_usb_host.u_async_wb.u_cmd_if._040_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .X(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_u_usb_host.u_async_wb.u_resp_if._018_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .X(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_u_usb_host.u_async_wb.u_resp_if._019_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .X(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_u_usb_host.u_core._200_  (.A(\clknet_0_u_usb_host.u_core._200_ ),
    .X(\clknet_2_1__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_u_usb_host.u_core.u_sie._00_  (.A(\clknet_0_u_usb_host.u_core.u_sie._00_ ),
    .X(\clknet_2_1__leaf_u_usb_host.u_core.u_sie._00_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_u_usb_host.u_async_wb.u_cmd_if._037_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .X(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_u_usb_host.u_async_wb.u_cmd_if._038_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .X(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_u_usb_host.u_async_wb.u_cmd_if._039_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .X(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_u_usb_host.u_async_wb.u_cmd_if._040_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .X(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_u_usb_host.u_async_wb.u_resp_if._018_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .X(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_u_usb_host.u_async_wb.u_resp_if._019_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .X(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_u_usb_host.u_core._200_  (.A(\clknet_0_u_usb_host.u_core._200_ ),
    .X(\clknet_2_2__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_u_usb_host.u_core.u_sie._00_  (.A(\clknet_0_u_usb_host.u_core.u_sie._00_ ),
    .X(\clknet_2_2__leaf_u_usb_host.u_core.u_sie._00_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_u_usb_host.u_async_wb.u_cmd_if._037_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .X(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_u_usb_host.u_async_wb.u_cmd_if._038_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .X(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_u_usb_host.u_async_wb.u_cmd_if._039_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .X(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_u_usb_host.u_async_wb.u_cmd_if._040_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .X(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_u_usb_host.u_async_wb.u_resp_if._018_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .X(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_u_usb_host.u_async_wb.u_resp_if._019_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .X(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_u_usb_host.u_core._200_  (.A(\clknet_0_u_usb_host.u_core._200_ ),
    .X(\clknet_2_3__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_u_usb_host.u_core.u_sie._00_  (.A(\clknet_0_u_usb_host.u_core.u_sie._00_ ),
    .X(\clknet_2_3__leaf_u_usb_host.u_core.u_sie._00_ ));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_usb_clk (.A(net382),
    .X(clknet_4_0_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_usb_clk (.A(net384),
    .X(clknet_4_10_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_usb_clk (.A(net384),
    .X(clknet_4_11_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_usb_clk (.A(net383),
    .X(clknet_4_12_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_usb_clk (.A(net383),
    .X(clknet_4_13_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_usb_clk (.A(net383),
    .X(clknet_4_14_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_usb_clk (.A(net383),
    .X(clknet_4_15_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_usb_clk (.A(net382),
    .X(clknet_4_1_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_usb_clk (.A(net382),
    .X(clknet_4_2_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_usb_clk (.A(net382),
    .X(clknet_4_3_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_usb_clk (.A(clknet_0_usb_clk),
    .X(clknet_4_4_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_usb_clk (.A(clknet_0_usb_clk),
    .X(clknet_4_5_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_usb_clk (.A(net384),
    .X(clknet_4_6_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_usb_clk (.A(clknet_0_usb_clk),
    .X(clknet_4_7_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_usb_clk (.A(net384),
    .X(clknet_4_8_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_usb_clk (.A(net384),
    .X(clknet_4_9_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_2 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 fanout101 (.A(\u_usb_host.u_async_wb.s_cmd_rd_empty ),
    .X(net101));
 sky130_fd_sc_hd__buf_2 fanout102 (.A(\u_usb_host.u_phy._050_ ),
    .X(net102));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout103 (.A(\u_usb_host.u_phy._050_ ),
    .X(net103));
 sky130_fd_sc_hd__buf_2 fanout104 (.A(net106),
    .X(net104));
 sky130_fd_sc_hd__buf_2 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_4 fanout106 (.A(\u_usb_host.u_core.fifo_rx_data_w[7] ),
    .X(net106));
 sky130_fd_sc_hd__buf_2 fanout107 (.A(net111),
    .X(net107));
 sky130_fd_sc_hd__buf_2 fanout108 (.A(net111),
    .X(net108));
 sky130_fd_sc_hd__buf_2 fanout109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__buf_2 fanout110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__buf_2 fanout111 (.A(\u_usb_host.u_core.fifo_rx_data_w[7] ),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_4 fanout112 (.A(net120),
    .X(net112));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout113 (.A(net120),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_4 fanout114 (.A(net120),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 fanout115 (.A(net120),
    .X(net115));
 sky130_fd_sc_hd__buf_2 fanout116 (.A(net120),
    .X(net116));
 sky130_fd_sc_hd__buf_2 fanout117 (.A(net120),
    .X(net117));
 sky130_fd_sc_hd__buf_2 fanout118 (.A(net119),
    .X(net118));
 sky130_fd_sc_hd__buf_2 fanout119 (.A(net120),
    .X(net119));
 sky130_fd_sc_hd__buf_4 fanout120 (.A(\u_usb_host.u_core.fifo_rx_data_w[6] ),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_4 fanout121 (.A(net124),
    .X(net121));
 sky130_fd_sc_hd__buf_2 fanout122 (.A(net124),
    .X(net122));
 sky130_fd_sc_hd__buf_2 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__buf_2 fanout124 (.A(\u_usb_host.u_core.fifo_rx_data_w[5] ),
    .X(net124));
 sky130_fd_sc_hd__buf_2 fanout125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__buf_2 fanout126 (.A(\u_usb_host.u_core.fifo_rx_data_w[5] ),
    .X(net126));
 sky130_fd_sc_hd__buf_2 fanout127 (.A(\u_usb_host.u_core.fifo_rx_data_w[5] ),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 fanout128 (.A(\u_usb_host.u_core.fifo_rx_data_w[5] ),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_4 fanout129 (.A(net132),
    .X(net129));
 sky130_fd_sc_hd__buf_2 fanout130 (.A(net132),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_4 fanout131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__buf_2 fanout132 (.A(\u_usb_host.u_core.fifo_rx_data_w[4] ),
    .X(net132));
 sky130_fd_sc_hd__buf_2 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_4 fanout134 (.A(net136),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_4 fanout135 (.A(net136),
    .X(net135));
 sky130_fd_sc_hd__buf_4 fanout136 (.A(\u_usb_host.u_core.fifo_rx_data_w[4] ),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_4 fanout137 (.A(net140),
    .X(net137));
 sky130_fd_sc_hd__buf_2 fanout138 (.A(net140),
    .X(net138));
 sky130_fd_sc_hd__buf_2 fanout139 (.A(net140),
    .X(net139));
 sky130_fd_sc_hd__buf_2 fanout140 (.A(\u_usb_host.u_core.fifo_rx_data_w[3] ),
    .X(net140));
 sky130_fd_sc_hd__buf_2 fanout141 (.A(net142),
    .X(net141));
 sky130_fd_sc_hd__buf_2 fanout142 (.A(\u_usb_host.u_core.fifo_rx_data_w[3] ),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_4 fanout143 (.A(\u_usb_host.u_core.fifo_rx_data_w[3] ),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 fanout144 (.A(\u_usb_host.u_core.fifo_rx_data_w[3] ),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_4 fanout145 (.A(net148),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 fanout146 (.A(net148),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_4 fanout147 (.A(net148),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 fanout148 (.A(\u_usb_host.u_core.fifo_rx_data_w[2] ),
    .X(net148));
 sky130_fd_sc_hd__buf_2 fanout149 (.A(net150),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 fanout150 (.A(\u_usb_host.u_core.fifo_rx_data_w[2] ),
    .X(net150));
 sky130_fd_sc_hd__buf_2 fanout151 (.A(\u_usb_host.u_core.fifo_rx_data_w[2] ),
    .X(net151));
 sky130_fd_sc_hd__buf_2 fanout152 (.A(\u_usb_host.u_core.fifo_rx_data_w[2] ),
    .X(net152));
 sky130_fd_sc_hd__buf_2 fanout153 (.A(net161),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_2 fanout154 (.A(net161),
    .X(net154));
 sky130_fd_sc_hd__buf_2 fanout155 (.A(net161),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 fanout156 (.A(net160),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 fanout157 (.A(net160),
    .X(net157));
 sky130_fd_sc_hd__buf_2 fanout158 (.A(net159),
    .X(net158));
 sky130_fd_sc_hd__buf_2 fanout159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_2 fanout160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_4 fanout161 (.A(\u_usb_host.u_core.fifo_rx_data_w[1] ),
    .X(net161));
 sky130_fd_sc_hd__buf_2 fanout162 (.A(net169),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 fanout163 (.A(net169),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_4 fanout164 (.A(net169),
    .X(net164));
 sky130_fd_sc_hd__buf_2 fanout165 (.A(net169),
    .X(net165));
 sky130_fd_sc_hd__buf_2 fanout166 (.A(net169),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_4 fanout167 (.A(net169),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_2 fanout168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__buf_4 fanout169 (.A(\u_usb_host.u_core.fifo_rx_data_w[0] ),
    .X(net169));
 sky130_fd_sc_hd__buf_2 fanout170 (.A(\u_usb_host.u_core.u_fifo_rx._0563_ ),
    .X(net170));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout171 (.A(\u_usb_host.u_core.u_fifo_rx._0563_ ),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_4 fanout172 (.A(\u_usb_host.u_core.u_fifo_rx._0560_ ),
    .X(net172));
 sky130_fd_sc_hd__buf_2 fanout173 (.A(\u_usb_host.u_core.u_fifo_rx._0559_ ),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 fanout174 (.A(\u_usb_host.u_core.u_fifo_rx._0559_ ),
    .X(net174));
 sky130_fd_sc_hd__buf_2 fanout175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__buf_2 fanout176 (.A(\u_usb_host.u_core.u_fifo_rx._0559_ ),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_2 fanout177 (.A(net179),
    .X(net177));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout178 (.A(net179),
    .X(net178));
 sky130_fd_sc_hd__buf_2 fanout179 (.A(\u_usb_host.u_core.u_fifo_rx._0556_ ),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_2 fanout181 (.A(\u_usb_host.u_core.u_fifo_rx._0554_ ),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_2 fanout182 (.A(\u_usb_host.u_core.u_fifo_rx._0554_ ),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 fanout183 (.A(\u_usb_host.u_core.u_fifo_rx._0554_ ),
    .X(net183));
 sky130_fd_sc_hd__buf_2 fanout184 (.A(net186),
    .X(net184));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout185 (.A(net186),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_2 fanout186 (.A(net188),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_4 fanout187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_2 fanout188 (.A(\u_usb_host.u_core.u_fifo_rx._0541_ ),
    .X(net188));
 sky130_fd_sc_hd__buf_2 fanout189 (.A(\u_usb_host.u_core.u_fifo_rx._0526_ ),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 fanout190 (.A(\u_usb_host.u_core.u_fifo_rx._0526_ ),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_4 fanout191 (.A(\u_usb_host.u_core.u_fifo_rx._0524_ ),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_2 fanout192 (.A(\u_usb_host.u_core.u_fifo_rx._0524_ ),
    .X(net192));
 sky130_fd_sc_hd__buf_2 fanout193 (.A(net195),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 fanout194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_4 fanout195 (.A(\u_usb_host.u_core.u_fifo_rx._0522_ ),
    .X(net195));
 sky130_fd_sc_hd__buf_2 fanout196 (.A(\u_usb_host.u_core.u_fifo_rx._0520_ ),
    .X(net196));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout197 (.A(\u_usb_host.u_core.u_fifo_rx._0520_ ),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 fanout198 (.A(net200),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 fanout199 (.A(net200),
    .X(net199));
 sky130_fd_sc_hd__buf_2 fanout200 (.A(\u_usb_host.u_core.u_fifo_rx._0518_ ),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_2 fanout201 (.A(net202),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_2 fanout202 (.A(net208),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 fanout203 (.A(net205),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_2 fanout204 (.A(net205),
    .X(net204));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout205 (.A(net208),
    .X(net205));
 sky130_fd_sc_hd__buf_2 fanout206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__buf_2 fanout207 (.A(net208),
    .X(net207));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout208 (.A(\u_usb_host.u_core.u_fifo_rx._0515_ ),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_2 fanout209 (.A(net215),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_2 fanout210 (.A(net215),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_2 fanout211 (.A(net215),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_2 fanout212 (.A(net214),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_2 fanout213 (.A(net214),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_2 fanout214 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_2 fanout215 (.A(net216),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_2 fanout216 (.A(\u_usb_host.u_core.u_fifo_rx._0515_ ),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_2 fanout217 (.A(\u_usb_host.u_core.u_fifo_rx._0514_ ),
    .X(net217));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout218 (.A(\u_usb_host.u_core.u_fifo_rx._0514_ ),
    .X(net218));
 sky130_fd_sc_hd__buf_2 fanout219 (.A(\u_usb_host.u_core.u_fifo_rx._0512_ ),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_2 fanout220 (.A(\u_usb_host.u_core.u_fifo_rx._0512_ ),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_2 fanout221 (.A(net223),
    .X(net221));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__buf_2 fanout223 (.A(net224),
    .X(net223));
 sky130_fd_sc_hd__buf_2 fanout224 (.A(\u_usb_host.u_core.u_fifo_rx._0509_ ),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_2 fanout225 (.A(net226),
    .X(net225));
 sky130_fd_sc_hd__buf_2 fanout226 (.A(\u_usb_host.u_core.u_fifo_rx._0509_ ),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_2 fanout227 (.A(net229),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_1 fanout228 (.A(net229),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_4 fanout229 (.A(\u_usb_host.u_core.u_fifo_rx._0508_ ),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_2 fanout230 (.A(net243),
    .X(net230));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout231 (.A(net243),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_2 fanout232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 fanout233 (.A(net243),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_2 fanout234 (.A(net243),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_2 fanout235 (.A(net243),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_2 fanout236 (.A(net237),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_2 fanout237 (.A(net242),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_2 fanout238 (.A(net240),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_1 fanout239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout240 (.A(net242),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 fanout241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_2 fanout242 (.A(net243),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_4 fanout243 (.A(\u_usb_host.u_core.u_fifo_rx._0502_ ),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_2 fanout244 (.A(net254),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_1 fanout245 (.A(net254),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_2 fanout246 (.A(net247),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 fanout247 (.A(net248),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_2 fanout248 (.A(net249),
    .X(net248));
 sky130_fd_sc_hd__buf_2 fanout249 (.A(net254),
    .X(net249));
 sky130_fd_sc_hd__buf_2 fanout250 (.A(net252),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_1 fanout251 (.A(net252),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_2 fanout252 (.A(net253),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_2 fanout253 (.A(net254),
    .X(net253));
 sky130_fd_sc_hd__buf_2 fanout254 (.A(\u_usb_host.u_core.u_fifo_rx._0501_ ),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_2 fanout255 (.A(net257),
    .X(net255));
 sky130_fd_sc_hd__buf_2 fanout256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__buf_2 fanout257 (.A(net258),
    .X(net257));
 sky130_fd_sc_hd__buf_2 fanout258 (.A(\u_usb_host.u_core.u_fifo_rx._0499_ ),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_4 fanout259 (.A(\u_usb_host.u_core.u_fifo_rx._0497_ ),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_4 fanout260 (.A(net261),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_4 fanout261 (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_reset_n ),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_4 fanout262 (.A(net264),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_2 fanout263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_4 fanout264 (.A(net292),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_4 fanout265 (.A(net271),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_4 fanout266 (.A(net271),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_4 fanout267 (.A(net268),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_2 fanout268 (.A(net271),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_4 fanout269 (.A(net270),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_4 fanout270 (.A(net271),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_4 fanout271 (.A(net292),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_4 fanout272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_2 fanout273 (.A(net291),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_4 fanout274 (.A(net277),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_4 fanout275 (.A(net277),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_4 fanout276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_2 fanout277 (.A(net291),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_4 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__buf_4 fanout279 (.A(net291),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_4 fanout280 (.A(net282),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_4 fanout281 (.A(net285),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_2 fanout282 (.A(net285),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_4 fanout283 (.A(net284),
    .X(net283));
 sky130_fd_sc_hd__buf_4 fanout284 (.A(net285),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_4 fanout285 (.A(net291),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_4 fanout286 (.A(net287),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_4 fanout287 (.A(net288),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_2 fanout288 (.A(net291),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_4 fanout289 (.A(net290),
    .X(net289));
 sky130_fd_sc_hd__buf_2 fanout290 (.A(net291),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_4 fanout291 (.A(net292),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_4 fanout292 (.A(\u_usb_host.u_async_wb.u_cmd_if.rd_reset_n ),
    .X(net292));
 sky130_fd_sc_hd__buf_2 fanout293 (.A(\u_usb_host.u_phy.state_q[3] ),
    .X(net293));
 sky130_fd_sc_hd__buf_2 fanout294 (.A(\u_usb_host.u_phy.state_q[1] ),
    .X(net294));
 sky130_fd_sc_hd__buf_2 fanout295 (.A(\u_usb_host.u_phy.state_q[0] ),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_2 fanout296 (.A(net297),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_2 fanout297 (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[3] ),
    .X(net297));
 sky130_fd_sc_hd__buf_2 fanout298 (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[2] ),
    .X(net298));
 sky130_fd_sc_hd__buf_2 fanout299 (.A(\u_usb_host.u_core.u_fifo_rx.rd_ptr[3] ),
    .X(net299));
 sky130_fd_sc_hd__buf_2 fanout300 (.A(\u_usb_host.u_core.u_fifo_rx.rd_ptr[3] ),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_2 fanout301 (.A(\u_usb_host.u_core.u_fifo_rx.rd_ptr[2] ),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_4 fanout302 (.A(\u_usb_host.u_core.u_fifo_rx.rd_ptr[2] ),
    .X(net302));
 sky130_fd_sc_hd__buf_2 fanout303 (.A(net304),
    .X(net303));
 sky130_fd_sc_hd__buf_2 fanout304 (.A(\u_usb_host.u_core.u_fifo_rx.rd_ptr[1] ),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_2 fanout305 (.A(net306),
    .X(net305));
 sky130_fd_sc_hd__buf_2 fanout306 (.A(\u_usb_host.u_core.u_fifo_rx.rd_ptr[0] ),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_4 fanout307 (.A(net308),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_4 fanout308 (.A(net386),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_4 fanout309 (.A(net386),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_2 fanout310 (.A(net386),
    .X(net310));
 sky130_fd_sc_hd__buf_4 fanout311 (.A(net385),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_4 fanout312 (.A(net313),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_4 fanout313 (.A(net316),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_4 fanout314 (.A(net315),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_4 fanout315 (.A(net316),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_4 fanout316 (.A(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[1] ),
    .X(net316));
 sky130_fd_sc_hd__buf_4 fanout317 (.A(net318),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_4 fanout318 (.A(net321),
    .X(net318));
 sky130_fd_sc_hd__buf_4 fanout319 (.A(net320),
    .X(net319));
 sky130_fd_sc_hd__buf_4 fanout320 (.A(net321),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_4 fanout321 (.A(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[0] ),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_4 fanout86 (.A(\u_usb_host.u_core._117_ ),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_4 fanout87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__buf_2 fanout88 (.A(\u_usb_host.u_core._117_ ),
    .X(net88));
 sky130_fd_sc_hd__buf_2 fanout89 (.A(net91),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_4 fanout90 (.A(net91),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 fanout91 (.A(\u_usb_host.u_core._086_ ),
    .X(net91));
 sky130_fd_sc_hd__buf_2 fanout92 (.A(net94),
    .X(net92));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout93 (.A(net94),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 fanout94 (.A(\u_usb_host.u_core._116_ ),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_4 fanout95 (.A(\u_usb_host.u_core._095_ ),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 fanout96 (.A(\u_usb_host.u_core._095_ ),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 fanout97 (.A(net99),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 fanout99 (.A(\u_usb_host.u_async_wb.s_cmd_rd_empty ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net388),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\u_usb_host.u_core._140_ ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_0[1] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_0[0] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_0[0] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_0[1] ),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_0[2] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\u_usb_host.u_wb_rst.in_data_s ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\u_usb_host.u_core.u_sie.utmi_data_i[0] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\u_usb_host.u_phy.rxd_ms ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\u_usb_host.u_phy.rx_dp_ms ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\u_usb_host.u_core.reg_rdata_r[2] ),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\u_usb_host.u_core.utmi_termselect_o ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\u_usb_host.u_core.intr_done_q ),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\u_usb_host.u_core.reg_rdata_r[1] ),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\u_usb_host.reg_rdata[17] ),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\u_usb_host.reg_rdata[16] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\u_usb_host.reg_rdata[24] ),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\u_usb_host.reg_rdata[26] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\u_usb_host.reg_rdata[13] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net311),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\u_usb_host.reg_rdata[9] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\u_usb_host.reg_rdata[29] ),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\u_usb_host.reg_rdata[14] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\u_usb_host.reg_rdata[10] ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\u_usb_host.reg_rdata[31] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\u_usb_host.u_core.utmi_dppulldown_o ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\u_usb_host.reg_rdata[7] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\u_usb_host.reg_rdata[23] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\u_usb_host.reg_rdata[28] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\u_usb_host.u_core.usb_irq_mask_device_detect_out_w ),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net310),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\u_usb_host.reg_rdata[12] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\u_usb_host.reg_rdata[15] ),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\u_usb_host.reg_rdata[21] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\u_usb_host.u_core.sof_irq_q ),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\u_usb_host.reg_rdata[18] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\u_usb_host.reg_rdata[3] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\u_usb_host.reg_rdata[4] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\u_usb_host.reg_rdata[30] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\u_usb_host.reg_rdata[5] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\u_usb_host.reg_rdata[11] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\u_usb_host.u_async_wb.u_resp_if.rd_ptr[0] ),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\u_usb_host.reg_rdata[0] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\u_usb_host.reg_rdata[8] ),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\u_usb_host.u_core.intr_sof_q ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\u_usb_host.u_core._131_ ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\u_usb_host.u_core.reg_rdata_r[0] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\u_usb_host.u_core.utmi_dmpulldown_o ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\u_usb_host.reg_rdata[6] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\u_usb_host.reg_rdata[27] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\u_usb_host.reg_rdata[2] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\u_usb_host.reg_rdata[1] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\u_usb_host.u_wb_rst.in_data_2s ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\u_usb_host.reg_rdata[25] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\u_usb_host.reg_rdata[20] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\u_usb_host.u_phy.sync_j_detected_q ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\u_usb_host.reg_rdata[19] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\u_usb_host.u_phy.rxd_last_q ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\u_usb_host.reg_rdata[22] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\u_usb_host.u_core.u_sie.utmi_data_i[6] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\u_usb_host.u_core.u_sie.utmi_data_i[4] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\u_usb_host.u_core.u_sie.utmi_data_i[2] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\u_usb_host.u_core.u_sie.utmi_data_i[7] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_reset_n ),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\u_usb_host.u_core.u_sie.utmi_data_i[1] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\u_usb_host.u_core.u_sie.utmi_data_i[3] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\u_usb_host.u_core.u_sie.utmi_data_i[5] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\u_usb_host.u_core.u_sie.data_idx_i ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\u_usb_host.u_core.usb_xfer_token_ack_out_w ),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\u_usb_host.u_core.usb_ctrl_wr_q ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\u_usb_host.u_core.usb_xfer_token_in_out_w ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\u_usb_host.u_core.usb_ctrl_enable_sof_out_w ),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[18] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\u_usb_host.u_core.transfer_start_q ),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\u_usb_host.u_usb_rst.in_data_2s ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[20] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[21] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[19] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[22] ),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[17] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[23] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[16] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\u_usb_host.u_phy.rxd_last_j_q ),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[28] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[10] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\u_usb_host.u_core.usb_rx_stat_start_pend_in_w ),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[12] ),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[11] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[27] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_0[1] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_0[0] ),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[31] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[14] ),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[9] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[13] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[26] ),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\u_usb_host.u_core.usb_irq_mask_err_out_w ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[25] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[15] ),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[29] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_0[2] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[24] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_0[1] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[30] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_0[0] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\u_usb_host.u_usb_rst.in_data_s ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[8] ),
    .X(net483));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(cfg_cska_usb[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(reg_addr[5]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(reg_addr[6]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(reg_addr[7]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(reg_addr[8]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(reg_cs),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(reg_wdata[0]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(reg_wdata[10]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(reg_wdata[11]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(reg_wdata[12]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(reg_wdata[13]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(cfg_cska_usb[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(reg_wdata[14]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(reg_wdata[15]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(reg_wdata[16]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(reg_wdata[17]),
    .X(net23));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(reg_wdata[18]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(reg_wdata[19]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(reg_wdata[1]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(reg_wdata[20]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(reg_wdata[21]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(reg_wdata[22]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(cfg_cska_usb[2]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input30 (.A(reg_wdata[23]),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(reg_wdata[28]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(reg_wdata[29]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(reg_wdata[2]),
    .X(net33));
 sky130_fd_sc_hd__dlymetal6s2s_1 input34 (.A(reg_wdata[30]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(reg_wdata[31]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(reg_wdata[3]),
    .X(net36));
 sky130_fd_sc_hd__dlymetal6s2s_1 input37 (.A(reg_wdata[4]),
    .X(net37));
 sky130_fd_sc_hd__dlymetal6s2s_1 input38 (.A(reg_wdata[5]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(reg_wdata[6]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(cfg_cska_usb[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(reg_wdata[7]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(reg_wdata[8]),
    .X(net41));
 sky130_fd_sc_hd__dlymetal6s2s_1 input42 (.A(reg_wdata[9]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(reg_wr),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(usb_in_dn),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(usb_in_dp),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 input46 (.A(usb_rstn),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(wbd_clk_int),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(reg_addr[0]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(reg_addr[1]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(reg_addr[2]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(reg_addr[3]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(reg_addr[4]),
    .X(net9));
 sky130_fd_sc_hd__buf_6 max_length3 (.A(net384),
    .X(net382));
 sky130_fd_sc_hd__buf_4 max_length4 (.A(clknet_0_usb_clk),
    .X(net383));
 sky130_fd_sc_hd__buf_6 max_length5 (.A(clknet_0_usb_clk),
    .X(net384));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(reg_ack));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(reg_rdata[0]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(reg_rdata[10]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(reg_rdata[11]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(reg_rdata[12]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(reg_rdata[13]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(reg_rdata[14]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(reg_rdata[15]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(reg_rdata[16]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(reg_rdata[17]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(reg_rdata[18]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(reg_rdata[19]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(reg_rdata[1]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(reg_rdata[20]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(reg_rdata[21]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(reg_rdata[22]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(reg_rdata[23]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(reg_rdata[24]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(reg_rdata[25]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(reg_rdata[26]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(reg_rdata[27]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(reg_rdata[28]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(reg_rdata[29]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(reg_rdata[2]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(reg_rdata[30]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(reg_rdata[31]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(reg_rdata[3]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(reg_rdata[4]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(reg_rdata[5]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(reg_rdata[6]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(reg_rdata[7]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(reg_rdata[8]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(reg_rdata[9]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(usb_intr_o));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(usb_out_dn));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(usb_out_dp));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(usb_out_tx_oen));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(wbd_clk_usb));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_1.u_dly0  (.A(\u_skew_usb.clk_inbuf ),
    .X(\u_skew_usb.clkbuf_1.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_1.u_dly1  (.A(\u_skew_usb.clkbuf_1.X1 ),
    .X(\u_skew_usb.clkbuf_1.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_1.u_dly2  (.A(\u_skew_usb.clkbuf_1.X2 ),
    .X(\u_skew_usb.clkbuf_1.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_1.u_dly3  (.A(\u_skew_usb.clkbuf_1.X3 ),
    .X(\u_skew_usb.clk_d1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_10.u_dly0  (.A(\u_skew_usb.clk_d9 ),
    .X(\u_skew_usb.clkbuf_10.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_10.u_dly1  (.A(\u_skew_usb.clkbuf_10.X1 ),
    .X(\u_skew_usb.clkbuf_10.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_10.u_dly2  (.A(\u_skew_usb.clkbuf_10.X2 ),
    .X(\u_skew_usb.clkbuf_10.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_10.u_dly3  (.A(\u_skew_usb.clkbuf_10.X3 ),
    .X(\u_skew_usb.clk_d10 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_11.u_dly0  (.A(\u_skew_usb.clk_d10 ),
    .X(\u_skew_usb.clkbuf_11.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_11.u_dly1  (.A(\u_skew_usb.clkbuf_11.X1 ),
    .X(\u_skew_usb.clkbuf_11.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_11.u_dly2  (.A(\u_skew_usb.clkbuf_11.X2 ),
    .X(\u_skew_usb.clkbuf_11.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_11.u_dly3  (.A(\u_skew_usb.clkbuf_11.X3 ),
    .X(\u_skew_usb.clk_d11 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_12.u_dly0  (.A(\u_skew_usb.clk_d11 ),
    .X(\u_skew_usb.clkbuf_12.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_12.u_dly1  (.A(\u_skew_usb.clkbuf_12.X1 ),
    .X(\u_skew_usb.clkbuf_12.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_12.u_dly2  (.A(\u_skew_usb.clkbuf_12.X2 ),
    .X(\u_skew_usb.clkbuf_12.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_12.u_dly3  (.A(\u_skew_usb.clkbuf_12.X3 ),
    .X(\u_skew_usb.clk_d12 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_13.u_dly0  (.A(\u_skew_usb.clk_d12 ),
    .X(\u_skew_usb.clkbuf_13.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_13.u_dly1  (.A(\u_skew_usb.clkbuf_13.X1 ),
    .X(\u_skew_usb.clkbuf_13.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_13.u_dly2  (.A(\u_skew_usb.clkbuf_13.X2 ),
    .X(\u_skew_usb.clkbuf_13.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_13.u_dly3  (.A(\u_skew_usb.clkbuf_13.X3 ),
    .X(\u_skew_usb.clk_d13 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_14.u_dly0  (.A(\u_skew_usb.clk_d13 ),
    .X(\u_skew_usb.clkbuf_14.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_14.u_dly1  (.A(\u_skew_usb.clkbuf_14.X1 ),
    .X(\u_skew_usb.clkbuf_14.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_14.u_dly2  (.A(\u_skew_usb.clkbuf_14.X2 ),
    .X(\u_skew_usb.clkbuf_14.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_14.u_dly3  (.A(\u_skew_usb.clkbuf_14.X3 ),
    .X(\u_skew_usb.clk_d14 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_15.u_dly0  (.A(\u_skew_usb.clk_d14 ),
    .X(\u_skew_usb.clkbuf_15.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_15.u_dly1  (.A(\u_skew_usb.clkbuf_15.X1 ),
    .X(\u_skew_usb.clkbuf_15.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_15.u_dly2  (.A(\u_skew_usb.clkbuf_15.X2 ),
    .X(\u_skew_usb.clkbuf_15.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_15.u_dly3  (.A(\u_skew_usb.clkbuf_15.X3 ),
    .X(\u_skew_usb.clk_d15 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_2.u_dly0  (.A(\u_skew_usb.clk_d1 ),
    .X(\u_skew_usb.clkbuf_2.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_2.u_dly1  (.A(\u_skew_usb.clkbuf_2.X1 ),
    .X(\u_skew_usb.clkbuf_2.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_2.u_dly2  (.A(\u_skew_usb.clkbuf_2.X2 ),
    .X(\u_skew_usb.clkbuf_2.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_2.u_dly3  (.A(\u_skew_usb.clkbuf_2.X3 ),
    .X(\u_skew_usb.clk_d2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_3.u_dly0  (.A(\u_skew_usb.clk_d2 ),
    .X(\u_skew_usb.clkbuf_3.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_3.u_dly1  (.A(\u_skew_usb.clkbuf_3.X1 ),
    .X(\u_skew_usb.clkbuf_3.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_3.u_dly2  (.A(\u_skew_usb.clkbuf_3.X2 ),
    .X(\u_skew_usb.clkbuf_3.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_3.u_dly3  (.A(\u_skew_usb.clkbuf_3.X3 ),
    .X(\u_skew_usb.clk_d3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_4.u_dly0  (.A(\u_skew_usb.clk_d3 ),
    .X(\u_skew_usb.clkbuf_4.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_4.u_dly1  (.A(\u_skew_usb.clkbuf_4.X1 ),
    .X(\u_skew_usb.clkbuf_4.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_4.u_dly2  (.A(\u_skew_usb.clkbuf_4.X2 ),
    .X(\u_skew_usb.clkbuf_4.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_4.u_dly3  (.A(\u_skew_usb.clkbuf_4.X3 ),
    .X(\u_skew_usb.clk_d4 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_5.u_dly0  (.A(\u_skew_usb.clk_d4 ),
    .X(\u_skew_usb.clkbuf_5.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_5.u_dly1  (.A(\u_skew_usb.clkbuf_5.X1 ),
    .X(\u_skew_usb.clkbuf_5.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_5.u_dly2  (.A(\u_skew_usb.clkbuf_5.X2 ),
    .X(\u_skew_usb.clkbuf_5.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_5.u_dly3  (.A(\u_skew_usb.clkbuf_5.X3 ),
    .X(\u_skew_usb.clk_d5 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_6.u_dly0  (.A(\u_skew_usb.clk_d5 ),
    .X(\u_skew_usb.clkbuf_6.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_6.u_dly1  (.A(\u_skew_usb.clkbuf_6.X1 ),
    .X(\u_skew_usb.clkbuf_6.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_6.u_dly2  (.A(\u_skew_usb.clkbuf_6.X2 ),
    .X(\u_skew_usb.clkbuf_6.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_6.u_dly3  (.A(\u_skew_usb.clkbuf_6.X3 ),
    .X(\u_skew_usb.clk_d6 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_7.u_dly0  (.A(\u_skew_usb.clk_d6 ),
    .X(\u_skew_usb.clkbuf_7.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_7.u_dly1  (.A(\u_skew_usb.clkbuf_7.X1 ),
    .X(\u_skew_usb.clkbuf_7.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_7.u_dly2  (.A(\u_skew_usb.clkbuf_7.X2 ),
    .X(\u_skew_usb.clkbuf_7.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_7.u_dly3  (.A(\u_skew_usb.clkbuf_7.X3 ),
    .X(\u_skew_usb.clk_d7 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_8.u_dly0  (.A(\u_skew_usb.clk_d7 ),
    .X(\u_skew_usb.clkbuf_8.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_8.u_dly1  (.A(\u_skew_usb.clkbuf_8.X1 ),
    .X(\u_skew_usb.clkbuf_8.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_8.u_dly2  (.A(\u_skew_usb.clkbuf_8.X2 ),
    .X(\u_skew_usb.clkbuf_8.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_8.u_dly3  (.A(\u_skew_usb.clkbuf_8.X3 ),
    .X(\u_skew_usb.clk_d8 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_9.u_dly0  (.A(\u_skew_usb.clk_d8 ),
    .X(\u_skew_usb.clkbuf_9.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_9.u_dly1  (.A(\u_skew_usb.clkbuf_9.X1 ),
    .X(\u_skew_usb.clkbuf_9.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_9.u_dly2  (.A(\u_skew_usb.clkbuf_9.X2 ),
    .X(\u_skew_usb.clkbuf_9.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_9.u_dly3  (.A(\u_skew_usb.clkbuf_9.X3 ),
    .X(\u_skew_usb.clk_d9 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_clkbuf_in.u_buf  (.A(net47),
    .X(\u_skew_usb.clk_inbuf ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_clkbuf_out.u_buf  (.A(\u_skew_usb.d30 ),
    .X(net85));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_00.genblk1.u_mux  (.A0(\u_skew_usb.in0 ),
    .A1(\u_skew_usb.in1 ),
    .S(net1),
    .X(\u_skew_usb.d00 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_01.genblk1.u_mux  (.A0(\u_skew_usb.in2 ),
    .A1(\u_skew_usb.in3 ),
    .S(net1),
    .X(\u_skew_usb.d01 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_02.genblk1.u_mux  (.A0(\u_skew_usb.in4 ),
    .A1(\u_skew_usb.in5 ),
    .S(net1),
    .X(\u_skew_usb.d02 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_03.genblk1.u_mux  (.A0(\u_skew_usb.in6 ),
    .A1(\u_skew_usb.in7 ),
    .S(net1),
    .X(\u_skew_usb.d03 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_04.genblk1.u_mux  (.A0(\u_skew_usb.in8 ),
    .A1(\u_skew_usb.in9 ),
    .S(net1),
    .X(\u_skew_usb.d04 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_05.genblk1.u_mux  (.A0(\u_skew_usb.in10 ),
    .A1(\u_skew_usb.in11 ),
    .S(net1),
    .X(\u_skew_usb.d05 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_06.genblk1.u_mux  (.A0(\u_skew_usb.in12 ),
    .A1(\u_skew_usb.in13 ),
    .S(net1),
    .X(\u_skew_usb.d06 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_07.genblk1.u_mux  (.A0(\u_skew_usb.in14 ),
    .A1(\u_skew_usb.in15 ),
    .S(net1),
    .X(\u_skew_usb.d07 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_10.genblk1.u_mux  (.A0(\u_skew_usb.d00 ),
    .A1(\u_skew_usb.d01 ),
    .S(net2),
    .X(\u_skew_usb.d10 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_11.genblk1.u_mux  (.A0(\u_skew_usb.d02 ),
    .A1(\u_skew_usb.d03 ),
    .S(net2),
    .X(\u_skew_usb.d11 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_12.genblk1.u_mux  (.A0(\u_skew_usb.d04 ),
    .A1(\u_skew_usb.d05 ),
    .S(net2),
    .X(\u_skew_usb.d12 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_13.genblk1.u_mux  (.A0(\u_skew_usb.d06 ),
    .A1(\u_skew_usb.d07 ),
    .S(net2),
    .X(\u_skew_usb.d13 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_20.genblk1.u_mux  (.A0(\u_skew_usb.d10 ),
    .A1(\u_skew_usb.d11 ),
    .S(net3),
    .X(\u_skew_usb.d20 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_21.genblk1.u_mux  (.A0(\u_skew_usb.d12 ),
    .A1(\u_skew_usb.d13 ),
    .S(net3),
    .X(\u_skew_usb.d21 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_30.genblk1.u_mux  (.A0(\u_skew_usb.d20 ),
    .A1(\u_skew_usb.d21 ),
    .S(net4),
    .X(\u_skew_usb.d30 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_0.u_buf  (.A(\u_skew_usb.clk_inbuf ),
    .X(\u_skew_usb.in0 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_1.u_buf  (.A(\u_skew_usb.clk_d1 ),
    .X(\u_skew_usb.in1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_10.u_buf  (.A(\u_skew_usb.clk_d10 ),
    .X(\u_skew_usb.in10 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_11.u_buf  (.A(\u_skew_usb.clk_d11 ),
    .X(\u_skew_usb.in11 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_12.u_buf  (.A(\u_skew_usb.clk_d12 ),
    .X(\u_skew_usb.in12 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_13.u_buf  (.A(\u_skew_usb.clk_d13 ),
    .X(\u_skew_usb.in13 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_14.u_buf  (.A(\u_skew_usb.clk_d14 ),
    .X(\u_skew_usb.in14 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_15.u_buf  (.A(\u_skew_usb.clk_d15 ),
    .X(\u_skew_usb.in15 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_2.u_buf  (.A(\u_skew_usb.clk_d2 ),
    .X(\u_skew_usb.in2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_3.u_buf  (.A(\u_skew_usb.clk_d3 ),
    .X(\u_skew_usb.in3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_4.u_buf  (.A(\u_skew_usb.clk_d4 ),
    .X(\u_skew_usb.in4 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_5.u_buf  (.A(\u_skew_usb.clk_d5 ),
    .X(\u_skew_usb.in5 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_6.u_buf  (.A(\u_skew_usb.clk_d6 ),
    .X(\u_skew_usb.in6 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_7.u_buf  (.A(\u_skew_usb.clk_d7 ),
    .X(\u_skew_usb.in7 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_8.u_buf  (.A(\u_skew_usb.clk_d8 ),
    .X(\u_skew_usb.in8 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_9.u_buf  (.A(\u_skew_usb.clk_d9 ),
    .X(\u_skew_usb.in9 ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_async_wb._06_  (.A(\u_usb_host.u_async_wb.PendingRd ),
    .Y(\u_usb_host.u_async_wb._02_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_async_wb._07_  (.A(\u_usb_host.u_async_wb.m_resp_rd_empty ),
    .Y(\u_usb_host.u_async_wb.m_resp_rd_en ));
 sky130_fd_sc_hd__or4b_2 \u_usb_host.u_async_wb._08_  (.A(\u_usb_host.u_async_wb.m_cmd_wr_full ),
    .B(\u_usb_host.u_async_wb.m_cmd_wr_afull ),
    .C(\u_usb_host.u_async_wb.PendingRd ),
    .D_N(\u_usb_host.u_async_wb.wbm_cyc_i ),
    .X(\u_usb_host.u_async_wb._03_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_async_wb._09_  (.A(\u_usb_host.u_async_wb._03_ ),
    .Y(\u_usb_host.u_async_wb.m_cmd_wr_en ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_async_wb._10_  (.A(net43),
    .B(\u_usb_host.u_async_wb._03_ ),
    .Y(\u_usb_host.u_async_wb._00_ ));
 sky130_fd_sc_hd__or3b_1 \u_usb_host.u_async_wb._11_  (.A(net43),
    .B(\u_usb_host.u_async_wb.m_resp_rd_empty ),
    .C_N(\u_usb_host.u_async_wb.wbm_cyc_i ),
    .X(\u_usb_host.u_async_wb._04_ ));
 sky130_fd_sc_hd__a21bo_1 \u_usb_host.u_async_wb._12_  (.A1(net43),
    .A2(\u_usb_host.u_async_wb.m_cmd_wr_en ),
    .B1_N(\u_usb_host.u_async_wb._04_ ),
    .X(net48));
 sky130_fd_sc_hd__o22ai_1 \u_usb_host.u_async_wb._13_  (.A1(net43),
    .A2(\u_usb_host.u_async_wb._03_ ),
    .B1(\u_usb_host.u_async_wb._04_ ),
    .B2(\u_usb_host.u_async_wb._02_ ),
    .Y(\u_usb_host.u_async_wb._01_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._14_  (.A_N(net97),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[36] ),
    .X(\u_usb_host.reg_wr ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._19_  (.A_N(net101),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[4] ),
    .X(\u_usb_host.reg_wdata[0] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._20_  (.A_N(net101),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[5] ),
    .X(\u_usb_host.reg_wdata[1] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._21_  (.A_N(net101),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[6] ),
    .X(\u_usb_host.reg_wdata[2] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._22_  (.A_N(net101),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[7] ),
    .X(\u_usb_host.reg_wdata[3] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._23_  (.A_N(net100),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[8] ),
    .X(\u_usb_host.reg_wdata[4] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._24_  (.A_N(net100),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[9] ),
    .X(\u_usb_host.reg_wdata[5] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._25_  (.A_N(net100),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[10] ),
    .X(\u_usb_host.reg_wdata[6] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._26_  (.A_N(net100),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[11] ),
    .X(\u_usb_host.reg_wdata[7] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._27_  (.A_N(net100),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[12] ),
    .X(\u_usb_host.reg_wdata[8] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._28_  (.A_N(net100),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[13] ),
    .X(\u_usb_host.reg_wdata[9] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._29_  (.A_N(net100),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[14] ),
    .X(\u_usb_host.reg_wdata[10] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._30_  (.A_N(net100),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[15] ),
    .X(\u_usb_host.reg_wdata[11] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._31_  (.A_N(net101),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[16] ),
    .X(\u_usb_host.reg_wdata[12] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._32_  (.A_N(net100),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[17] ),
    .X(\u_usb_host.reg_wdata[13] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._33_  (.A_N(net101),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[18] ),
    .X(\u_usb_host.reg_wdata[14] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._34_  (.A_N(net100),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[19] ),
    .X(\u_usb_host.reg_wdata[15] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._35_  (.A_N(net99),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[20] ),
    .X(\u_usb_host.reg_wdata[16] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._36_  (.A_N(net99),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[21] ),
    .X(\u_usb_host.reg_wdata[17] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._37_  (.A_N(net97),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[22] ),
    .X(\u_usb_host.reg_wdata[18] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._38_  (.A_N(net99),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[23] ),
    .X(\u_usb_host.reg_wdata[19] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._39_  (.A_N(net99),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[24] ),
    .X(\u_usb_host.reg_wdata[20] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._40_  (.A_N(net98),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[25] ),
    .X(\u_usb_host.reg_wdata[21] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._41_  (.A_N(net98),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[26] ),
    .X(\u_usb_host.reg_wdata[22] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._42_  (.A_N(net97),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[27] ),
    .X(\u_usb_host.reg_wdata[23] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._47_  (.A_N(net97),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[32] ),
    .X(\u_usb_host.reg_wdata[28] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._48_  (.A_N(net98),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[33] ),
    .X(\u_usb_host.reg_wdata[29] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._49_  (.A_N(net97),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[34] ),
    .X(\u_usb_host.reg_wdata[30] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._50_  (.A_N(net99),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[35] ),
    .X(\u_usb_host.reg_wdata[31] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._51_  (.A_N(net98),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[37] ),
    .X(\u_usb_host.reg_addr[0] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._52_  (.A_N(net98),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[38] ),
    .X(\u_usb_host.reg_addr[1] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._53_  (.A_N(net97),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[39] ),
    .X(\u_usb_host.reg_addr[2] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._54_  (.A_N(net97),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[40] ),
    .X(\u_usb_host.reg_addr[3] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._55_  (.A_N(net97),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[41] ),
    .X(\u_usb_host.reg_addr[4] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._56_  (.A_N(net97),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[42] ),
    .X(\u_usb_host.reg_addr[5] ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_async_wb._57_  (.A(net97),
    .B(\u_usb_host.u_async_wb.wbs_ack_f ),
    .Y(\u_usb_host.u_async_wb.wbs_cyc_o ));
 sky130_fd_sc_hd__and4bb_1 \u_usb_host.u_async_wb._58_  (.A_N(\u_usb_host.u_async_wb.s_resp_wr_full ),
    .B_N(\u_usb_host.reg_wr ),
    .C(\u_usb_host.u_async_wb.wbs_cyc_o ),
    .D(\u_usb_host.reg_ack ),
    .X(\u_usb_host.u_async_wb.s_resp_wr_en ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb._59_  (.CLK(\u_usb_host.u_async_wb._05_ ),
    .D(\u_usb_host.u_async_wb._00_ ),
    .RESET_B(net260),
    .Q(\u_usb_host.u_async_wb.PendingRd ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb._60_  (.CLK(clknet_4_3_0_usb_clk),
    .D(\u_usb_host.reg_ack ),
    .RESET_B(net292),
    .Q(\u_usb_host.u_async_wb.wbs_ack_f ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_async_wb._61_  (.CLK(clknet_1_1__leaf_app_clk),
    .GATE(\u_usb_host.u_async_wb._01_ ),
    .GCLK(\u_usb_host.u_async_wb._05_ ));
 sky130_fd_sc_hd__clkbuf_1 \u_usb_host.u_async_wb._62_  (.A(\u_usb_host.u_async_wb.wbs_cyc_o ),
    .X(\u_usb_host.reg_cs ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_async_wb.u_cmd_if._041_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[1] ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._000_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_async_wb.u_cmd_if._042_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[0] ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[0] ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_async_wb.u_cmd_if._043_  (.A(net318),
    .Y(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[0] ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_async_wb.u_cmd_if._044_  (.A(net313),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._002_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_async_wb.u_cmd_if._045_  (.A(net318),
    .B(net313),
    .X(\u_usb_host.u_async_wb.u_cmd_if._008_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_async_wb.u_cmd_if._046_  (.A(net318),
    .B(net313),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._009_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_async_wb.u_cmd_if._047_  (.A(\u_usb_host.u_async_wb.u_cmd_if._008_ ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._009_ ),
    .X(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[1] ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_async_wb.u_cmd_if._048_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[1] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[0] ),
    .X(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[1] ));
 sky130_fd_sc_hd__xor2_2 \u_usb_host.u_async_wb.u_cmd_if._049_  (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_1[1] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr[2] ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._010_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_async_wb.u_cmd_if._050_  (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_1[0] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._010_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._011_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_async_wb.u_cmd_if._051_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[0] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._011_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._012_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_async_wb.u_cmd_if._052_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[0] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._011_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._013_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_async_wb.u_cmd_if._053_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[1] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._010_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._014_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_async_wb.u_cmd_if._054_  (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr[2] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[2] ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._015_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_async_wb.u_cmd_if._055_  (.A(\u_usb_host.u_async_wb.u_cmd_if._013_ ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._014_ ),
    .C(\u_usb_host.u_async_wb.u_cmd_if._015_ ),
    .X(\u_usb_host.u_async_wb.m_cmd_wr_full ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_async_wb.u_cmd_if._056_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[1] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[0] ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._016_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_async_wb.u_cmd_if._057_  (.A(\u_usb_host.u_async_wb.u_cmd_if._016_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._017_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_async_wb.u_cmd_if._058_  (.A1(\u_usb_host.u_async_wb.u_cmd_if._013_ ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if._017_ ),
    .B1(\u_usb_host.u_async_wb.u_cmd_if._015_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._018_ ));
 sky130_fd_sc_hd__or3b_1 \u_usb_host.u_async_wb.u_cmd_if._059_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[0] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._011_ ),
    .C_N(\u_usb_host.u_async_wb.u_cmd_if._014_ ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._019_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_async_wb.u_cmd_if._060_  (.A1(\u_usb_host.u_async_wb.u_cmd_if._012_ ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if._014_ ),
    .B1(\u_usb_host.u_async_wb.u_cmd_if._019_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._020_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_async_wb.u_cmd_if._061_  (.A(\u_usb_host.u_async_wb.u_cmd_if._013_ ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._015_ ),
    .C(\u_usb_host.u_async_wb.u_cmd_if._017_ ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._021_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_async_wb.u_cmd_if._062_  (.A(\u_usb_host.u_async_wb.u_cmd_if._018_ ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._020_ ),
    .C(\u_usb_host.u_async_wb.u_cmd_if._021_ ),
    .X(\u_usb_host.u_async_wb.m_cmd_wr_afull ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_async_wb.u_cmd_if._063_  (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_1[1] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr[2] ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._022_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_async_wb.u_cmd_if._064_  (.A(net313),
    .B(\u_usb_host.u_async_wb.u_cmd_if._022_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._023_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_async_wb.u_cmd_if._065_  (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr[2] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[2] ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._024_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_async_wb.u_cmd_if._066_  (.A1(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_1[0] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if._023_ ),
    .B1(\u_usb_host.u_async_wb.u_cmd_if._024_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._025_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_async_wb.u_cmd_if._067_  (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_1[0] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._023_ ),
    .C(\u_usb_host.u_async_wb.u_cmd_if._024_ ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._026_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_async_wb.u_cmd_if._068_  (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_1[0] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._022_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._027_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_async_wb.u_cmd_if._069_  (.A1(net318),
    .A2(\u_usb_host.u_async_wb.u_cmd_if._027_ ),
    .B1(\u_usb_host.u_async_wb.u_cmd_if._023_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._028_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_async_wb.u_cmd_if._070_  (.A1(net318),
    .A2(\u_usb_host.u_async_wb.u_cmd_if._027_ ),
    .B1(\u_usb_host.u_async_wb.u_cmd_if._028_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._029_ ));
 sky130_fd_sc_hd__and3_2 \u_usb_host.u_async_wb.u_cmd_if._071_  (.A(\u_usb_host.u_async_wb.u_cmd_if._025_ ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._026_ ),
    .C(\u_usb_host.u_async_wb.u_cmd_if._029_ ),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_empty ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_async_wb.u_cmd_if._074_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[2] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._016_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[2] ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_async_wb.u_cmd_if._075_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[1] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[2] ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._031_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_async_wb.u_cmd_if._076_  (.A1(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[2] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[1] ),
    .B1(\u_usb_host.u_async_wb.u_cmd_if._031_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._001_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_async_wb.u_cmd_if._077_  (.A(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[2] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._009_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[2] ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_async_wb.u_cmd_if._078_  (.A(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[1] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[2] ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._032_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_async_wb.u_cmd_if._079_  (.A1(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[2] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[1] ),
    .B1(\u_usb_host.u_async_wb.u_cmd_if._032_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._003_ ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._084_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][4] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][4] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][4] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][4] ),
    .S0(net320),
    .S1(net315),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[4] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._085_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][5] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][5] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][5] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][5] ),
    .S0(net320),
    .S1(net315),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[5] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._086_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][6] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][6] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][6] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][6] ),
    .S0(net319),
    .S1(net314),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[6] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._087_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][7] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][7] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][7] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][7] ),
    .S0(net321),
    .S1(net316),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[7] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._088_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][8] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][8] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][8] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][8] ),
    .S0(net320),
    .S1(net316),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[8] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._089_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][9] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][9] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][9] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][9] ),
    .S0(net320),
    .S1(net315),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[9] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._090_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][10] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][10] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][10] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][10] ),
    .S0(net319),
    .S1(net315),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[10] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._091_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][11] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][11] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][11] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][11] ),
    .S0(net321),
    .S1(net316),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[11] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._092_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][12] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][12] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][12] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][12] ),
    .S0(net321),
    .S1(net316),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[12] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._093_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][13] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][13] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][13] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][13] ),
    .S0(net321),
    .S1(net315),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[13] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._094_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][14] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][14] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][14] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][14] ),
    .S0(net320),
    .S1(net315),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[14] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._095_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][15] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][15] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][15] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][15] ),
    .S0(net320),
    .S1(net315),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[15] ));
 sky130_fd_sc_hd__mux4_2 \u_usb_host.u_async_wb.u_cmd_if._096_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][16] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][16] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][16] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][16] ),
    .S0(net319),
    .S1(net314),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[16] ));
 sky130_fd_sc_hd__mux4_2 \u_usb_host.u_async_wb.u_cmd_if._097_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][17] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][17] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][17] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][17] ),
    .S0(net319),
    .S1(net314),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[17] ));
 sky130_fd_sc_hd__mux4_2 \u_usb_host.u_async_wb.u_cmd_if._098_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][18] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][18] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][18] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][18] ),
    .S0(net319),
    .S1(net314),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[18] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._099_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][19] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][19] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][19] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][19] ),
    .S0(net319),
    .S1(net315),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[19] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._100_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][20] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][20] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][20] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][20] ),
    .S0(net319),
    .S1(net314),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[20] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._101_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][21] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][21] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][21] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][21] ),
    .S0(net320),
    .S1(net315),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[21] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._102_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][22] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][22] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][22] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][22] ),
    .S0(net320),
    .S1(net314),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[22] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._103_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][23] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][23] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][23] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][23] ),
    .S0(net319),
    .S1(net314),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[23] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._104_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][24] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][24] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][24] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][24] ),
    .S0(net319),
    .S1(net314),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[24] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._105_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][25] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][25] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][25] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][25] ),
    .S0(net319),
    .S1(net314),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[25] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._106_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][26] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][26] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][26] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][26] ),
    .S0(net317),
    .S1(net312),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[26] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._107_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][27] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][27] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][27] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][27] ),
    .S0(net317),
    .S1(net312),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[27] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._112_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][32] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][32] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][32] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][32] ),
    .S0(net318),
    .S1(net312),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[32] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._113_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][33] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][33] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][33] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][33] ),
    .S0(net318),
    .S1(net313),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[33] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._114_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][34] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][34] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][34] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][34] ),
    .S0(net317),
    .S1(net312),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[34] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._115_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][35] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][35] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][35] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][35] ),
    .S0(net320),
    .S1(net314),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[35] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._116_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][36] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][36] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][36] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][36] ),
    .S0(net317),
    .S1(net312),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[36] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._117_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][37] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][37] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][37] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][37] ),
    .S0(net317),
    .S1(net312),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[37] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._118_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][38] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][38] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][38] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][38] ),
    .S0(net317),
    .S1(net313),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[38] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._119_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][39] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][39] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][39] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][39] ),
    .S0(net317),
    .S1(net312),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[39] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._120_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][40] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][40] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][40] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][40] ),
    .S0(net317),
    .S1(net312),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[40] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._121_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][41] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][41] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][41] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][41] ),
    .S0(net317),
    .S1(net312),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[41] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._122_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][42] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][42] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][42] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][42] ),
    .S0(net317),
    .S1(net312),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[42] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_async_wb.u_cmd_if._123_  (.A(\u_usb_host.u_async_wb.u_cmd_if._000_ ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[0] ),
    .C(\u_usb_host.u_async_wb.m_cmd_wr_en ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._007_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_async_wb.u_cmd_if._124_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[1] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[0] ),
    .C(\u_usb_host.u_async_wb.m_cmd_wr_en ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._005_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_async_wb.u_cmd_if._125_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[1] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[0] ),
    .C(\u_usb_host.u_async_wb.m_cmd_wr_en ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._004_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_async_wb.u_cmd_if._126_  (.A(\u_usb_host.u_async_wb.u_cmd_if._000_ ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[0] ),
    .C(\u_usb_host.u_async_wb.m_cmd_wr_en ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._006_ ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._131_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net15),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._132_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net26),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._133_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net33),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._134_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net36),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._135_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net37),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._136_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net38),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._137_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net39),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._138_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net40),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._139_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net41),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._140_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net42),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._141_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net16),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._142_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net17),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._143_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net18),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._144_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net19),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._145_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net20),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._146_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net21),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._147_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net22),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._148_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net23),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._149_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net24),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._150_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net25),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._151_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net27),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._152_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net28),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._153_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net29),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._154_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net30),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._159_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net31),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._160_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net32),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._161_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net34),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._162_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net35),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._163_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net43),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._164_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net5),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._165_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net6),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._166_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net7),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._167_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net8),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._168_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net9),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._169_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net10),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._174_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net15),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._175_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net26),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._176_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net33),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._177_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net36),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._178_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net37),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._179_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net38),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._180_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net39),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._181_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net40),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._182_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net41),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._183_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net42),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._184_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net16),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._185_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net17),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._186_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net18),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._187_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net19),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._188_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net20),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._189_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net21),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._190_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net22),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._191_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net23),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._192_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net24),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._193_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net25),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._194_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net27),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._195_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net28),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._196_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net29),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._197_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net30),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._202_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net31),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._203_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net32),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._204_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net34),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._205_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net35),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._206_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net43),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._207_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net5),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._208_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net6),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._209_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net7),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._210_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net8),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._211_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net9),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._212_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(net10),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._217_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net15),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._218_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net26),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._219_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net33),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._220_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net36),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._221_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net37),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._222_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net38),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._223_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net39),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._224_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net40),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._225_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net41),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._226_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net42),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._227_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net16),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._228_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net17),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._229_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net18),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._230_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net19),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._231_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net20),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._232_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net21),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._233_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net22),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._234_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net23),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._235_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net24),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._236_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net25),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._237_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net27),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._238_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net28),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._239_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net29),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._240_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net30),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._245_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net31),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][32] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._246_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net32),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][33] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._247_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net34),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][34] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._248_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net35),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][35] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._249_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net43),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][36] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._250_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net5),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][37] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._251_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net6),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][38] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._252_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net7),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][39] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._253_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net8),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][40] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._254_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net9),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][41] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._255_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(net10),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][42] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._260_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net15),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._261_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net26),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._262_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net33),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._263_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net36),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._264_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net37),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._265_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net38),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._266_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net39),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._267_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net40),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._268_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net41),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._269_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net42),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._270_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net16),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._271_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net17),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._272_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net18),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._273_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net19),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._274_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net20),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._275_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net21),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._276_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net22),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._277_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net23),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._278_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net24),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._279_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net25),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._280_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net27),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._281_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net28),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._282_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net29),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._283_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net30),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._288_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net31),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._289_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net32),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._290_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net34),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._291_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net35),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._292_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net43),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._293_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net5),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._294_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net6),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._295_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net7),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._296_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net8),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._297_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net9),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._298_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net10),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][42] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._299_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._033_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[0] ),
    .RESET_B(net263),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._300_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._033_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[1] ),
    .RESET_B(net263),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._301_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._033_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[2] ),
    .RESET_B(net263),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_async_wb.u_cmd_if._302_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._034_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[0] ),
    .RESET_B(net260),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_async_wb.u_cmd_if._303_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._034_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[1] ),
    .RESET_B(net260),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._304_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._034_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[2] ),
    .RESET_B(net261),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._305_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._036_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if._002_ ),
    .RESET_B(net262),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.grey_rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._306_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._036_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if._003_ ),
    .RESET_B(net262),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.grey_rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._307_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._036_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[2] ),
    .RESET_B(net262),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.grey_rd_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._308_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._035_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if._000_ ),
    .RESET_B(net390),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.grey_wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._309_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._035_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if._001_ ),
    .RESET_B(net261),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.grey_wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._310_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._035_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[2] ),
    .RESET_B(net261),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.grey_wr_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._311_  (.CLK(clknet_1_0__leaf_app_clk),
    .D(\u_usb_host.u_async_wb.u_cmd_if.grey_rd_ptr[0] ),
    .RESET_B(net261),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_0[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._312_  (.CLK(clknet_1_0__leaf_app_clk),
    .D(\u_usb_host.u_async_wb.u_cmd_if.grey_rd_ptr[1] ),
    .RESET_B(net261),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_0[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._313_  (.CLK(clknet_1_0__leaf_app_clk),
    .D(\u_usb_host.u_async_wb.u_cmd_if.grey_rd_ptr[2] ),
    .RESET_B(net261),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_0[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._314_  (.CLK(clknet_1_0__leaf_app_clk),
    .D(net485),
    .RESET_B(net261),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._315_  (.CLK(clknet_1_0__leaf_app_clk),
    .D(net467),
    .RESET_B(net261),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._316_  (.CLK(clknet_1_0__leaf_app_clk),
    .D(net477),
    .RESET_B(net261),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._317_  (.CLK(clknet_4_0_0_usb_clk),
    .D(\u_usb_host.u_async_wb.u_cmd_if.grey_wr_ptr[0] ),
    .RESET_B(net262),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_0[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._318_  (.CLK(clknet_4_0_0_usb_clk),
    .D(\u_usb_host.u_async_wb.u_cmd_if.grey_wr_ptr[1] ),
    .RESET_B(net262),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_0[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._319_  (.CLK(clknet_4_0_0_usb_clk),
    .D(\u_usb_host.u_async_wb.u_cmd_if.grey_wr_ptr[2] ),
    .RESET_B(net262),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_0[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._320_  (.CLK(clknet_4_0_0_usb_clk),
    .D(net486),
    .RESET_B(net263),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._321_  (.CLK(clknet_4_0_0_usb_clk),
    .D(net484),
    .RESET_B(net263),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._322_  (.CLK(clknet_4_0_0_usb_clk),
    .D(net488),
    .RESET_B(net263),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr[2] ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_async_wb.u_cmd_if._323_  (.CLK(clknet_4_0_0_usb_clk),
    .GATE(\u_usb_host.reg_ack ),
    .GCLK(\u_usb_host.u_async_wb.u_cmd_if._033_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_async_wb.u_cmd_if._324_  (.CLK(clknet_1_0__leaf_app_clk),
    .GATE(\u_usb_host.u_async_wb.m_cmd_wr_en ),
    .GCLK(\u_usb_host.u_async_wb.u_cmd_if._034_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_async_wb.u_cmd_if._325_  (.CLK(clknet_1_1__leaf_app_clk),
    .GATE(\u_usb_host.u_async_wb.m_cmd_wr_en ),
    .GCLK(\u_usb_host.u_async_wb.u_cmd_if._035_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_async_wb.u_cmd_if._326_  (.CLK(clknet_4_0_0_usb_clk),
    .GATE(\u_usb_host.reg_ack ),
    .GCLK(\u_usb_host.u_async_wb.u_cmd_if._036_ ));
 sky130_fd_sc_hd__dlclkp_4 \u_usb_host.u_async_wb.u_cmd_if._327_  (.CLK(clknet_1_1__leaf_app_clk),
    .GATE(\u_usb_host.u_async_wb.u_cmd_if._004_ ),
    .GCLK(\u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__dlclkp_4 \u_usb_host.u_async_wb.u_cmd_if._328_  (.CLK(clknet_1_1__leaf_app_clk),
    .GATE(\u_usb_host.u_async_wb.u_cmd_if._005_ ),
    .GCLK(\u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__dlclkp_4 \u_usb_host.u_async_wb.u_cmd_if._329_  (.CLK(clknet_1_1__leaf_app_clk),
    .GATE(\u_usb_host.u_async_wb.u_cmd_if._006_ ),
    .GCLK(\u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__dlclkp_4 \u_usb_host.u_async_wb.u_cmd_if._330_  (.CLK(clknet_1_1__leaf_app_clk),
    .GATE(\u_usb_host.u_async_wb.u_cmd_if._007_ ),
    .GCLK(\u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_async_wb.u_resp_if._020_  (.A(\u_usb_host.u_async_wb.u_resp_if.rd_ptr[1] ),
    .Y(\u_usb_host.u_async_wb.u_resp_if._012_ ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_async_wb.u_resp_if._021_  (.A(net311),
    .Y(\u_usb_host.u_async_wb.u_resp_if.rd_ptr_inc[0] ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_async_wb.u_resp_if._022_  (.A(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[0] ),
    .Y(\u_usb_host.u_async_wb.u_resp_if.wr_ptr_inc[0] ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_async_wb.u_resp_if._023_  (.A(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[1] ),
    .Y(\u_usb_host.u_async_wb.u_resp_if._010_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_async_wb.u_resp_if._024_  (.A(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[0] ),
    .B(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[1] ),
    .X(\u_usb_host.u_async_wb.u_resp_if.wr_ptr_inc[1] ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_async_wb.u_resp_if._025_  (.A(\u_usb_host.u_async_wb.u_resp_if.rd_ptr[1] ),
    .B(net311),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_ptr_inc[1] ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_async_wb.u_resp_if._026_  (.A(\u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_1[0] ),
    .B(\u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_1[1] ),
    .Y(\u_usb_host.u_async_wb.u_resp_if._002_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_async_wb.u_resp_if._027_  (.A(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[0] ),
    .B(\u_usb_host.u_async_wb.u_resp_if._002_ ),
    .X(\u_usb_host.u_async_wb.u_resp_if._003_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_async_wb.u_resp_if._028_  (.A(\u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_1[1] ),
    .B(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[1] ),
    .X(\u_usb_host.u_async_wb.u_resp_if._004_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_async_wb.u_resp_if._029_  (.A1(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[0] ),
    .A2(\u_usb_host.u_async_wb.u_resp_if._002_ ),
    .B1(\u_usb_host.u_async_wb.u_resp_if._004_ ),
    .Y(\u_usb_host.u_async_wb.u_resp_if._005_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_async_wb.u_resp_if._030_  (.A(\u_usb_host.u_async_wb.u_resp_if._003_ ),
    .B(\u_usb_host.u_async_wb.u_resp_if._005_ ),
    .Y(\u_usb_host.u_async_wb.s_resp_wr_full ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_async_wb.u_resp_if._032_  (.A(\u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_1[1] ),
    .B(\u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_1[0] ),
    .Y(\u_usb_host.u_async_wb.u_resp_if._006_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_async_wb.u_resp_if._033_  (.A(net311),
    .B(\u_usb_host.u_async_wb.u_resp_if._006_ ),
    .X(\u_usb_host.u_async_wb.u_resp_if._007_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_async_wb.u_resp_if._034_  (.A(\u_usb_host.u_async_wb.u_resp_if.rd_ptr[1] ),
    .B(\u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_1[1] ),
    .Y(\u_usb_host.u_async_wb.u_resp_if._008_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_async_wb.u_resp_if._035_  (.A1(net311),
    .A2(\u_usb_host.u_async_wb.u_resp_if._006_ ),
    .B1(\u_usb_host.u_async_wb.u_resp_if._008_ ),
    .Y(\u_usb_host.u_async_wb.u_resp_if._009_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_async_wb.u_resp_if._036_  (.A(\u_usb_host.u_async_wb.u_resp_if._007_ ),
    .B(\u_usb_host.u_async_wb.u_resp_if._009_ ),
    .Y(\u_usb_host.u_async_wb.m_resp_rd_empty ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._038_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][0] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][0] ),
    .S(net309),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[0] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._039_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][1] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][1] ),
    .S(net309),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[1] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._040_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][2] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][2] ),
    .S(net309),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[2] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._041_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][3] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][3] ),
    .S(net309),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[3] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._042_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][4] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][4] ),
    .S(net387),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[4] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._043_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][5] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][5] ),
    .S(net309),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[5] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._044_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][6] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][6] ),
    .S(net308),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[6] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._045_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][7] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][7] ),
    .S(net309),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[7] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._046_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][8] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][8] ),
    .S(net309),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[8] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._047_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][9] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][9] ),
    .S(net309),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[9] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._048_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][10] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][10] ),
    .S(net387),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[10] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._049_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][11] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][11] ),
    .S(net387),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[11] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._050_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][12] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][12] ),
    .S(net387),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[12] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._051_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][13] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][13] ),
    .S(net387),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[13] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._052_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][14] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][14] ),
    .S(net309),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[14] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._053_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][15] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][15] ),
    .S(net309),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[15] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._054_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][16] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][16] ),
    .S(net307),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[16] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._055_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][17] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][17] ),
    .S(net307),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[17] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._056_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][18] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][18] ),
    .S(net308),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[18] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._057_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][19] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][19] ),
    .S(net308),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[19] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._058_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][20] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][20] ),
    .S(net308),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[20] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._059_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][21] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][21] ),
    .S(net307),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[21] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._060_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][22] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][22] ),
    .S(net308),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[22] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._061_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][23] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][23] ),
    .S(net307),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[23] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._062_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][24] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][24] ),
    .S(net307),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[24] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._063_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][25] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][25] ),
    .S(net308),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[25] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._064_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][26] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][26] ),
    .S(net307),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[26] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._065_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][27] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][27] ),
    .S(net308),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[27] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._066_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][28] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][28] ),
    .S(net307),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[28] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._067_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][29] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][29] ),
    .S(net307),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[29] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._068_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][30] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][30] ),
    .S(net307),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[30] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._069_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][31] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][31] ),
    .S(net307),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[31] ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_async_wb.u_resp_if._071_  (.A(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[0] ),
    .B(\u_usb_host.u_async_wb.s_resp_wr_en ),
    .X(\u_usb_host.u_async_wb.u_resp_if._000_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_async_wb.u_resp_if._072_  (.A(\u_usb_host.u_async_wb.u_resp_if.wr_ptr_inc[0] ),
    .B(\u_usb_host.u_async_wb.s_resp_wr_en ),
    .X(\u_usb_host.u_async_wb.u_resp_if._001_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_async_wb.u_resp_if._073_  (.A(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[0] ),
    .B(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[1] ),
    .X(\u_usb_host.u_async_wb.u_resp_if._011_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_async_wb.u_resp_if._074_  (.A(\u_usb_host.u_async_wb.u_resp_if.rd_ptr[1] ),
    .B(net311),
    .X(\u_usb_host.u_async_wb.u_resp_if._013_ ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._075_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._014_ ),
    .D(\u_usb_host.u_async_wb.u_resp_if.rd_ptr_inc[0] ),
    .RESET_B(net260),
    .Q(\u_usb_host.u_async_wb.u_resp_if.rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_async_wb.u_resp_if._076_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._014_ ),
    .D(\u_usb_host.u_async_wb.u_resp_if.rd_ptr_inc[1] ),
    .RESET_B(net260),
    .Q(\u_usb_host.u_async_wb.u_resp_if.rd_ptr[1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._077_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net424),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._078_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net433),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._079_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net432),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._080_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net419),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._081_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net420),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._082_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net422),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._083_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net430),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._084_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net410),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._085_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net425),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._086_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net404),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._087_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net407),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._088_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net423),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._089_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net414),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._090_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net403),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._091_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net406),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._092_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net415),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._093_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net400),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._094_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net399),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._095_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net418),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._096_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net437),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._097_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net435),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._098_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net416),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._099_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net439),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._100_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net411),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._101_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net401),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._102_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net434),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._103_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net402),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._104_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net431),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._105_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net412),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._106_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net405),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._107_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net421),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._108_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net408),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._110_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net424),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._111_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net433),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._112_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net432),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._113_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net419),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._114_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net420),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._115_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net422),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._116_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net430),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._117_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net410),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._118_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net425),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._119_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net404),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._120_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net407),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._121_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net423),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._122_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net414),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._123_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net403),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._124_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net406),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._125_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net415),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._126_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net400),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._127_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net399),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._128_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net418),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._129_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net437),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._130_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net435),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._131_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net416),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._132_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net439),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._133_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net411),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._134_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net401),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._135_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net434),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._136_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net402),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._137_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net431),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._138_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net412),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._139_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net405),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._140_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net421),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._141_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net408),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][31] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._143_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._016_ ),
    .D(\u_usb_host.u_async_wb.u_resp_if._010_ ),
    .RESET_B(net264),
    .Q(\u_usb_host.u_async_wb.u_resp_if.grey_wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._144_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._016_ ),
    .D(\u_usb_host.u_async_wb.u_resp_if._011_ ),
    .RESET_B(net264),
    .Q(\u_usb_host.u_async_wb.u_resp_if.grey_wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._145_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._017_ ),
    .D(\u_usb_host.u_async_wb.u_resp_if._012_ ),
    .RESET_B(net260),
    .Q(\u_usb_host.u_async_wb.u_resp_if.grey_rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._146_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._017_ ),
    .D(\u_usb_host.u_async_wb.u_resp_if._013_ ),
    .RESET_B(net260),
    .Q(\u_usb_host.u_async_wb.u_resp_if.grey_rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_async_wb.u_resp_if._147_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._015_ ),
    .D(\u_usb_host.u_async_wb.u_resp_if.wr_ptr_inc[0] ),
    .RESET_B(net264),
    .Q(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_async_wb.u_resp_if._148_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._015_ ),
    .D(\u_usb_host.u_async_wb.u_resp_if.wr_ptr_inc[1] ),
    .RESET_B(net264),
    .Q(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._149_  (.CLK(clknet_4_1_0_usb_clk),
    .D(\u_usb_host.u_async_wb.u_resp_if.grey_rd_ptr[0] ),
    .RESET_B(net262),
    .Q(\u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_0[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._150_  (.CLK(clknet_4_1_0_usb_clk),
    .D(\u_usb_host.u_async_wb.u_resp_if.grey_rd_ptr[1] ),
    .RESET_B(net262),
    .Q(\u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_0[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._151_  (.CLK(clknet_4_1_0_usb_clk),
    .D(net468),
    .RESET_B(net262),
    .Q(\u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._152_  (.CLK(clknet_4_1_0_usb_clk),
    .D(net479),
    .RESET_B(net262),
    .Q(\u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._153_  (.CLK(clknet_1_1__leaf_app_clk),
    .D(\u_usb_host.u_async_wb.u_resp_if.grey_wr_ptr[0] ),
    .RESET_B(\u_usb_host.u_async_wb.u_cmd_if.wr_reset_n ),
    .Q(\u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_0[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._154_  (.CLK(clknet_1_1__leaf_app_clk),
    .D(\u_usb_host.u_async_wb.u_resp_if.grey_wr_ptr[1] ),
    .RESET_B(net260),
    .Q(\u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_0[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._155_  (.CLK(clknet_1_1__leaf_app_clk),
    .D(net481),
    .RESET_B(net260),
    .Q(\u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._156_  (.CLK(clknet_1_1__leaf_app_clk),
    .D(net487),
    .RESET_B(net260),
    .Q(\u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_1[1] ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_async_wb.u_resp_if._157_  (.CLK(clknet_1_1__leaf_app_clk),
    .GATE(\u_usb_host.u_async_wb.m_resp_rd_en ),
    .GCLK(\u_usb_host.u_async_wb.u_resp_if._014_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_async_wb.u_resp_if._158_  (.CLK(clknet_4_3_0_usb_clk),
    .GATE(\u_usb_host.u_async_wb.s_resp_wr_en ),
    .GCLK(\u_usb_host.u_async_wb.u_resp_if._015_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_async_wb.u_resp_if._159_  (.CLK(clknet_4_1_0_usb_clk),
    .GATE(\u_usb_host.u_async_wb.s_resp_wr_en ),
    .GCLK(\u_usb_host.u_async_wb.u_resp_if._016_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_async_wb.u_resp_if._160_  (.CLK(clknet_1_1__leaf_app_clk),
    .GATE(\u_usb_host.u_async_wb.m_resp_rd_en ),
    .GCLK(\u_usb_host.u_async_wb.u_resp_if._017_ ));
 sky130_fd_sc_hd__dlclkp_4 \u_usb_host.u_async_wb.u_resp_if._161_  (.CLK(clknet_4_2_0_usb_clk),
    .GATE(\u_usb_host.u_async_wb.u_resp_if._000_ ),
    .GCLK(\u_usb_host.u_async_wb.u_resp_if._018_ ));
 sky130_fd_sc_hd__dlclkp_4 \u_usb_host.u_async_wb.u_resp_if._162_  (.CLK(clknet_4_2_0_usb_clk),
    .GATE(\u_usb_host.u_async_wb.u_resp_if._001_ ),
    .GCLK(\u_usb_host.u_async_wb.u_resp_if._019_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core._203_  (.A(\u_usb_host.u_core.sof_time_q[12] ),
    .Y(\u_usb_host.u_core._061_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core._205_  (.A(net453),
    .Y(\u_usb_host.u_core._002_ ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_core._206_  (.A(\u_usb_host.u_core.sof_time_q[0] ),
    .Y(\u_usb_host.u_core._007_ ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_core._207_  (.A(net449),
    .Y(\u_usb_host.u_core._026_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core._208_  (.A(\u_usb_host.u_core.sof_time_q[2] ),
    .B(\u_usb_host.u_core.sof_time_q[1] ),
    .C(\u_usb_host.u_core.sof_time_q[0] ),
    .X(\u_usb_host.u_core._062_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_core._209_  (.A(\u_usb_host.u_core.sof_time_q[3] ),
    .B(\u_usb_host.u_core.sof_time_q[2] ),
    .C(\u_usb_host.u_core.sof_time_q[1] ),
    .D(\u_usb_host.u_core.sof_time_q[0] ),
    .X(\u_usb_host.u_core._063_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._210_  (.A(\u_usb_host.u_core.sof_time_q[4] ),
    .B(\u_usb_host.u_core._063_ ),
    .X(\u_usb_host.u_core._064_ ));
 sky130_fd_sc_hd__and4b_1 \u_usb_host.u_core._211_  (.A_N(\u_usb_host.u_core.sof_time_q[10] ),
    .B(\u_usb_host.u_core.sof_time_q[11] ),
    .C(\u_usb_host.u_core.sof_time_q[14] ),
    .D(\u_usb_host.u_core.sof_time_q[15] ),
    .X(\u_usb_host.u_core._065_ ));
 sky130_fd_sc_hd__nor4b_1 \u_usb_host.u_core._212_  (.A(\u_usb_host.u_core.sof_time_q[5] ),
    .B(\u_usb_host.u_core.sof_time_q[7] ),
    .C(\u_usb_host.u_core.sof_time_q[8] ),
    .D_N(\u_usb_host.u_core.sof_time_q[6] ),
    .Y(\u_usb_host.u_core._066_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_core._213_  (.A(\u_usb_host.u_core.sof_time_q[9] ),
    .B(\u_usb_host.u_core._061_ ),
    .C(\u_usb_host.u_core.sof_time_q[13] ),
    .D(\u_usb_host.u_core._066_ ),
    .X(\u_usb_host.u_core._067_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core._214_  (.A(\u_usb_host.u_core._064_ ),
    .B(\u_usb_host.u_core._065_ ),
    .C(\u_usb_host.u_core._067_ ),
    .X(\u_usb_host.u_core._068_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core._215_  (.A(\u_usb_host.u_core.usb_ctrl_enable_sof_out_w ),
    .B(net372),
    .C(\u_usb_host.u_core._068_ ),
    .X(\u_usb_host.u_core.send_sof_w ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._215__372  (.HI(net372));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_core._216_  (.A1(\u_usb_host.u_core.sof_time_q[1] ),
    .A2(\u_usb_host.u_core.sof_time_q[0] ),
    .B1(\u_usb_host.u_core.sof_time_q[2] ),
    .X(\u_usb_host.u_core._069_ ));
 sky130_fd_sc_hd__o311a_1 \u_usb_host.u_core._217_  (.A1(\u_usb_host.u_core.sof_time_q[3] ),
    .A2(\u_usb_host.u_core.sof_time_q[4] ),
    .A3(\u_usb_host.u_core._069_ ),
    .B1(\u_usb_host.u_core.sof_time_q[6] ),
    .C1(\u_usb_host.u_core.sof_time_q[5] ),
    .X(\u_usb_host.u_core._070_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_core._218_  (.A(\u_usb_host.u_core.sof_time_q[13] ),
    .B(\u_usb_host.u_core.sof_time_q[14] ),
    .C(\u_usb_host.u_core.sof_time_q[15] ),
    .X(\u_usb_host.u_core._071_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core._219_  (.A(\u_usb_host.u_core.sof_time_q[9] ),
    .B(\u_usb_host.u_core.sof_time_q[10] ),
    .C(\u_usb_host.u_core.sof_time_q[11] ),
    .D(\u_usb_host.u_core.sof_time_q[12] ),
    .X(\u_usb_host.u_core._072_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core._220_  (.A(\u_usb_host.u_core.sof_time_q[7] ),
    .B(\u_usb_host.u_core.sof_time_q[8] ),
    .C(\u_usb_host.u_core._071_ ),
    .D(\u_usb_host.u_core._072_ ),
    .X(\u_usb_host.u_core._073_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._221_  (.A(\u_usb_host.u_core._070_ ),
    .B(\u_usb_host.u_core._073_ ),
    .Y(\u_usb_host.u_core._074_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core._222_  (.A(\u_usb_host.u_core.sof_time_q[10] ),
    .B(\u_usb_host.u_core.sof_time_q[11] ),
    .C(\u_usb_host.u_core.sof_time_q[12] ),
    .X(\u_usb_host.u_core._075_ ));
 sky130_fd_sc_hd__o211a_1 \u_usb_host.u_core._223_  (.A1(\u_usb_host.u_core.sof_time_q[13] ),
    .A2(\u_usb_host.u_core._075_ ),
    .B1(\u_usb_host.u_core.sof_time_q[15] ),
    .C1(\u_usb_host.u_core.sof_time_q[14] ),
    .X(\u_usb_host.u_core._076_ ));
 sky130_fd_sc_hd__o31a_1 \u_usb_host.u_core._224_  (.A1(\u_usb_host.u_core.sof_time_q[2] ),
    .A2(\u_usb_host.u_core.sof_time_q[1] ),
    .A3(\u_usb_host.u_core.sof_time_q[0] ),
    .B1(\u_usb_host.u_core.sof_time_q[4] ),
    .X(\u_usb_host.u_core._077_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core._225_  (.A1(\u_usb_host.u_core.sof_time_q[3] ),
    .A2(\u_usb_host.u_core.sof_time_q[5] ),
    .A3(\u_usb_host.u_core._077_ ),
    .B1(\u_usb_host.u_core.sof_time_q[6] ),
    .X(\u_usb_host.u_core._078_ ));
 sky130_fd_sc_hd__and4b_1 \u_usb_host.u_core._226_  (.A_N(\u_usb_host.u_core.sof_time_q[13] ),
    .B(\u_usb_host.u_core.sof_time_q[9] ),
    .C(\u_usb_host.u_core.sof_time_q[8] ),
    .D(\u_usb_host.u_core.sof_time_q[7] ),
    .X(\u_usb_host.u_core._079_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_core._227_  (.A(\u_usb_host.u_core.sof_time_q[12] ),
    .B(\u_usb_host.u_core._065_ ),
    .C(\u_usb_host.u_core._078_ ),
    .D(\u_usb_host.u_core._079_ ),
    .X(\u_usb_host.u_core._080_ ));
 sky130_fd_sc_hd__o31ai_1 \u_usb_host.u_core._228_  (.A1(\u_usb_host.u_core._074_ ),
    .A2(\u_usb_host.u_core._076_ ),
    .A3(\u_usb_host.u_core._080_ ),
    .B1(\u_usb_host.u_core.usb_ctrl_enable_sof_out_w ),
    .Y(\u_usb_host.u_core._081_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core._229_  (.A1(net373),
    .A2(\u_usb_host.u_core.usb_rx_stat_start_pend_in_w ),
    .A3(\u_usb_host.u_core._081_ ),
    .B1(\u_usb_host.u_core.transfer_start_q ),
    .X(\u_usb_host.u_core._038_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._229__373  (.HI(net373));
 sky130_fd_sc_hd__nand2b_1 \u_usb_host.u_core._230_  (.A_N(\u_usb_host.reg_addr[5] ),
    .B(\u_usb_host.reg_addr[4] ),
    .Y(\u_usb_host.u_core._082_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core._231_  (.A(\u_usb_host.u_core._082_ ),
    .Y(\u_usb_host.u_core._083_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._232_  (.A(\u_usb_host.reg_addr[1] ),
    .B(\u_usb_host.reg_addr[0] ),
    .Y(\u_usb_host.u_core._084_ ));
 sky130_fd_sc_hd__and3b_1 \u_usb_host.u_core._233_  (.A_N(\u_usb_host.reg_addr[2] ),
    .B(\u_usb_host.reg_addr[3] ),
    .C(\u_usb_host.u_core._084_ ),
    .X(\u_usb_host.u_core._085_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._234_  (.A(\u_usb_host.u_core._083_ ),
    .B(\u_usb_host.u_core._085_ ),
    .X(\u_usb_host.u_core._086_ ));
 sky130_fd_sc_hd__and3_2 \u_usb_host.u_core._235_  (.A(\u_usb_host.u_core.cfg_wr ),
    .B(\u_usb_host.u_core._083_ ),
    .C(\u_usb_host.u_core._085_ ),
    .X(\u_usb_host.u_core._037_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._236_  (.A(\u_usb_host.u_core.fifo_flush_q ),
    .B(\u_usb_host.u_core._037_ ),
    .X(\u_usb_host.u_core._036_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._237_  (.A(\u_usb_host.u_core.u_sie.utmi_linestate_i[1] ),
    .B(\u_usb_host.u_core.u_sie.utmi_linestate_i[0] ),
    .X(\u_usb_host.u_core._000_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._238_  (.A(\u_usb_host.u_core.usb_irq_ack_device_detect_out_w ),
    .B(\u_usb_host.u_core._000_ ),
    .X(\u_usb_host.u_core._045_ ));
 sky130_fd_sc_hd__or2_2 \u_usb_host.u_core._239_  (.A(net349),
    .B(net352),
    .X(\u_usb_host.u_core._001_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._239__349  (.LO(net349));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._239__352  (.LO(net352));
 sky130_fd_sc_hd__and2b_2 \u_usb_host.u_core._240_  (.A_N(\u_usb_host.u_core.err_cond_q ),
    .B(\u_usb_host.u_core._001_ ),
    .X(\u_usb_host.u_core._004_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._241_  (.A(\u_usb_host.u_core.usb_irq_ack_err_out_w ),
    .B(\u_usb_host.u_core._004_ ),
    .X(\u_usb_host.u_core._044_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._242_  (.A(\u_usb_host.u_core.sof_irq_q ),
    .B(\u_usb_host.u_core.usb_irq_ack_sof_out_w ),
    .X(\u_usb_host.u_core._043_ ));
 sky130_fd_sc_hd__or2_2 \u_usb_host.u_core._243_  (.A(net354),
    .B(net351),
    .X(\u_usb_host.u_core._003_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._243__351  (.LO(net351));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._243__354  (.LO(net354));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._244_  (.A(\u_usb_host.u_core.usb_irq_ack_done_out_w ),
    .B(\u_usb_host.u_core._003_ ),
    .X(\u_usb_host.u_core._042_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._245_  (.A(\u_usb_host.u_core.usb_ctrl_wr_q ),
    .B(\u_usb_host.u_core.utmi_rxerror_i ),
    .X(\u_usb_host.u_core._041_ ));
 sky130_fd_sc_hd__a21bo_1 \u_usb_host.u_core._246_  (.A1(\u_usb_host.u_core.usb_ctrl_enable_sof_out_w ),
    .A2(net374),
    .B1_N(\u_usb_host.u_core._068_ ),
    .X(\u_usb_host.u_core._040_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._246__374  (.HI(net374));
 sky130_fd_sc_hd__nand3_2 \u_usb_host.u_core._247_  (.A(net451),
    .B(net375),
    .C(\u_usb_host.u_core._068_ ),
    .Y(\u_usb_host.u_core._087_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._247__375  (.HI(net375));
 sky130_fd_sc_hd__a31oi_1 \u_usb_host.u_core._248_  (.A1(net376),
    .A2(\u_usb_host.u_core.usb_rx_stat_start_pend_in_w ),
    .A3(\u_usb_host.u_core._081_ ),
    .B1(\u_usb_host.u_core.send_sof_w ),
    .Y(\u_usb_host.u_core._088_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._248__376  (.HI(net376));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_core._250_  (.A_N(\u_usb_host.reg_ack ),
    .B(\u_usb_host.reg_cs ),
    .X(\u_usb_host.u_core._006_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._251_  (.A(\u_usb_host.reg_wr ),
    .B(\u_usb_host.u_core._006_ ),
    .X(\u_usb_host.u_core._047_ ));
 sky130_fd_sc_hd__or4_4 \u_usb_host.u_core._252_  (.A(\u_usb_host.reg_addr[1] ),
    .B(\u_usb_host.reg_addr[0] ),
    .C(\u_usb_host.reg_addr[2] ),
    .D(\u_usb_host.reg_addr[3] ),
    .X(\u_usb_host.u_core._089_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._253_  (.A(\u_usb_host.reg_addr[5] ),
    .B(\u_usb_host.reg_addr[4] ),
    .Y(\u_usb_host.u_core._090_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._254_  (.A(\u_usb_host.reg_addr[5] ),
    .B(\u_usb_host.reg_addr[4] ),
    .X(\u_usb_host.u_core._091_ ));
 sky130_fd_sc_hd__nor2_4 \u_usb_host.u_core._255_  (.A(\u_usb_host.u_core._089_ ),
    .B(\u_usb_host.u_core._091_ ),
    .Y(\u_usb_host.u_core._092_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core._256_  (.A(\u_usb_host.u_core.cfg_wr ),
    .B(\u_usb_host.u_core._092_ ),
    .X(\u_usb_host.u_core._025_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core._257_  (.A(\u_usb_host.u_core._082_ ),
    .B(\u_usb_host.u_core._089_ ),
    .Y(\u_usb_host.u_core._093_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._258_  (.A(\u_usb_host.u_core.cfg_wr ),
    .B(\u_usb_host.u_core._093_ ),
    .X(\u_usb_host.u_core._034_ ));
 sky130_fd_sc_hd__or4b_1 \u_usb_host.u_core._259_  (.A(\u_usb_host.reg_addr[1] ),
    .B(\u_usb_host.reg_addr[0] ),
    .C(\u_usb_host.reg_addr[3] ),
    .D_N(\u_usb_host.reg_addr[2] ),
    .X(\u_usb_host.u_core._094_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core._260_  (.A(\u_usb_host.u_core._082_ ),
    .B(\u_usb_host.u_core._094_ ),
    .Y(\u_usb_host.u_core._095_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._261_  (.A(\u_usb_host.u_core.cfg_wr ),
    .B(net95),
    .X(\u_usb_host.u_core._035_ ));
 sky130_fd_sc_hd__nor3b_4 \u_usb_host.u_core._262_  (.A(\u_usb_host.reg_addr[4] ),
    .B(\u_usb_host.u_core._089_ ),
    .C_N(\u_usb_host.reg_addr[5] ),
    .Y(\u_usb_host.u_core._096_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core._264_  (.A(\u_usb_host.u_core.sof_time_q[1] ),
    .B(\u_usb_host.u_core.sof_time_q[0] ),
    .X(\u_usb_host.u_core._014_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_core._265_  (.A1(\u_usb_host.u_core.sof_time_q[1] ),
    .A2(\u_usb_host.u_core.sof_time_q[0] ),
    .B1(\u_usb_host.u_core.sof_time_q[2] ),
    .Y(\u_usb_host.u_core._097_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._266_  (.A(\u_usb_host.u_core._062_ ),
    .B(\u_usb_host.u_core._097_ ),
    .Y(\u_usb_host.u_core._015_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._267_  (.A(\u_usb_host.u_core.sof_time_q[3] ),
    .B(\u_usb_host.u_core._062_ ),
    .Y(\u_usb_host.u_core._098_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._268_  (.A(\u_usb_host.u_core._063_ ),
    .B(\u_usb_host.u_core._098_ ),
    .Y(\u_usb_host.u_core._016_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._269_  (.A(\u_usb_host.u_core.sof_time_q[4] ),
    .B(\u_usb_host.u_core._063_ ),
    .Y(\u_usb_host.u_core._099_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._270_  (.A(\u_usb_host.u_core._064_ ),
    .B(\u_usb_host.u_core._099_ ),
    .Y(\u_usb_host.u_core._017_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core._271_  (.A1(\u_usb_host.u_core.sof_time_q[5] ),
    .A2(\u_usb_host.u_core._064_ ),
    .B1(\u_usb_host.u_core._087_ ),
    .Y(\u_usb_host.u_core._100_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_core._272_  (.A1(\u_usb_host.u_core.sof_time_q[5] ),
    .A2(\u_usb_host.u_core._064_ ),
    .B1(\u_usb_host.u_core._100_ ),
    .Y(\u_usb_host.u_core._018_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_core._273_  (.A(\u_usb_host.u_core.sof_time_q[5] ),
    .B(\u_usb_host.u_core.sof_time_q[4] ),
    .C(\u_usb_host.u_core.sof_time_q[6] ),
    .D(\u_usb_host.u_core._063_ ),
    .X(\u_usb_host.u_core._101_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_core._274_  (.A1(\u_usb_host.u_core.sof_time_q[5] ),
    .A2(\u_usb_host.u_core._064_ ),
    .B1(\u_usb_host.u_core.sof_time_q[6] ),
    .Y(\u_usb_host.u_core._102_ ));
 sky130_fd_sc_hd__nor3_1 \u_usb_host.u_core._275_  (.A(\u_usb_host.u_core.send_sof_w ),
    .B(\u_usb_host.u_core._101_ ),
    .C(\u_usb_host.u_core._102_ ),
    .Y(\u_usb_host.u_core._019_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core._276_  (.A(\u_usb_host.u_core.sof_time_q[7] ),
    .B(\u_usb_host.u_core._101_ ),
    .Y(\u_usb_host.u_core._103_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core._277_  (.A(\u_usb_host.u_core.sof_time_q[7] ),
    .B(\u_usb_host.u_core._101_ ),
    .X(\u_usb_host.u_core._020_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core._278_  (.A(\u_usb_host.u_core.sof_time_q[8] ),
    .B(\u_usb_host.u_core._103_ ),
    .Y(\u_usb_host.u_core._021_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core._279_  (.A1(\u_usb_host.u_core.sof_time_q[7] ),
    .A2(\u_usb_host.u_core.sof_time_q[8] ),
    .A3(\u_usb_host.u_core._101_ ),
    .B1(\u_usb_host.u_core.sof_time_q[9] ),
    .X(\u_usb_host.u_core._104_ ));
 sky130_fd_sc_hd__and4_2 \u_usb_host.u_core._280_  (.A(\u_usb_host.u_core.sof_time_q[7] ),
    .B(\u_usb_host.u_core.sof_time_q[8] ),
    .C(\u_usb_host.u_core.sof_time_q[9] ),
    .D(\u_usb_host.u_core._101_ ),
    .X(\u_usb_host.u_core._105_ ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_core._281_  (.A(\u_usb_host.u_core._105_ ),
    .Y(\u_usb_host.u_core._106_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core._282_  (.A(\u_usb_host.u_core._087_ ),
    .B(\u_usb_host.u_core._104_ ),
    .C(\u_usb_host.u_core._106_ ),
    .X(\u_usb_host.u_core._022_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._283_  (.A(\u_usb_host.u_core.sof_time_q[10] ),
    .B(\u_usb_host.u_core._105_ ),
    .X(\u_usb_host.u_core._107_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._284_  (.A(\u_usb_host.u_core.sof_time_q[10] ),
    .B(\u_usb_host.u_core._105_ ),
    .Y(\u_usb_host.u_core._108_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._285_  (.A(\u_usb_host.u_core._107_ ),
    .B(\u_usb_host.u_core._108_ ),
    .Y(\u_usb_host.u_core._008_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core._286_  (.A(\u_usb_host.u_core.sof_time_q[11] ),
    .B(\u_usb_host.u_core._107_ ),
    .Y(\u_usb_host.u_core._109_ ));
 sky130_fd_sc_hd__o211a_1 \u_usb_host.u_core._287_  (.A1(\u_usb_host.u_core.sof_time_q[11] ),
    .A2(\u_usb_host.u_core._107_ ),
    .B1(\u_usb_host.u_core._109_ ),
    .C1(\u_usb_host.u_core._087_ ),
    .X(\u_usb_host.u_core._009_ ));
 sky130_fd_sc_hd__a22oi_1 \u_usb_host.u_core._288_  (.A1(\u_usb_host.u_core._075_ ),
    .A2(\u_usb_host.u_core._105_ ),
    .B1(\u_usb_host.u_core._109_ ),
    .B2(\u_usb_host.u_core._061_ ),
    .Y(\u_usb_host.u_core._010_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._289_  (.A1(\u_usb_host.u_core._075_ ),
    .A2(\u_usb_host.u_core._105_ ),
    .B1(\u_usb_host.u_core.sof_time_q[13] ),
    .X(\u_usb_host.u_core._110_ ));
 sky130_fd_sc_hd__nand3_1 \u_usb_host.u_core._290_  (.A(\u_usb_host.u_core.sof_time_q[13] ),
    .B(\u_usb_host.u_core._075_ ),
    .C(\u_usb_host.u_core._105_ ),
    .Y(\u_usb_host.u_core._111_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core._291_  (.A(\u_usb_host.u_core._087_ ),
    .B(\u_usb_host.u_core._110_ ),
    .C(\u_usb_host.u_core._111_ ),
    .X(\u_usb_host.u_core._011_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core._292_  (.A1(\u_usb_host.u_core.sof_time_q[13] ),
    .A2(\u_usb_host.u_core._075_ ),
    .A3(\u_usb_host.u_core._105_ ),
    .B1(\u_usb_host.u_core.sof_time_q[14] ),
    .X(\u_usb_host.u_core._112_ ));
 sky130_fd_sc_hd__nand4_1 \u_usb_host.u_core._293_  (.A(\u_usb_host.u_core.sof_time_q[13] ),
    .B(\u_usb_host.u_core.sof_time_q[14] ),
    .C(\u_usb_host.u_core._075_ ),
    .D(\u_usb_host.u_core._105_ ),
    .Y(\u_usb_host.u_core._113_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core._294_  (.A(\u_usb_host.u_core._087_ ),
    .B(\u_usb_host.u_core._112_ ),
    .C(\u_usb_host.u_core._113_ ),
    .X(\u_usb_host.u_core._012_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core._295_  (.A(\u_usb_host.u_core.sof_time_q[15] ),
    .B(\u_usb_host.u_core._113_ ),
    .Y(\u_usb_host.u_core._114_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._296_  (.A(\u_usb_host.u_core._087_ ),
    .B(\u_usb_host.u_core._114_ ),
    .X(\u_usb_host.u_core._013_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._297_  (.A(\u_usb_host.u_core._002_ ),
    .B(net368),
    .X(\u_usb_host.u_core._115_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._297__368  (.LO(net368));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core._298_  (.A1(\u_usb_host.u_core.transfer_start_q ),
    .A2(\u_usb_host.u_core._088_ ),
    .B1(\u_usb_host.u_core._115_ ),
    .Y(\u_usb_host.u_core._023_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._301_  (.A(\u_usb_host.u_core._091_ ),
    .B(\u_usb_host.u_core._094_ ),
    .Y(\u_usb_host.u_core._116_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._302_  (.A(\u_usb_host.u_core.sof_time_q[8] ),
    .B(net92),
    .X(\u_usb_host.u_core.reg_rdata_r[24] ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._303_  (.A(\u_usb_host.u_core.sof_time_q[9] ),
    .B(net93),
    .X(\u_usb_host.u_core.reg_rdata_r[25] ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._304_  (.A(\u_usb_host.u_core.sof_time_q[10] ),
    .B(net93),
    .X(\u_usb_host.u_core.reg_rdata_r[26] ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._305_  (.A(\u_usb_host.u_core.sof_time_q[11] ),
    .B(net93),
    .X(\u_usb_host.u_core.reg_rdata_r[27] ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_core._325_  (.A(\u_usb_host.reg_addr[2] ),
    .B(\u_usb_host.reg_addr[3] ),
    .C(\u_usb_host.u_core._083_ ),
    .D(\u_usb_host.u_core._084_ ),
    .X(\u_usb_host.u_core._117_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._326_  (.A1(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[0] ),
    .A2(net89),
    .B1(net92),
    .B2(\u_usb_host.u_core.sof_time_q[0] ),
    .X(\u_usb_host.u_core._118_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._327_  (.A1(net325),
    .A2(net86),
    .B1(\u_usb_host.u_core._118_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[16] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._327__325  (.LO(net325));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._328_  (.A1(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[1] ),
    .A2(net89),
    .B1(net92),
    .B2(\u_usb_host.u_core.sof_time_q[1] ),
    .X(\u_usb_host.u_core._119_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._329_  (.A1(net326),
    .A2(net86),
    .B1(\u_usb_host.u_core._119_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[17] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._329__326  (.LO(net326));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._330_  (.A1(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[2] ),
    .A2(net89),
    .B1(net92),
    .B2(\u_usb_host.u_core.sof_time_q[2] ),
    .X(\u_usb_host.u_core._120_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._331_  (.A1(net327),
    .A2(net86),
    .B1(\u_usb_host.u_core._120_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[18] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._331__327  (.LO(net327));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._332_  (.A(\u_usb_host.u_core.sof_time_q[3] ),
    .B(net92),
    .X(\u_usb_host.u_core._121_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core._333_  (.A1(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[3] ),
    .A2(net89),
    .B1(net86),
    .B2(net328),
    .C1(\u_usb_host.u_core._121_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[19] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._333__328  (.LO(net328));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._334_  (.A(\u_usb_host.u_core.sof_time_q[4] ),
    .B(net92),
    .X(\u_usb_host.u_core._122_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core._335_  (.A1(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[4] ),
    .A2(net89),
    .B1(net86),
    .B2(net329),
    .C1(\u_usb_host.u_core._122_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[20] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._335__329  (.LO(net329));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._336_  (.A1(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[5] ),
    .A2(net89),
    .B1(net92),
    .B2(\u_usb_host.u_core.sof_time_q[5] ),
    .X(\u_usb_host.u_core._123_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._337_  (.A1(net330),
    .A2(net86),
    .B1(\u_usb_host.u_core._123_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[21] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._337__330  (.LO(net330));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._338_  (.A1(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[6] ),
    .A2(net89),
    .B1(net92),
    .B2(\u_usb_host.u_core.sof_time_q[6] ),
    .X(\u_usb_host.u_core._124_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._339_  (.A1(net331),
    .A2(net86),
    .B1(\u_usb_host.u_core._124_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[22] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._339__331  (.LO(net331));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._340_  (.A1(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[7] ),
    .A2(net89),
    .B1(net92),
    .B2(\u_usb_host.u_core.sof_time_q[7] ),
    .X(\u_usb_host.u_core._125_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._341_  (.A1(net332),
    .A2(net86),
    .B1(\u_usb_host.u_core._125_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[23] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._341__332  (.LO(net332));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._342_  (.A1(\u_usb_host.u_core.utmi_xcvrselect_o[1] ),
    .A2(\u_usb_host.u_core._092_ ),
    .B1(\u_usb_host.u_core._096_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.data_o[4] ),
    .X(\u_usb_host.u_core._126_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._343_  (.A1(\u_usb_host.u_core.u_sie.data_len_i[4] ),
    .A2(net96),
    .B1(net87),
    .B2(net337),
    .X(\u_usb_host.u_core._127_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._343__337  (.LO(net337));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._344_  (.A(\u_usb_host.u_core._126_ ),
    .B(\u_usb_host.u_core._127_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[4] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._345_  (.A1(\u_usb_host.u_core.sof_time_q[15] ),
    .A2(net93),
    .B1(net86),
    .B2(net392),
    .X(\u_usb_host.u_core.reg_rdata_r[31] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._346_  (.A1(\u_usb_host.u_core.usb_ctrl_enable_sof_out_w ),
    .A2(\u_usb_host.u_core._092_ ),
    .B1(net94),
    .B2(\u_usb_host.u_core.u_sie.utmi_linestate_i[0] ),
    .X(\u_usb_host.u_core._128_ ));
 sky130_fd_sc_hd__and4_2 \u_usb_host.u_core._347_  (.A(\u_usb_host.reg_addr[2] ),
    .B(\u_usb_host.reg_addr[3] ),
    .C(\u_usb_host.u_core._084_ ),
    .D(\u_usb_host.u_core._090_ ),
    .X(\u_usb_host.u_core._129_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._348_  (.A1(\u_usb_host.u_core.usb_irq_mask_sof_out_w ),
    .A2(\u_usb_host.u_core._093_ ),
    .B1(net95),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[0] ),
    .X(\u_usb_host.u_core._130_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core._349_  (.A1(net333),
    .A2(net88),
    .B1(\u_usb_host.u_core._129_ ),
    .B2(net426),
    .C1(\u_usb_host.u_core._130_ ),
    .X(\u_usb_host.u_core._131_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._349__333  (.LO(net333));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core._350_  (.A1(\u_usb_host.u_core.u_fifo_rx.data_o[0] ),
    .A2(\u_usb_host.u_core._096_ ),
    .B1(\u_usb_host.u_core._128_ ),
    .C1(net427),
    .X(\u_usb_host.u_core.reg_rdata_r[0] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._351_  (.A1(net409),
    .A2(\u_usb_host.u_core._092_ ),
    .B1(net95),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[6] ),
    .X(\u_usb_host.u_core._132_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._352_  (.A1(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[1] ),
    .A2(net90),
    .B1(net88),
    .B2(net339),
    .X(\u_usb_host.u_core._133_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._352__339  (.LO(net339));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core._353_  (.A1(\u_usb_host.u_core.u_fifo_rx.data_o[6] ),
    .A2(\u_usb_host.u_core._096_ ),
    .B1(\u_usb_host.u_core._132_ ),
    .C1(\u_usb_host.u_core._133_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[6] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._354_  (.A1(\u_usb_host.u_core.utmi_xcvrselect_o[0] ),
    .A2(\u_usb_host.u_core._092_ ),
    .B1(net95),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[3] ),
    .X(\u_usb_host.u_core._134_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._355_  (.A1(net413),
    .A2(\u_usb_host.u_core._093_ ),
    .B1(\u_usb_host.u_core._096_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.data_o[3] ),
    .X(\u_usb_host.u_core._135_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core._356_  (.A1(net336),
    .A2(net87),
    .B1(\u_usb_host.u_core._134_ ),
    .C1(\u_usb_host.u_core._135_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[3] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._356__336  (.LO(net336));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._357_  (.A1(net396),
    .A2(\u_usb_host.u_core._092_ ),
    .B1(net95),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[5] ),
    .X(\u_usb_host.u_core._136_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._358_  (.A1(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[0] ),
    .A2(net91),
    .B1(net87),
    .B2(net338),
    .X(\u_usb_host.u_core._137_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._358__338  (.LO(net338));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core._359_  (.A1(\u_usb_host.u_core.u_fifo_rx.data_o[5] ),
    .A2(\u_usb_host.u_core._096_ ),
    .B1(\u_usb_host.u_core._136_ ),
    .C1(\u_usb_host.u_core._137_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[5] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._360_  (.A1(\u_usb_host.u_core.u_sie.data_len_i[2] ),
    .A2(net95),
    .B1(net94),
    .B2(\u_usb_host.u_core.usb_err_q ),
    .X(\u_usb_host.u_core._138_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._361_  (.A1(net335),
    .A2(net88),
    .B1(\u_usb_host.u_core._129_ ),
    .B2(\u_usb_host.u_core.intr_err_q ),
    .X(\u_usb_host.u_core._139_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._361__335  (.LO(net335));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core._362_  (.A1(\u_usb_host.u_core.utmi_op_mode_o[1] ),
    .A2(\u_usb_host.u_core._092_ ),
    .B1(\u_usb_host.u_core._093_ ),
    .B2(net393),
    .C1(\u_usb_host.u_core._139_ ),
    .X(\u_usb_host.u_core._140_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core._363_  (.A1(\u_usb_host.u_core.u_fifo_rx.data_o[2] ),
    .A2(\u_usb_host.u_core._096_ ),
    .B1(\u_usb_host.u_core._138_ ),
    .C1(net394),
    .X(\u_usb_host.u_core.reg_rdata_r[2] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._364_  (.A1(net429),
    .A2(\u_usb_host.u_core._092_ ),
    .B1(net95),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[7] ),
    .X(\u_usb_host.u_core._141_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._365_  (.A1(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[2] ),
    .A2(net90),
    .B1(net88),
    .B2(net340),
    .X(\u_usb_host.u_core._142_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._365__340  (.LO(net340));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core._366_  (.A1(\u_usb_host.u_core.u_fifo_rx.data_o[7] ),
    .A2(\u_usb_host.u_core._096_ ),
    .B1(\u_usb_host.u_core._141_ ),
    .C1(\u_usb_host.u_core._142_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[7] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._367_  (.A1(\u_usb_host.u_core.usb_irq_mask_done_out_w ),
    .A2(\u_usb_host.u_core._093_ ),
    .B1(net96),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[1] ),
    .X(\u_usb_host.u_core._143_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._368_  (.A1(\u_usb_host.u_core.utmi_op_mode_o[0] ),
    .A2(\u_usb_host.u_core._092_ ),
    .B1(net94),
    .B2(\u_usb_host.u_core.u_sie.utmi_linestate_i[1] ),
    .X(\u_usb_host.u_core._144_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core._369_  (.A1(net334),
    .A2(net87),
    .B1(\u_usb_host.u_core._129_ ),
    .B2(net397),
    .C1(\u_usb_host.u_core._144_ ),
    .X(\u_usb_host.u_core._145_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._369__334  (.LO(net334));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core._370_  (.A1(\u_usb_host.u_core.u_fifo_rx.data_o[1] ),
    .A2(\u_usb_host.u_core._096_ ),
    .B1(\u_usb_host.u_core._143_ ),
    .C1(\u_usb_host.u_core._145_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[1] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._371_  (.A1(net450),
    .A2(net89),
    .B1(net93),
    .B2(\u_usb_host.u_core.sof_time_q[14] ),
    .X(\u_usb_host.u_core._146_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._372_  (.A1(net353),
    .A2(net86),
    .B1(\u_usb_host.u_core._146_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[30] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._372__353  (.LO(net353));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._373_  (.A1(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[3] ),
    .A2(net90),
    .B1(net95),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[8] ),
    .X(\u_usb_host.u_core._147_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._374_  (.A1(net341),
    .A2(net88),
    .B1(\u_usb_host.u_core._147_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[8] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._374__341  (.LO(net341));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._375_  (.A1(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[0] ),
    .A2(net90),
    .B1(net96),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[9] ),
    .X(\u_usb_host.u_core._148_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._376_  (.A1(net342),
    .A2(net87),
    .B1(\u_usb_host.u_core._148_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[9] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._376__342  (.LO(net342));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._377_  (.A1(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[1] ),
    .A2(net90),
    .B1(net96),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[10] ),
    .X(\u_usb_host.u_core._149_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._378_  (.A1(net343),
    .A2(net87),
    .B1(\u_usb_host.u_core._149_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[10] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._378__343  (.LO(net343));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._379_  (.A1(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[2] ),
    .A2(net90),
    .B1(net96),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[11] ),
    .X(\u_usb_host.u_core._150_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._380_  (.A1(net344),
    .A2(net87),
    .B1(\u_usb_host.u_core._150_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[11] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._380__344  (.LO(net344));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._381_  (.A1(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[3] ),
    .A2(net90),
    .B1(net96),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[12] ),
    .X(\u_usb_host.u_core._151_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._382_  (.A1(net345),
    .A2(net87),
    .B1(\u_usb_host.u_core._151_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[12] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._382__345  (.LO(net345));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._383_  (.A1(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[4] ),
    .A2(net90),
    .B1(net96),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[13] ),
    .X(\u_usb_host.u_core._152_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._384_  (.A1(net346),
    .A2(net87),
    .B1(\u_usb_host.u_core._152_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[13] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._384__346  (.LO(net346));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._385_  (.A1(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[5] ),
    .A2(net90),
    .B1(net95),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[14] ),
    .X(\u_usb_host.u_core._153_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._386_  (.A1(net347),
    .A2(net87),
    .B1(\u_usb_host.u_core._153_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[14] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._386__347  (.LO(net347));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._387_  (.A1(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[6] ),
    .A2(net90),
    .B1(net95),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[15] ),
    .X(\u_usb_host.u_core._154_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._388_  (.A1(net348),
    .A2(net88),
    .B1(\u_usb_host.u_core._154_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[15] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._388__348  (.LO(net348));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._389_  (.A1(net448),
    .A2(net91),
    .B1(net92),
    .B2(\u_usb_host.u_core.sof_time_q[13] ),
    .X(\u_usb_host.u_core._155_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._390_  (.A1(net350),
    .A2(net88),
    .B1(\u_usb_host.u_core._155_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[29] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._390__350  (.LO(net350));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._391_  (.A1(net447),
    .A2(net91),
    .B1(net93),
    .B2(\u_usb_host.u_core.sof_time_q[12] ),
    .X(\u_usb_host.u_core._156_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._392_  (.A1(net377),
    .A2(\u_usb_host.u_core._117_ ),
    .B1(\u_usb_host.u_core._156_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[28] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core._392__377  (.HI(net377));
 sky130_fd_sc_hd__or3b_1 \u_usb_host.u_core._393_  (.A(\u_usb_host.reg_ack ),
    .B(\u_usb_host.reg_wr ),
    .C_N(\u_usb_host.reg_cs ),
    .X(\u_usb_host.u_core._046_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core._394_  (.A(\u_usb_host.u_core._046_ ),
    .Y(\u_usb_host.u_core._033_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core._395_  (.A(\u_usb_host.u_core.cfg_wr ),
    .B(\u_usb_host.reg_wdata[31] ),
    .C(net89),
    .X(\u_usb_host.u_core._032_ ));
 sky130_fd_sc_hd__and3_2 \u_usb_host.u_core._396_  (.A(\u_usb_host.u_core.cfg_wr ),
    .B(\u_usb_host.u_core._085_ ),
    .C(\u_usb_host.u_core._090_ ),
    .X(\u_usb_host.u_core._157_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._397_  (.A(\u_usb_host.reg_wdata[0] ),
    .B(\u_usb_host.u_core._157_ ),
    .X(\u_usb_host.u_core._030_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._398_  (.A(\u_usb_host.reg_wdata[1] ),
    .B(\u_usb_host.u_core._157_ ),
    .X(\u_usb_host.u_core._028_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._399_  (.A(\u_usb_host.reg_wdata[2] ),
    .B(\u_usb_host.u_core._157_ ),
    .X(\u_usb_host.u_core._029_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._400_  (.A(\u_usb_host.reg_wdata[3] ),
    .B(\u_usb_host.u_core._157_ ),
    .X(\u_usb_host.u_core._027_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._402_  (.A(\u_usb_host.u_core._096_ ),
    .B(\u_usb_host.u_core._033_ ),
    .X(\u_usb_host.u_core.u_fifo_rx.pop_i ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._403_  (.A1(\u_usb_host.u_core.usb_irq_mask_done_out_w ),
    .A2(\u_usb_host.u_core.intr_done_q ),
    .B1(\u_usb_host.u_core.device_det_q ),
    .B2(\u_usb_host.u_core.usb_irq_mask_device_detect_out_w ),
    .X(\u_usb_host.u_core._158_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core._404_  (.A1(\u_usb_host.u_core.usb_irq_mask_sof_out_w ),
    .A2(\u_usb_host.u_core.intr_sof_q ),
    .B1(\u_usb_host.u_core.usb_irq_mask_err_out_w ),
    .B2(\u_usb_host.u_core.intr_err_q ),
    .C1(\u_usb_host.u_core._158_ ),
    .X(\u_usb_host.u_core._005_ ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._427_  (.CLK(\u_usb_host.u_core._179_ ),
    .D(\u_usb_host.u_core._032_ ),
    .RESET_B(net265),
    .Q(\u_usb_host.u_core.usb_rx_stat_start_pend_in_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._428_  (.CLK(\u_usb_host.u_core._181_ ),
    .D(\u_usb_host.reg_wdata[29] ),
    .RESET_B(net264),
    .Q(\u_usb_host.u_core.usb_xfer_token_ack_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._429_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[0] ),
    .RESET_B(net273),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._430_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[1] ),
    .RESET_B(net276),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._431_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[2] ),
    .RESET_B(net275),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._432_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[3] ),
    .RESET_B(net276),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._433_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[4] ),
    .RESET_B(net276),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._434_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[5] ),
    .RESET_B(net276),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._435_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[6] ),
    .RESET_B(net272),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[6] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._436_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[7] ),
    .RESET_B(net275),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[7] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._437_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[8] ),
    .RESET_B(net272),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[8] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._438_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[9] ),
    .RESET_B(net274),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[9] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._439_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[10] ),
    .RESET_B(net277),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[10] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._440_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[11] ),
    .RESET_B(net274),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[11] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._441_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[12] ),
    .RESET_B(net281),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[12] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._442_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[13] ),
    .RESET_B(net281),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[13] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._443_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[14] ),
    .RESET_B(net274),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[14] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._444_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[15] ),
    .RESET_B(net274),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[15] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._445_  (.CLK(\u_usb_host.u_core._180_ ),
    .D(\u_usb_host.reg_wdata[30] ),
    .RESET_B(net264),
    .Q(\u_usb_host.u_core.usb_xfer_token_in_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._446_  (.CLK(\u_usb_host.u_core._175_ ),
    .D(\u_usb_host.reg_wdata[2] ),
    .RESET_B(net279),
    .Q(\u_usb_host.u_core.usb_irq_mask_err_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._447_  (.CLK(\u_usb_host.u_core._176_ ),
    .D(\u_usb_host.reg_wdata[1] ),
    .RESET_B(net279),
    .Q(\u_usb_host.u_core.usb_irq_mask_done_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._448_  (.CLK(\u_usb_host.u_core._177_ ),
    .D(\u_usb_host.reg_wdata[0] ),
    .RESET_B(net278),
    .Q(\u_usb_host.u_core.usb_irq_mask_sof_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._449_  (.CLK(\u_usb_host.u_core._182_ ),
    .D(\u_usb_host.reg_wdata[28] ),
    .RESET_B(net264),
    .Q(\u_usb_host.u_core.u_sie.data_idx_i ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._450_  (.CLK(\u_usb_host.u_core._199_ ),
    .D(\u_usb_host.reg_wdata[5] ),
    .RESET_B(net276),
    .Q(\u_usb_host.u_core.utmi_termselect_o ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._451_  (.CLK(\u_usb_host.u_core._198_ ),
    .D(\u_usb_host.u_core._000_ ),
    .RESET_B(net287),
    .Q(\u_usb_host.u_core.device_det_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._452_  (.CLK(\u_usb_host.u_core._197_ ),
    .D(\u_usb_host.u_core._004_ ),
    .RESET_B(net278),
    .Q(\u_usb_host.u_core.intr_err_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._453_  (.CLK(\u_usb_host.u_core._196_ ),
    .D(net417),
    .RESET_B(net278),
    .Q(\u_usb_host.u_core.intr_sof_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._454_  (.CLK(\u_usb_host.u_core._195_ ),
    .D(\u_usb_host.u_core._003_ ),
    .RESET_B(net279),
    .Q(\u_usb_host.u_core.intr_done_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._455_  (.CLK(\u_usb_host.u_core._194_ ),
    .D(\u_usb_host.u_core._026_ ),
    .RESET_B(net280),
    .Q(\u_usb_host.u_core.usb_err_q ));
 sky130_fd_sc_hd__dfrtp_4 \u_usb_host.u_core._456_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._007_ ),
    .RESET_B(net267),
    .Q(\u_usb_host.u_core.sof_time_q[0] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core._457_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._014_ ),
    .RESET_B(net267),
    .Q(\u_usb_host.u_core.sof_time_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._458_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._015_ ),
    .RESET_B(net267),
    .Q(\u_usb_host.u_core.sof_time_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._459_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._016_ ),
    .RESET_B(net267),
    .Q(\u_usb_host.u_core.sof_time_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._460_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._017_ ),
    .RESET_B(net267),
    .Q(\u_usb_host.u_core.sof_time_q[4] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core._461_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._018_ ),
    .RESET_B(net268),
    .Q(\u_usb_host.u_core.sof_time_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._462_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._019_ ),
    .RESET_B(net267),
    .Q(\u_usb_host.u_core.sof_time_q[6] ));
 sky130_fd_sc_hd__dfrtp_4 \u_usb_host.u_core._463_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._020_ ),
    .RESET_B(net267),
    .Q(\u_usb_host.u_core.sof_time_q[7] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core._464_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._021_ ),
    .RESET_B(net268),
    .Q(\u_usb_host.u_core.sof_time_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._465_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._022_ ),
    .RESET_B(net268),
    .Q(\u_usb_host.u_core.sof_time_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._466_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._008_ ),
    .RESET_B(net270),
    .Q(\u_usb_host.u_core.sof_time_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._467_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._009_ ),
    .RESET_B(net270),
    .Q(\u_usb_host.u_core.sof_time_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._468_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._010_ ),
    .RESET_B(net270),
    .Q(\u_usb_host.u_core.sof_time_q[12] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core._469_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._011_ ),
    .RESET_B(net270),
    .Q(\u_usb_host.u_core.sof_time_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._470_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._012_ ),
    .RESET_B(net270),
    .Q(\u_usb_host.u_core.sof_time_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._471_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._013_ ),
    .RESET_B(net270),
    .Q(\u_usb_host.u_core.sof_time_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._486_  (.CLK(\u_usb_host.u_core._187_ ),
    .D(\u_usb_host.reg_wdata[6] ),
    .RESET_B(net273),
    .Q(\u_usb_host.u_core.utmi_dppulldown_o ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._495_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._185_ ),
    .D(\u_usb_host.reg_wdata[5] ),
    .RESET_B(net275),
    .Q(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._496_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._185_ ),
    .D(\u_usb_host.reg_wdata[6] ),
    .RESET_B(net272),
    .Q(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._497_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._185_ ),
    .D(\u_usb_host.reg_wdata[7] ),
    .RESET_B(net275),
    .Q(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._498_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._185_ ),
    .D(\u_usb_host.reg_wdata[8] ),
    .RESET_B(net273),
    .Q(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._499_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._184_ ),
    .D(\u_usb_host.reg_wdata[9] ),
    .RESET_B(net274),
    .Q(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._500_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._184_ ),
    .D(\u_usb_host.reg_wdata[10] ),
    .RESET_B(net277),
    .Q(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._501_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._184_ ),
    .D(\u_usb_host.reg_wdata[11] ),
    .RESET_B(net274),
    .Q(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._502_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._184_ ),
    .D(\u_usb_host.reg_wdata[12] ),
    .RESET_B(net281),
    .Q(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._503_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._184_ ),
    .D(\u_usb_host.reg_wdata[13] ),
    .RESET_B(net281),
    .Q(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._504_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._184_ ),
    .D(\u_usb_host.reg_wdata[14] ),
    .RESET_B(net274),
    .Q(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._505_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._184_ ),
    .D(\u_usb_host.reg_wdata[15] ),
    .RESET_B(net274),
    .Q(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[6] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._506_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._183_ ),
    .D(\u_usb_host.reg_wdata[16] ),
    .RESET_B(net266),
    .Q(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._507_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._183_ ),
    .D(\u_usb_host.reg_wdata[17] ),
    .RESET_B(net266),
    .Q(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._508_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._183_ ),
    .D(\u_usb_host.reg_wdata[18] ),
    .RESET_B(net266),
    .Q(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._509_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._183_ ),
    .D(\u_usb_host.reg_wdata[19] ),
    .RESET_B(net266),
    .Q(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._510_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._183_ ),
    .D(\u_usb_host.reg_wdata[20] ),
    .RESET_B(net266),
    .Q(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._511_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._183_ ),
    .D(\u_usb_host.reg_wdata[21] ),
    .RESET_B(net266),
    .Q(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._512_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._183_ ),
    .D(\u_usb_host.reg_wdata[22] ),
    .RESET_B(net266),
    .Q(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[6] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._513_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._183_ ),
    .D(\u_usb_host.reg_wdata[23] ),
    .RESET_B(net266),
    .Q(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[7] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._514_  (.CLK(\u_usb_host.u_core._174_ ),
    .D(\u_usb_host.reg_wdata[3] ),
    .RESET_B(net279),
    .Q(\u_usb_host.u_core.usb_irq_mask_device_detect_out_w ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core._515_  (.CLK(\u_usb_host.u_core._173_ ),
    .D(\u_usb_host.reg_wdata[0] ),
    .RESET_B(net278),
    .Q(\u_usb_host.u_core.usb_ctrl_enable_sof_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._516_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._172_ ),
    .D(\u_usb_host.reg_wdata[1] ),
    .RESET_B(net275),
    .Q(\u_usb_host.u_core.utmi_op_mode_o[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._517_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._172_ ),
    .D(\u_usb_host.reg_wdata[2] ),
    .RESET_B(net275),
    .Q(\u_usb_host.u_core.utmi_op_mode_o[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._518_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core._200_ ),
    .D(net428),
    .RESET_B(net272),
    .Q(\u_usb_host.reg_rdata[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._519_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core._200_ ),
    .D(net398),
    .RESET_B(net291),
    .Q(\u_usb_host.reg_rdata[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._520_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core._200_ ),
    .D(net395),
    .RESET_B(net275),
    .Q(\u_usb_host.reg_rdata[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._521_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[3] ),
    .RESET_B(net276),
    .Q(\u_usb_host.reg_rdata[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._522_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[4] ),
    .RESET_B(net276),
    .Q(\u_usb_host.reg_rdata[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._523_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[5] ),
    .RESET_B(net275),
    .Q(\u_usb_host.reg_rdata[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._524_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[6] ),
    .RESET_B(net272),
    .Q(\u_usb_host.reg_rdata[6] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._525_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[7] ),
    .RESET_B(net275),
    .Q(\u_usb_host.reg_rdata[7] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._526_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[8] ),
    .RESET_B(net273),
    .Q(\u_usb_host.reg_rdata[8] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._527_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[9] ),
    .RESET_B(net277),
    .Q(\u_usb_host.reg_rdata[9] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._528_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[10] ),
    .RESET_B(net281),
    .Q(\u_usb_host.reg_rdata[10] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._529_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[11] ),
    .RESET_B(net276),
    .Q(\u_usb_host.reg_rdata[11] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._530_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[12] ),
    .RESET_B(net281),
    .Q(\u_usb_host.reg_rdata[12] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._531_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[13] ),
    .RESET_B(net281),
    .Q(\u_usb_host.reg_rdata[13] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._532_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[14] ),
    .RESET_B(net274),
    .Q(\u_usb_host.reg_rdata[14] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._533_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[15] ),
    .RESET_B(net274),
    .Q(\u_usb_host.reg_rdata[15] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._534_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[16] ),
    .RESET_B(net272),
    .Q(\u_usb_host.reg_rdata[16] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._535_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[17] ),
    .RESET_B(net272),
    .Q(\u_usb_host.reg_rdata[17] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._536_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[18] ),
    .RESET_B(net265),
    .Q(\u_usb_host.reg_rdata[18] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._537_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[19] ),
    .RESET_B(net265),
    .Q(\u_usb_host.reg_rdata[19] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._538_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[20] ),
    .RESET_B(net265),
    .Q(\u_usb_host.reg_rdata[20] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._539_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[21] ),
    .RESET_B(net265),
    .Q(\u_usb_host.reg_rdata[21] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._540_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[22] ),
    .RESET_B(net265),
    .Q(\u_usb_host.reg_rdata[22] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._541_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[23] ),
    .RESET_B(net265),
    .Q(\u_usb_host.reg_rdata[23] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._542_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[24] ),
    .RESET_B(net266),
    .Q(\u_usb_host.reg_rdata[24] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._543_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[25] ),
    .RESET_B(net266),
    .Q(\u_usb_host.reg_rdata[25] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._544_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[26] ),
    .RESET_B(net265),
    .Q(\u_usb_host.reg_rdata[26] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._545_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[27] ),
    .RESET_B(net265),
    .Q(\u_usb_host.reg_rdata[27] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._546_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[28] ),
    .RESET_B(net272),
    .Q(\u_usb_host.reg_rdata[28] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._547_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[29] ),
    .RESET_B(net272),
    .Q(\u_usb_host.reg_rdata[29] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._548_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[30] ),
    .RESET_B(net272),
    .Q(\u_usb_host.reg_rdata[30] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._549_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[31] ),
    .RESET_B(net265),
    .Q(\u_usb_host.reg_rdata[31] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._550_  (.CLK(\u_usb_host.u_core._188_ ),
    .D(\u_usb_host.u_core._002_ ),
    .RESET_B(net278),
    .Q(\u_usb_host.u_core.fifo_flush_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._551_  (.CLK(\u_usb_host.u_core._202_ ),
    .D(\u_usb_host.reg_wdata[7] ),
    .RESET_B(net275),
    .Q(\u_usb_host.u_core.utmi_dmpulldown_o ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core._552_  (.CLK(\u_usb_host.u_core._201_ ),
    .D(\u_usb_host.u_core._047_ ),
    .RESET_B(net264),
    .Q(\u_usb_host.u_core.cfg_wr ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._553_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._171_ ),
    .D(\u_usb_host.reg_wdata[3] ),
    .RESET_B(net276),
    .Q(\u_usb_host.u_core.utmi_xcvrselect_o[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._554_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._171_ ),
    .D(\u_usb_host.reg_wdata[4] ),
    .RESET_B(net276),
    .Q(\u_usb_host.u_core.utmi_xcvrselect_o[1] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core._555_  (.CLK(clknet_4_3_0_usb_clk),
    .D(\u_usb_host.u_core._006_ ),
    .RESET_B(net292),
    .Q(\u_usb_host.reg_ack ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._556_  (.CLK(clknet_4_11_0_usb_clk),
    .D(\u_usb_host.u_core._025_ ),
    .RESET_B(net280),
    .Q(\u_usb_host.u_core.usb_ctrl_wr_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._558_  (.CLK(clknet_4_8_0_usb_clk),
    .D(\u_usb_host.u_core._027_ ),
    .RESET_B(net280),
    .Q(\u_usb_host.u_core.usb_irq_ack_device_detect_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._559_  (.CLK(clknet_4_6_0_usb_clk),
    .D(\u_usb_host.u_core._029_ ),
    .RESET_B(net278),
    .Q(\u_usb_host.u_core.usb_irq_ack_err_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._560_  (.CLK(clknet_4_9_0_usb_clk),
    .D(\u_usb_host.u_core._028_ ),
    .RESET_B(net279),
    .Q(\u_usb_host.u_core.usb_irq_ack_done_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._561_  (.CLK(clknet_4_9_0_usb_clk),
    .D(\u_usb_host.u_core._030_ ),
    .RESET_B(net278),
    .Q(\u_usb_host.u_core.usb_irq_ack_sof_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._563_  (.CLK(clknet_4_6_0_usb_clk),
    .D(\u_usb_host.u_core._023_ ),
    .RESET_B(net278),
    .Q(\u_usb_host.u_core.transfer_start_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._564_  (.CLK(clknet_4_9_0_usb_clk),
    .D(\u_usb_host.u_core.send_sof_w ),
    .RESET_B(net278),
    .Q(\u_usb_host.u_core.sof_irq_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._565_  (.CLK(clknet_4_6_0_usb_clk),
    .D(\u_usb_host.u_core._001_ ),
    .RESET_B(net278),
    .Q(\u_usb_host.u_core.err_cond_q ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core._566_  (.CLK(clknet_4_9_0_usb_clk),
    .D(\u_usb_host.u_core._005_ ),
    .RESET_B(net279),
    .Q(net81));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._567_  (.CLK(clknet_4_10_0_usb_clk),
    .GATE(\u_usb_host.u_core._025_ ),
    .GCLK(\u_usb_host.u_core._171_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._568_  (.CLK(clknet_4_8_0_usb_clk),
    .GATE(\u_usb_host.u_core._025_ ),
    .GCLK(\u_usb_host.u_core._172_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._569_  (.CLK(clknet_4_8_0_usb_clk),
    .GATE(\u_usb_host.u_core._025_ ),
    .GCLK(\u_usb_host.u_core._173_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._570_  (.CLK(clknet_4_8_0_usb_clk),
    .GATE(\u_usb_host.u_core._034_ ),
    .GCLK(\u_usb_host.u_core._174_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._571_  (.CLK(clknet_4_9_0_usb_clk),
    .GATE(\u_usb_host.u_core._034_ ),
    .GCLK(\u_usb_host.u_core._175_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._572_  (.CLK(clknet_4_8_0_usb_clk),
    .GATE(\u_usb_host.u_core._034_ ),
    .GCLK(\u_usb_host.u_core._176_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._573_  (.CLK(clknet_4_9_0_usb_clk),
    .GATE(\u_usb_host.u_core._034_ ),
    .GCLK(\u_usb_host.u_core._177_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core._574_  (.CLK(clknet_4_8_0_usb_clk),
    .GATE(\u_usb_host.u_core._035_ ),
    .GCLK(\u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._575_  (.CLK(clknet_4_6_0_usb_clk),
    .GATE(\u_usb_host.u_core._036_ ),
    .GCLK(\u_usb_host.u_core._179_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._576_  (.CLK(clknet_4_3_0_usb_clk),
    .GATE(\u_usb_host.u_core._037_ ),
    .GCLK(\u_usb_host.u_core._180_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._577_  (.CLK(clknet_4_3_0_usb_clk),
    .GATE(\u_usb_host.u_core._037_ ),
    .GCLK(\u_usb_host.u_core._181_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._578_  (.CLK(clknet_4_3_0_usb_clk),
    .GATE(\u_usb_host.u_core._037_ ),
    .GCLK(\u_usb_host.u_core._182_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core._579_  (.CLK(clknet_4_2_0_usb_clk),
    .GATE(\u_usb_host.u_core._037_ ),
    .GCLK(\u_usb_host.u_core._183_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core._580_  (.CLK(clknet_4_8_0_usb_clk),
    .GATE(\u_usb_host.u_core._037_ ),
    .GCLK(\u_usb_host.u_core._184_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._581_  (.CLK(clknet_4_8_0_usb_clk),
    .GATE(\u_usb_host.u_core._037_ ),
    .GCLK(\u_usb_host.u_core._185_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._583_  (.CLK(clknet_4_8_0_usb_clk),
    .GATE(\u_usb_host.u_core._025_ ),
    .GCLK(\u_usb_host.u_core._187_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._584_  (.CLK(clknet_4_6_0_usb_clk),
    .GATE(\u_usb_host.u_core._038_ ),
    .GCLK(\u_usb_host.u_core._188_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core._589_  (.CLK(clknet_4_6_0_usb_clk),
    .GATE(\u_usb_host.u_core._040_ ),
    .GCLK(\u_usb_host.u_core._193_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._590_  (.CLK(clknet_4_11_0_usb_clk),
    .GATE(\u_usb_host.u_core._041_ ),
    .GCLK(\u_usb_host.u_core._194_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._591_  (.CLK(clknet_4_9_0_usb_clk),
    .GATE(\u_usb_host.u_core._042_ ),
    .GCLK(\u_usb_host.u_core._195_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._592_  (.CLK(clknet_4_6_0_usb_clk),
    .GATE(\u_usb_host.u_core._043_ ),
    .GCLK(\u_usb_host.u_core._196_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._593_  (.CLK(clknet_4_6_0_usb_clk),
    .GATE(\u_usb_host.u_core._044_ ),
    .GCLK(\u_usb_host.u_core._197_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._594_  (.CLK(clknet_4_9_0_usb_clk),
    .GATE(\u_usb_host.u_core._045_ ),
    .GCLK(\u_usb_host.u_core._198_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._595_  (.CLK(clknet_4_8_0_usb_clk),
    .GATE(\u_usb_host.u_core._025_ ),
    .GCLK(\u_usb_host.u_core._199_ ));
 sky130_fd_sc_hd__dlclkp_4 \u_usb_host.u_core._596_  (.CLK(clknet_4_6_0_usb_clk),
    .GATE(\u_usb_host.u_core._033_ ),
    .GCLK(\u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._597_  (.CLK(clknet_4_2_0_usb_clk),
    .GATE(\u_usb_host.u_core._046_ ),
    .GCLK(\u_usb_host.u_core._201_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._598_  (.CLK(clknet_4_8_0_usb_clk),
    .GATE(\u_usb_host.u_core._025_ ),
    .GCLK(\u_usb_host.u_core._202_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_fifo_rx._0784_  (.A(\u_usb_host.u_core.u_fifo_rx.count[6] ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0438_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_core.u_fifo_rx._0785_  (.A(\u_usb_host.u_core.u_fifo_rx.count[2] ),
    .B(\u_usb_host.u_core.u_fifo_rx.count[0] ),
    .C(\u_usb_host.u_core.u_fifo_rx.count[1] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0439_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_rx._0786_  (.A(\u_usb_host.u_core.u_fifo_rx.count[3] ),
    .B(\u_usb_host.u_core.u_fifo_rx.count[2] ),
    .C(\u_usb_host.u_core.u_fifo_rx.count[0] ),
    .D(\u_usb_host.u_core.u_fifo_rx.count[1] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0440_ ));
 sky130_fd_sc_hd__or3_2 \u_usb_host.u_core.u_fifo_rx._0787_  (.A(\u_usb_host.u_core.u_fifo_rx.count[5] ),
    .B(\u_usb_host.u_core.u_fifo_rx.count[4] ),
    .C(\u_usb_host.u_core.u_fifo_rx._0440_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0441_ ));
 sky130_fd_sc_hd__o21a_2 \u_usb_host.u_core.u_fifo_rx._0789_  (.A1(\u_usb_host.u_core.u_fifo_rx._0438_ ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0441_ ),
    .B1(net367),
    .X(\u_usb_host.u_core.u_fifo_rx._0442_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core.u_fifo_rx._0789__367  (.LO(net367));
 sky130_fd_sc_hd__nand2_2 \u_usb_host.u_core.u_fifo_rx._0790_  (.A(net269),
    .B(\u_usb_host.u_core.u_fifo_rx._0442_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0443_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_rx._0791_  (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[0] ),
    .B(\u_usb_host.u_core.u_fifo_rx.wr_ptr[1] ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0444_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_rx._0792_  (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[2] ),
    .B(net296),
    .Y(\u_usb_host.u_core.u_fifo_rx._0445_ ));
 sky130_fd_sc_hd__and3_2 \u_usb_host.u_core.u_fifo_rx._0793_  (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[0] ),
    .B(\u_usb_host.u_core.u_fifo_rx.wr_ptr[1] ),
    .C(net298),
    .X(\u_usb_host.u_core.u_fifo_rx._0446_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0794_  (.A(\u_usb_host.u_core.u_fifo_rx._0444_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0445_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0447_ ));
 sky130_fd_sc_hd__nand2_2 \u_usb_host.u_core.u_fifo_rx._0795_  (.A(net297),
    .B(\u_usb_host.u_core.u_fifo_rx._0446_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0448_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0796_  (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[5] ),
    .B(\u_usb_host.u_core.u_fifo_rx.wr_ptr[4] ),
    .C(\u_usb_host.u_core.u_fifo_rx._0447_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0449_ ));
 sky130_fd_sc_hd__and3_2 \u_usb_host.u_core.u_fifo_rx._0797_  (.A(net279),
    .B(\u_usb_host.u_core.u_fifo_rx._0442_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0449_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0019_ ));
 sky130_fd_sc_hd__nand4_2 \u_usb_host.u_core.u_fifo_rx._0798_  (.A(net271),
    .B(\u_usb_host.u_core.u_fifo_rx.wr_ptr[5] ),
    .C(\u_usb_host.u_core.u_fifo_rx.wr_ptr[4] ),
    .D(\u_usb_host.u_core.u_fifo_rx._0442_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__nand2b_2 \u_usb_host.u_core.u_fifo_rx._0799_  (.A_N(\u_usb_host.u_core.u_fifo_rx.wr_ptr[1] ),
    .B(\u_usb_host.u_core.u_fifo_rx.wr_ptr[0] ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0451_ ));
 sky130_fd_sc_hd__or2_4 \u_usb_host.u_core.u_fifo_rx._0800_  (.A(\u_usb_host.u_core.u_fifo_rx._0445_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0451_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0452_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0801_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0452_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0020_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_fifo_rx._0802_  (.A(\u_usb_host.u_core.fifo_flush_q ),
    .B(\u_usb_host.u_core.u_fifo_rx._0442_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0023_ ));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_core.u_fifo_rx._0804_  (.A1(\u_usb_host.u_core.u_fifo_rx.count[6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0441_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx.pop_i ),
    .X(\u_usb_host.u_core.u_fifo_rx._0453_ ));
 sky130_fd_sc_hd__o21ai_2 \u_usb_host.u_core.u_fifo_rx._0805_  (.A1(\u_usb_host.u_core.u_fifo_rx.count[6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0441_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx.pop_i ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0454_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_fifo_rx._0806_  (.A(\u_usb_host.u_core.fifo_flush_q ),
    .B(\u_usb_host.u_core.u_fifo_rx._0453_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0024_ ));
 sky130_fd_sc_hd__or4_4 \u_usb_host.u_core.u_fifo_rx._0807_  (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[0] ),
    .B(\u_usb_host.u_core.u_fifo_rx.wr_ptr[1] ),
    .C(\u_usb_host.u_core.u_fifo_rx.wr_ptr[2] ),
    .D(net297),
    .X(\u_usb_host.u_core.u_fifo_rx._0455_ ));
 sky130_fd_sc_hd__or3_2 \u_usb_host.u_core.u_fifo_rx._0808_  (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[5] ),
    .B(\u_usb_host.u_core.u_fifo_rx.wr_ptr[4] ),
    .C(\u_usb_host.u_core.u_fifo_rx._0443_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0809_  (.A(\u_usb_host.u_core.u_fifo_rx._0455_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0456_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0026_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0810_  (.A(\u_usb_host.u_core.u_fifo_rx._0442_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0454_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0457_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0811_  (.A(\u_usb_host.u_core.u_fifo_rx._0442_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0454_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0458_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_core.u_fifo_rx._0812_  (.A(\u_usb_host.u_core.fifo_flush_q ),
    .B(\u_usb_host.u_core.u_fifo_rx._0457_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0458_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0025_ ));
 sky130_fd_sc_hd__nand2b_2 \u_usb_host.u_core.u_fifo_rx._0813_  (.A_N(\u_usb_host.u_core.u_fifo_rx.wr_ptr[0] ),
    .B(\u_usb_host.u_core.u_fifo_rx.wr_ptr[1] ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0459_ ));
 sky130_fd_sc_hd__or2_4 \u_usb_host.u_core.u_fifo_rx._0814_  (.A(\u_usb_host.u_core.u_fifo_rx._0445_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0459_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0460_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0815_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0460_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0021_ ));
 sky130_fd_sc_hd__or3_4 \u_usb_host.u_core.u_fifo_rx._0816_  (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[0] ),
    .B(\u_usb_host.u_core.u_fifo_rx.wr_ptr[1] ),
    .C(\u_usb_host.u_core.u_fifo_rx._0445_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0461_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0817_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0461_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0022_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0818_  (.A(\u_usb_host.u_core.u_fifo_rx._0452_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0456_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0039_ ));
 sky130_fd_sc_hd__or3b_2 \u_usb_host.u_core.u_fifo_rx._0819_  (.A(\u_usb_host.u_core.u_fifo_rx._0443_ ),
    .B(\u_usb_host.u_core.u_fifo_rx.wr_ptr[5] ),
    .C_N(\u_usb_host.u_core.u_fifo_rx.wr_ptr[4] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0820_  (.A(\u_usb_host.u_core.u_fifo_rx._0455_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0462_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0042_ ));
 sky130_fd_sc_hd__or3b_4 \u_usb_host.u_core.u_fifo_rx._0821_  (.A(\u_usb_host.u_core.u_fifo_rx._0444_ ),
    .B(net298),
    .C_N(net297),
    .X(\u_usb_host.u_core.u_fifo_rx._0463_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0822_  (.A(\u_usb_host.u_core.u_fifo_rx._0456_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0463_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0037_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0823_  (.A(\u_usb_host.u_core.u_fifo_rx._0448_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0456_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0041_ ));
 sky130_fd_sc_hd__or3_4 \u_usb_host.u_core.u_fifo_rx._0824_  (.A(net298),
    .B(net296),
    .C(\u_usb_host.u_core.u_fifo_rx._0459_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0464_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0825_  (.A(\u_usb_host.u_core.u_fifo_rx._0462_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0464_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0044_ ));
 sky130_fd_sc_hd__or3_4 \u_usb_host.u_core.u_fifo_rx._0826_  (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[2] ),
    .B(net296),
    .C(\u_usb_host.u_core.u_fifo_rx._0451_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0465_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0827_  (.A(\u_usb_host.u_core.u_fifo_rx._0462_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0465_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0043_ ));
 sky130_fd_sc_hd__or3_4 \u_usb_host.u_core.u_fifo_rx._0828_  (.A(net298),
    .B(net296),
    .C(\u_usb_host.u_core.u_fifo_rx._0444_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0466_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0829_  (.A(\u_usb_host.u_core.u_fifo_rx._0462_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0466_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0045_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0830_  (.A(\u_usb_host.u_core.u_fifo_rx._0461_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0462_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0054_ ));
 sky130_fd_sc_hd__or3b_4 \u_usb_host.u_core.u_fifo_rx._0831_  (.A(net296),
    .B(\u_usb_host.u_core.u_fifo_rx._0459_ ),
    .C_N(net298),
    .X(\u_usb_host.u_core.u_fifo_rx._0467_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0832_  (.A(\u_usb_host.u_core.u_fifo_rx._0462_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0467_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0048_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0833_  (.A(\u_usb_host.u_core.u_fifo_rx._0462_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0463_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0053_ ));
 sky130_fd_sc_hd__or3b_4 \u_usb_host.u_core.u_fifo_rx._0834_  (.A(net296),
    .B(\u_usb_host.u_core.u_fifo_rx._0451_ ),
    .C_N(\u_usb_host.u_core.u_fifo_rx.wr_ptr[2] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0468_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0835_  (.A(\u_usb_host.u_core.u_fifo_rx._0462_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0468_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0047_ ));
 sky130_fd_sc_hd__or3b_4 \u_usb_host.u_core.u_fifo_rx._0836_  (.A(\u_usb_host.u_core.u_fifo_rx._0459_ ),
    .B(net298),
    .C_N(net296),
    .X(\u_usb_host.u_core.u_fifo_rx._0469_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0837_  (.A(\u_usb_host.u_core.u_fifo_rx._0462_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0469_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0052_ ));
 sky130_fd_sc_hd__or3b_4 \u_usb_host.u_core.u_fifo_rx._0838_  (.A(\u_usb_host.u_core.u_fifo_rx._0451_ ),
    .B(net298),
    .C_N(net296),
    .X(\u_usb_host.u_core.u_fifo_rx._0470_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0839_  (.A(\u_usb_host.u_core.u_fifo_rx._0462_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0470_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0051_ ));
 sky130_fd_sc_hd__or4b_4 \u_usb_host.u_core.u_fifo_rx._0840_  (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[0] ),
    .B(\u_usb_host.u_core.u_fifo_rx.wr_ptr[1] ),
    .C(net298),
    .D_N(net296),
    .X(\u_usb_host.u_core.u_fifo_rx._0471_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0841_  (.A(\u_usb_host.u_core.u_fifo_rx._0462_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0471_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0050_ ));
 sky130_fd_sc_hd__or4b_4 \u_usb_host.u_core.u_fifo_rx._0842_  (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[0] ),
    .B(\u_usb_host.u_core.u_fifo_rx.wr_ptr[1] ),
    .C(net296),
    .D_N(net298),
    .X(\u_usb_host.u_core.u_fifo_rx._0472_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0843_  (.A(\u_usb_host.u_core.u_fifo_rx._0462_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0472_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0046_ ));
 sky130_fd_sc_hd__nand2b_4 \u_usb_host.u_core.u_fifo_rx._0844_  (.A_N(net297),
    .B(\u_usb_host.u_core.u_fifo_rx._0446_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0473_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0845_  (.A(\u_usb_host.u_core.u_fifo_rx._0462_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0473_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0049_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0846_  (.A(\u_usb_host.u_core.u_fifo_rx._0456_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0460_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0040_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0847_  (.A(\u_usb_host.u_core.u_fifo_rx._0456_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0461_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0038_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0848_  (.A(\u_usb_host.u_core.u_fifo_rx._0456_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0469_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0036_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0849_  (.A(\u_usb_host.u_core.u_fifo_rx._0456_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0470_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0035_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0850_  (.A(\u_usb_host.u_core.u_fifo_rx._0456_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0471_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0034_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0851_  (.A(\u_usb_host.u_core.u_fifo_rx._0456_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0473_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0033_ ));
 sky130_fd_sc_hd__or3b_2 \u_usb_host.u_core.u_fifo_rx._0852_  (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[4] ),
    .B(\u_usb_host.u_core.u_fifo_rx._0443_ ),
    .C_N(\u_usb_host.u_core.u_fifo_rx.wr_ptr[5] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0853_  (.A(\u_usb_host.u_core.u_fifo_rx._0472_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0062_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0854_  (.A(\u_usb_host.u_core.u_fifo_rx._0466_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0061_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0855_  (.A(\u_usb_host.u_core.u_fifo_rx._0464_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0060_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0856_  (.A(\u_usb_host.u_core.u_fifo_rx._0465_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0059_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0857_  (.A(\u_usb_host.u_core.u_fifo_rx._0455_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0058_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0858_  (.A(\u_usb_host.u_core.u_fifo_rx._0448_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0462_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0057_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0859_  (.A(\u_usb_host.u_core.u_fifo_rx._0460_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0462_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0056_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0860_  (.A(\u_usb_host.u_core.u_fifo_rx._0452_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0462_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0055_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0861_  (.A(\u_usb_host.u_core.u_fifo_rx._0456_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0467_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0032_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0862_  (.A(\u_usb_host.u_core.u_fifo_rx._0456_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0468_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0031_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0863_  (.A(\u_usb_host.u_core.u_fifo_rx._0456_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0472_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0030_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0864_  (.A(\u_usb_host.u_core.u_fifo_rx._0456_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0466_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0029_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0865_  (.A(\u_usb_host.u_core.u_fifo_rx._0456_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0464_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0028_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0866_  (.A(\u_usb_host.u_core.u_fifo_rx._0456_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0465_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0027_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0867_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0464_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0076_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0868_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0465_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0075_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0869_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0455_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0074_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0870_  (.A(\u_usb_host.u_core.u_fifo_rx._0448_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0073_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0871_  (.A(\u_usb_host.u_core.u_fifo_rx._0460_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0072_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0872_  (.A(\u_usb_host.u_core.u_fifo_rx._0452_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0071_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0873_  (.A(\u_usb_host.u_core.u_fifo_rx._0461_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0070_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0874_  (.A(\u_usb_host.u_core.u_fifo_rx._0463_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0069_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0875_  (.A(\u_usb_host.u_core.u_fifo_rx._0469_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0068_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0876_  (.A(\u_usb_host.u_core.u_fifo_rx._0470_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0067_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0877_  (.A(\u_usb_host.u_core.u_fifo_rx._0471_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0066_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0878_  (.A(\u_usb_host.u_core.u_fifo_rx._0467_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0064_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0879_  (.A(\u_usb_host.u_core.u_fifo_rx._0473_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0065_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0880_  (.A(\u_usb_host.u_core.u_fifo_rx._0468_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0063_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0881_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0473_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0081_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0882_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0472_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0078_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0883_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0467_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0080_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0884_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0468_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0079_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0885_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0466_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0077_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0886_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0469_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0084_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0887_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0463_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0085_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0888_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0471_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0082_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0889_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0470_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0083_ ));
 sky130_fd_sc_hd__o21ba_1 \u_usb_host.u_core.u_fifo_rx._0890_  (.A1(\u_usb_host.u_core.u_fifo_rx._0457_ ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0458_ ),
    .B1_N(\u_usb_host.u_core.u_fifo_rx.count[0] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0000_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_fifo_rx._0891_  (.A(\u_usb_host.u_core.u_fifo_rx.count[0] ),
    .B(\u_usb_host.u_core.u_fifo_rx.count[1] ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0475_ ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core.u_fifo_rx._0892_  (.A0(\u_usb_host.u_core.u_fifo_rx._0457_ ),
    .A1(\u_usb_host.u_core.u_fifo_rx._0458_ ),
    .S(\u_usb_host.u_core.u_fifo_rx._0475_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0001_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_fifo_rx._0893_  (.A1(\u_usb_host.u_core.u_fifo_rx.count[0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx.count[1] ),
    .B1(\u_usb_host.u_core.u_fifo_rx.count[2] ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0476_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_rx._0894_  (.A(\u_usb_host.u_core.u_fifo_rx._0439_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0476_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0477_ ));
 sky130_fd_sc_hd__nand3_1 \u_usb_host.u_core.u_fifo_rx._0895_  (.A(\u_usb_host.u_core.u_fifo_rx.count[2] ),
    .B(\u_usb_host.u_core.u_fifo_rx.count[0] ),
    .C(\u_usb_host.u_core.u_fifo_rx.count[1] ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0478_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_fifo_rx._0896_  (.A1(\u_usb_host.u_core.u_fifo_rx.count[0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx.count[1] ),
    .B1(\u_usb_host.u_core.u_fifo_rx.count[2] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0479_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._0897_  (.A1(\u_usb_host.u_core.u_fifo_rx._0457_ ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0478_ ),
    .A3(\u_usb_host.u_core.u_fifo_rx._0479_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0458_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0477_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0002_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_rx._0898_  (.A(\u_usb_host.u_core.u_fifo_rx.count[3] ),
    .B(\u_usb_host.u_core.u_fifo_rx._0439_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0480_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_rx._0899_  (.A(\u_usb_host.u_core.u_fifo_rx._0440_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0480_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0481_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_core.u_fifo_rx._0900_  (.A(\u_usb_host.u_core.u_fifo_rx.count[3] ),
    .B(\u_usb_host.u_core.u_fifo_rx.count[2] ),
    .C(\u_usb_host.u_core.u_fifo_rx.count[0] ),
    .D(\u_usb_host.u_core.u_fifo_rx.count[1] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0482_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_fifo_rx._0901_  (.A(\u_usb_host.u_core.u_fifo_rx._0482_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0483_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_rx._0902_  (.A1(\u_usb_host.u_core.u_fifo_rx.count[2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx.count[0] ),
    .A3(\u_usb_host.u_core.u_fifo_rx.count[1] ),
    .B1(\u_usb_host.u_core.u_fifo_rx.count[3] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0484_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._0903_  (.A1(\u_usb_host.u_core.u_fifo_rx._0457_ ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0483_ ),
    .A3(\u_usb_host.u_core.u_fifo_rx._0484_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0458_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0481_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0003_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_fifo_rx._0904_  (.A(\u_usb_host.u_core.u_fifo_rx.count[4] ),
    .B(\u_usb_host.u_core.u_fifo_rx._0440_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0485_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_fifo_rx._0905_  (.A(\u_usb_host.u_core.u_fifo_rx.count[4] ),
    .B(\u_usb_host.u_core.u_fifo_rx._0482_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0486_ ));
 sky130_fd_sc_hd__o21ai_2 \u_usb_host.u_core.u_fifo_rx._0906_  (.A1(\u_usb_host.u_core.u_fifo_rx.count[4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0482_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0457_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0487_ ));
 sky130_fd_sc_hd__a2bb2o_1 \u_usb_host.u_core.u_fifo_rx._0907_  (.A1_N(\u_usb_host.u_core.u_fifo_rx._0486_ ),
    .A2_N(\u_usb_host.u_core.u_fifo_rx._0487_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0458_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0485_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0004_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_fifo_rx._0908_  (.A1(\u_usb_host.u_core.u_fifo_rx.count[4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0440_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx.count[5] ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0488_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_rx._0909_  (.A(\u_usb_host.u_core.u_fifo_rx._0441_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0488_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0489_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0910_  (.A(\u_usb_host.u_core.u_fifo_rx.count[5] ),
    .B(\u_usb_host.u_core.u_fifo_rx.count[4] ),
    .C(\u_usb_host.u_core.u_fifo_rx._0482_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0490_ ));
 sky130_fd_sc_hd__o21ai_2 \u_usb_host.u_core.u_fifo_rx._0911_  (.A1(\u_usb_host.u_core.u_fifo_rx.count[5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0486_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0457_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0491_ ));
 sky130_fd_sc_hd__a2bb2o_1 \u_usb_host.u_core.u_fifo_rx._0912_  (.A1_N(\u_usb_host.u_core.u_fifo_rx._0490_ ),
    .A2_N(\u_usb_host.u_core.u_fifo_rx._0491_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0458_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0489_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0005_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_fifo_rx._0913_  (.A(\u_usb_host.u_core.u_fifo_rx._0438_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0490_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0492_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._0914_  (.A1(\u_usb_host.u_core.u_fifo_rx.count[6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0441_ ),
    .A3(\u_usb_host.u_core.u_fifo_rx._0458_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0492_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0457_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0006_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0915_  (.A(net305),
    .B(\u_usb_host.u_core.u_fifo_rx._0454_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0007_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_rx._0916_  (.A(net305),
    .B(net303),
    .Y(\u_usb_host.u_core.u_fifo_rx._0493_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_fifo_rx._0917_  (.A(net305),
    .B(net303),
    .X(\u_usb_host.u_core.u_fifo_rx._0494_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0918_  (.A(\u_usb_host.u_core.u_fifo_rx._0453_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0493_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0494_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0008_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_fifo_rx._0919_  (.A1(net305),
    .A2(net303),
    .B1(net301),
    .X(\u_usb_host.u_core.u_fifo_rx._0495_ ));
 sky130_fd_sc_hd__nand3_1 \u_usb_host.u_core.u_fifo_rx._0920_  (.A(net305),
    .B(net303),
    .C(net301),
    .Y(\u_usb_host.u_core.u_fifo_rx._0496_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0921_  (.A(\u_usb_host.u_core.u_fifo_rx._0453_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0495_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0496_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0009_ ));
 sky130_fd_sc_hd__and4b_2 \u_usb_host.u_core.u_fifo_rx._0922_  (.A_N(net299),
    .B(net301),
    .C(net304),
    .D(net305),
    .X(\u_usb_host.u_core.u_fifo_rx._0497_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_fifo_rx._0923_  (.A(net299),
    .B(\u_usb_host.u_core.u_fifo_rx._0496_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0498_ ));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_core.u_fifo_rx._0924_  (.A1(net259),
    .A2(\u_usb_host.u_core.u_fifo_rx._0498_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0453_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0010_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_core.u_fifo_rx._0925_  (.A(net306),
    .B(net303),
    .C(net301),
    .D(net299),
    .X(\u_usb_host.u_core.u_fifo_rx._0499_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_fifo_rx._0926_  (.A1(\u_usb_host.u_core.u_fifo_rx.rd_ptr[4] ),
    .A2(net256),
    .B1(\u_usb_host.u_core.u_fifo_rx._0453_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0500_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_core.u_fifo_rx._0927_  (.A1(\u_usb_host.u_core.u_fifo_rx.rd_ptr[4] ),
    .A2(net256),
    .B1(\u_usb_host.u_core.u_fifo_rx._0500_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0011_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_core.u_fifo_rx._0928_  (.A_N(\u_usb_host.u_core.u_fifo_rx.rd_ptr[5] ),
    .B(\u_usb_host.u_core.u_fifo_rx.rd_ptr[4] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0501_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_fifo_rx._0929_  (.A(\u_usb_host.u_core.u_fifo_rx.rd_ptr[4] ),
    .B(\u_usb_host.u_core.u_fifo_rx.rd_ptr[5] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0502_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_core.u_fifo_rx._0930_  (.A1(\u_usb_host.u_core.u_fifo_rx.rd_ptr[4] ),
    .A2(net256),
    .B1(\u_usb_host.u_core.u_fifo_rx.rd_ptr[5] ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0503_ ));
 sky130_fd_sc_hd__a211oi_1 \u_usb_host.u_core.u_fifo_rx._0931_  (.A1(net256),
    .A2(net243),
    .B1(\u_usb_host.u_core.u_fifo_rx._0503_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0454_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0012_ ));
 sky130_fd_sc_hd__and2b_2 \u_usb_host.u_core.u_fifo_rx._0932_  (.A_N(\u_usb_host.u_core.u_fifo_rx.wr_ptr[0] ),
    .B(\u_usb_host.u_core.u_fifo_rx._0442_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0013_ ));
 sky130_fd_sc_hd__a21boi_2 \u_usb_host.u_core.u_fifo_rx._0933_  (.A1(\u_usb_host.u_core.u_fifo_rx._0451_ ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0459_ ),
    .B1_N(\u_usb_host.u_core.u_fifo_rx._0442_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0014_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_fifo_rx._0934_  (.A1(\u_usb_host.u_core.u_fifo_rx.wr_ptr[0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx.wr_ptr[1] ),
    .B1(net298),
    .X(\u_usb_host.u_core.u_fifo_rx._0504_ ));
 sky130_fd_sc_hd__and3b_2 \u_usb_host.u_core.u_fifo_rx._0935_  (.A_N(\u_usb_host.u_core.u_fifo_rx._0446_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0504_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0442_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0015_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_fifo_rx._0936_  (.A(net297),
    .B(\u_usb_host.u_core.u_fifo_rx._0446_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0505_ ));
 sky130_fd_sc_hd__and3_2 \u_usb_host.u_core.u_fifo_rx._0937_  (.A(\u_usb_host.u_core.u_fifo_rx._0442_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0448_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0505_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0016_ ));
 sky130_fd_sc_hd__o21ai_2 \u_usb_host.u_core.u_fifo_rx._0938_  (.A1(\u_usb_host.u_core.u_fifo_rx.wr_ptr[4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0447_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0442_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0506_ ));
 sky130_fd_sc_hd__a21oi_2 \u_usb_host.u_core.u_fifo_rx._0939_  (.A1(\u_usb_host.u_core.u_fifo_rx.wr_ptr[4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0447_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0506_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0017_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_rx._0940_  (.A1(net297),
    .A2(\u_usb_host.u_core.u_fifo_rx.wr_ptr[4] ),
    .A3(\u_usb_host.u_core.u_fifo_rx._0446_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx.wr_ptr[5] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0507_ ));
 sky130_fd_sc_hd__and3b_2 \u_usb_host.u_core.u_fifo_rx._0941_  (.A_N(\u_usb_host.u_core.u_fifo_rx._0449_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0507_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0442_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0018_ ));
 sky130_fd_sc_hd__nor4_2 \u_usb_host.u_core.u_fifo_rx._0942_  (.A(net306),
    .B(net303),
    .C(net301),
    .D(net299),
    .Y(\u_usb_host.u_core.u_fifo_rx._0508_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0943_  (.A(\u_usb_host.u_core.u_fifo_rx.rd_ptr[4] ),
    .B(\u_usb_host.u_core.u_fifo_rx.rd_ptr[5] ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0509_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0944_  (.A(net229),
    .B(net226),
    .X(\u_usb_host.u_core.u_fifo_rx._0510_ ));
 sky130_fd_sc_hd__nand2_2 \u_usb_host.u_core.u_fifo_rx._0945_  (.A(net229),
    .B(net226),
    .Y(\u_usb_host.u_core.u_fifo_rx._0511_ ));
 sky130_fd_sc_hd__and4bb_2 \u_usb_host.u_core.u_fifo_rx._0946_  (.A_N(net303),
    .B_N(net301),
    .C(net299),
    .D(net305),
    .X(\u_usb_host.u_core.u_fifo_rx._0512_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0947_  (.A(net252),
    .B(net219),
    .X(\u_usb_host.u_core.u_fifo_rx._0513_ ));
 sky130_fd_sc_hd__nor4b_4 \u_usb_host.u_core.u_fifo_rx._0948_  (.A(net306),
    .B(net304),
    .C(net302),
    .D_N(net299),
    .Y(\u_usb_host.u_core.u_fifo_rx._0514_ ));
 sky130_fd_sc_hd__and2b_2 \u_usb_host.u_core.u_fifo_rx._0949_  (.A_N(\u_usb_host.u_core.u_fifo_rx.rd_ptr[4] ),
    .B(\u_usb_host.u_core.u_fifo_rx.rd_ptr[5] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0515_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0950_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[40][0] ),
    .B(net217),
    .C(net212),
    .X(\u_usb_host.u_core.u_fifo_rx._0516_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0951_  (.A(net252),
    .B(\u_usb_host.u_core.u_fifo_rx._0514_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0517_ ));
 sky130_fd_sc_hd__nor4b_4 \u_usb_host.u_core.u_fifo_rx._0952_  (.A(\u_usb_host.u_core.u_fifo_rx.rd_ptr[0] ),
    .B(net302),
    .C(net300),
    .D_N(net304),
    .Y(\u_usb_host.u_core.u_fifo_rx._0518_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0953_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[34][0] ),
    .B(net210),
    .C(net200),
    .X(\u_usb_host.u_core.u_fifo_rx._0519_ ));
 sky130_fd_sc_hd__and4b_1 \u_usb_host.u_core.u_fifo_rx._0954_  (.A_N(net301),
    .B(net299),
    .C(net305),
    .D(net304),
    .X(\u_usb_host.u_core.u_fifo_rx._0520_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0955_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[43][0] ),
    .B(net206),
    .C(net196),
    .X(\u_usb_host.u_core.u_fifo_rx._0521_ ));
 sky130_fd_sc_hd__nor4b_4 \u_usb_host.u_core.u_fifo_rx._0956_  (.A(\u_usb_host.u_core.u_fifo_rx.rd_ptr[1] ),
    .B(net302),
    .C(net300),
    .D_N(net306),
    .Y(\u_usb_host.u_core.u_fifo_rx._0522_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0957_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[17][0] ),
    .B(net244),
    .C(net193),
    .X(\u_usb_host.u_core.u_fifo_rx._0523_ ));
 sky130_fd_sc_hd__and4bb_1 \u_usb_host.u_core.u_fifo_rx._0958_  (.A_N(net306),
    .B_N(net302),
    .C(net300),
    .D(net304),
    .X(\u_usb_host.u_core.u_fifo_rx._0524_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0959_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[58][0] ),
    .B(net237),
    .C(net191),
    .X(\u_usb_host.u_core.u_fifo_rx._0525_ ));
 sky130_fd_sc_hd__and4bb_4 \u_usb_host.u_core.u_fifo_rx._0960_  (.A_N(net302),
    .B_N(net300),
    .C(net306),
    .D(net304),
    .X(\u_usb_host.u_core.u_fifo_rx._0526_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0961_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[35][0] ),
    .B(net214),
    .C(net189),
    .X(\u_usb_host.u_core.u_fifo_rx._0527_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0962_  (.A(net224),
    .B(net219),
    .X(\u_usb_host.u_core.u_fifo_rx._0528_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0963_  (.A(net224),
    .B(net196),
    .X(\u_usb_host.u_core.u_fifo_rx._0529_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0964_  (.A(net235),
    .B(\u_usb_host.u_core.u_fifo_rx._0514_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0530_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0965_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[50][0] ),
    .B(net234),
    .C(net198),
    .X(\u_usb_host.u_core.u_fifo_rx._0531_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0966_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[16][0] ),
    .B(net244),
    .C(net227),
    .X(\u_usb_host.u_core.u_fifo_rx._0532_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0967_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[57][0] ),
    .B(net239),
    .C(net220),
    .X(\u_usb_host.u_core.u_fifo_rx._0533_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0968_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[48][0] ),
    .B(net230),
    .C(net227),
    .X(\u_usb_host.u_core.u_fifo_rx._0534_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0969_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[18][0] ),
    .B(net246),
    .C(net198),
    .X(\u_usb_host.u_core.u_fifo_rx._0535_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0970_  (.A(net252),
    .B(net196),
    .X(\u_usb_host.u_core.u_fifo_rx._0536_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0971_  (.A(net225),
    .B(\u_usb_host.u_core.u_fifo_rx._0522_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0537_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0972_  (.A(net252),
    .B(\u_usb_host.u_core.u_fifo_rx._0526_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0538_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0973_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[32][0] ),
    .B(net229),
    .C(net206),
    .X(\u_usb_host.u_core.u_fifo_rx._0539_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0974_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[59][0] ),
    .B(net236),
    .C(net197),
    .X(\u_usb_host.u_core.u_fifo_rx._0540_ ));
 sky130_fd_sc_hd__and4b_1 \u_usb_host.u_core.u_fifo_rx._0975_  (.A_N(net305),
    .B(net303),
    .C(net301),
    .D(net299),
    .X(\u_usb_host.u_core.u_fifo_rx._0541_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0976_  (.A(net225),
    .B(\u_usb_host.u_core.u_fifo_rx._0518_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0542_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0977_  (.A(net225),
    .B(\u_usb_host.u_core.u_fifo_rx._0526_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0543_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0978_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[51][0] ),
    .B(net235),
    .C(net189),
    .X(\u_usb_host.u_core.u_fifo_rx._0544_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0979_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[49][0] ),
    .B(net230),
    .C(net193),
    .X(\u_usb_host.u_core.u_fifo_rx._0545_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0980_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[8][0] ),
    .B(net226),
    .C(net217),
    .X(\u_usb_host.u_core.u_fifo_rx._0546_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0981_  (.A(net224),
    .B(net191),
    .X(\u_usb_host.u_core.u_fifo_rx._0547_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0982_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[41][0] ),
    .B(net219),
    .C(net202),
    .X(\u_usb_host.u_core.u_fifo_rx._0548_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0983_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[33][0] ),
    .B(net211),
    .C(net195),
    .X(\u_usb_host.u_core.u_fifo_rx._0549_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0984_  (.A(net252),
    .B(net192),
    .X(\u_usb_host.u_core.u_fifo_rx._0550_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0985_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[42][0] ),
    .B(net202),
    .C(net191),
    .X(\u_usb_host.u_core.u_fifo_rx._0551_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0986_  (.A(net259),
    .B(net246),
    .X(\u_usb_host.u_core.u_fifo_rx._0552_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0987_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[63][0] ),
    .B(net258),
    .C(net240),
    .X(\u_usb_host.u_core.u_fifo_rx._0553_ ));
 sky130_fd_sc_hd__and4bb_1 \u_usb_host.u_core.u_fifo_rx._0988_  (.A_N(\u_usb_host.u_core.u_fifo_rx.rd_ptr[0] ),
    .B_N(net304),
    .C(net302),
    .D(net300),
    .X(\u_usb_host.u_core.u_fifo_rx._0554_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0989_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[44][0] ),
    .B(net202),
    .C(net180),
    .X(\u_usb_host.u_core.u_fifo_rx._0555_ ));
 sky130_fd_sc_hd__nor4b_2 \u_usb_host.u_core.u_fifo_rx._0990_  (.A(net305),
    .B(net303),
    .C(net299),
    .D_N(net301),
    .Y(\u_usb_host.u_core.u_fifo_rx._0556_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0991_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[36][0] ),
    .B(net210),
    .C(net177),
    .X(\u_usb_host.u_core.u_fifo_rx._0557_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0992_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[20][0] ),
    .B(net248),
    .C(net179),
    .X(\u_usb_host.u_core.u_fifo_rx._0558_ ));
 sky130_fd_sc_hd__and4b_2 \u_usb_host.u_core.u_fifo_rx._0993_  (.A_N(net303),
    .B(net301),
    .C(net299),
    .D(net306),
    .X(\u_usb_host.u_core.u_fifo_rx._0559_ ));
 sky130_fd_sc_hd__and4bb_2 \u_usb_host.u_core.u_fifo_rx._0994_  (.A_N(net306),
    .B_N(net300),
    .C(net302),
    .D(net304),
    .X(\u_usb_host.u_core.u_fifo_rx._0560_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0995_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[38][0] ),
    .B(net209),
    .C(net172),
    .X(\u_usb_host.u_core.u_fifo_rx._0561_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0996_  (.A(net259),
    .B(net241),
    .X(\u_usb_host.u_core.u_fifo_rx._0562_ ));
 sky130_fd_sc_hd__and4bb_2 \u_usb_host.u_core.u_fifo_rx._0997_  (.A_N(net304),
    .B_N(net300),
    .C(net302),
    .D(net306),
    .X(\u_usb_host.u_core.u_fifo_rx._0563_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0998_  (.A(net226),
    .B(net170),
    .X(\u_usb_host.u_core.u_fifo_rx._0564_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0999_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[14][0] ),
    .B(net222),
    .C(net184),
    .X(\u_usb_host.u_core.u_fifo_rx._0565_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1000_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[15][0] ),
    .B(net255),
    .C(net224),
    .X(\u_usb_host.u_core.u_fifo_rx._0566_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._1001_  (.A(net226),
    .B(net172),
    .X(\u_usb_host.u_core.u_fifo_rx._0567_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._1002_  (.A(net226),
    .B(\u_usb_host.u_core.u_fifo_rx._0556_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0568_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._1003_  (.A(net259),
    .B(net225),
    .X(\u_usb_host.u_core.u_fifo_rx._0569_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1004_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[60][0] ),
    .B(net232),
    .C(net182),
    .X(\u_usb_host.u_core.u_fifo_rx._0570_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1005_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[47][0] ),
    .B(net255),
    .C(net201),
    .X(\u_usb_host.u_core.u_fifo_rx._0571_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1006_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[31][0] ),
    .B(net257),
    .C(net248),
    .X(\u_usb_host.u_core.u_fifo_rx._0572_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1007_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[39][0] ),
    .B(net259),
    .C(net209),
    .X(\u_usb_host.u_core.u_fifo_rx._0573_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1008_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[46][0] ),
    .B(net201),
    .C(net184),
    .X(\u_usb_host.u_core.u_fifo_rx._0574_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1009_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[61][0] ),
    .B(net236),
    .C(net175),
    .X(\u_usb_host.u_core.u_fifo_rx._0575_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1010_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[45][0] ),
    .B(net202),
    .C(net173),
    .X(\u_usb_host.u_core.u_fifo_rx._0576_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._1011_  (.A(net241),
    .B(net172),
    .X(\u_usb_host.u_core.u_fifo_rx._0577_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._1012_  (.A(net235),
    .B(net170),
    .X(\u_usb_host.u_core.u_fifo_rx._0578_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1013_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[52][0] ),
    .B(net241),
    .C(net177),
    .X(\u_usb_host.u_core.u_fifo_rx._0579_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1014_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[21][0] ),
    .B(net253),
    .C(net170),
    .X(\u_usb_host.u_core.u_fifo_rx._0580_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1015_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[28][0] ),
    .B(net250),
    .C(net182),
    .X(\u_usb_host.u_core.u_fifo_rx._0581_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1016_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[62][0] ),
    .B(net240),
    .C(net187),
    .X(\u_usb_host.u_core.u_fifo_rx._0582_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._1017_  (.A(net253),
    .B(net172),
    .X(\u_usb_host.u_core.u_fifo_rx._0583_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1018_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[37][0] ),
    .B(net212),
    .C(net171),
    .X(\u_usb_host.u_core.u_fifo_rx._0584_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1019_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[19][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0538_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0550_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[26][0] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0585_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1020_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[13][0] ),
    .A2(net222),
    .A3(net173),
    .B1(\u_usb_host.u_core.u_fifo_rx._0565_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0545_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0586_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1021_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[5][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0564_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0567_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[6][0] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0587_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1022_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[1][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0543_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[3][0] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0588_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1023_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[27][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0536_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0568_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[4][0] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0587_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0589_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1024_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[2][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0542_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0569_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[7][0] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0588_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0590_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1025_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[25][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0513_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0517_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[24][0] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0585_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0591_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_rx._1026_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[29][0] ),
    .A2(net250),
    .A3(net175),
    .B1(\u_usb_host.u_core.u_fifo_rx._0581_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0592_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1027_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[30][0] ),
    .A2(net250),
    .A3(net187),
    .B1(\u_usb_host.u_core.u_fifo_rx._0592_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0539_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0593_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1028_  (.A(\u_usb_host.u_core.u_fifo_rx._0589_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0590_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0591_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0593_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0594_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1029_  (.A(\u_usb_host.u_core.u_fifo_rx._0534_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0571_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0574_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0576_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0595_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1030_  (.A(\u_usb_host.u_core.u_fifo_rx._0521_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0548_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0551_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0555_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0596_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1031_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[23][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0552_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0535_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0532_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0523_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0597_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1032_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[22][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0583_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0580_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0572_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0558_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0598_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1033_  (.A(\u_usb_host.u_core.u_fifo_rx._0595_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0596_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0597_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0598_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0599_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1034_  (.A(\u_usb_host.u_core.u_fifo_rx._0533_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0546_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0553_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0582_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0600_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1035_  (.A(\u_usb_host.u_core.u_fifo_rx._0525_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0540_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0570_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0575_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0601_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1036_  (.A(\u_usb_host.u_core.u_fifo_rx._0519_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0527_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0549_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0557_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0602_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1037_  (.A(\u_usb_host.u_core.u_fifo_rx._0516_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0561_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0573_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0584_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0603_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1038_  (.A(\u_usb_host.u_core.u_fifo_rx._0600_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0601_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0602_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0603_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0604_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1039_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[55][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0562_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[54][0] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0605_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1040_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[53][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0578_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0579_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0531_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0544_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0606_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1041_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[56][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0530_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0605_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0606_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0510_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0607_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1042_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[9][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0547_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[10][0] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0608_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._1043_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[12][0] ),
    .A2(net223),
    .A3(net181),
    .B1(\u_usb_host.u_core.u_fifo_rx._0529_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[11][0] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0609_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_rx._1044_  (.A(\u_usb_host.u_core.u_fifo_rx._0566_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0586_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0608_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0609_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0610_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1045_  (.A(\u_usb_host.u_core.u_fifo_rx._0599_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0604_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0607_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0610_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0611_ ));
 sky130_fd_sc_hd__o22a_1 \u_usb_host.u_core.u_fifo_rx._1046_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[0][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0511_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0594_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0611_ ),
    .X(\u_usb_host.u_core.u_fifo_rx.data_o[0] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1047_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[40][1] ),
    .B(net218),
    .C(net212),
    .X(\u_usb_host.u_core.u_fifo_rx._0612_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1048_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[33][1] ),
    .B(net211),
    .C(net195),
    .X(\u_usb_host.u_core.u_fifo_rx._0613_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1049_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[43][1] ),
    .B(net207),
    .C(net196),
    .X(\u_usb_host.u_core.u_fifo_rx._0614_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1050_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[17][1] ),
    .B(net244),
    .C(net193),
    .X(\u_usb_host.u_core.u_fifo_rx._0615_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1051_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[59][1] ),
    .B(net232),
    .C(net197),
    .X(\u_usb_host.u_core.u_fifo_rx._0616_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1052_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[35][1] ),
    .B(net214),
    .C(net189),
    .X(\u_usb_host.u_core.u_fifo_rx._0617_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1053_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[50][1] ),
    .B(net234),
    .C(net198),
    .X(\u_usb_host.u_core.u_fifo_rx._0618_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1054_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[16][1] ),
    .B(net245),
    .C(net227),
    .X(\u_usb_host.u_core.u_fifo_rx._0619_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1055_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[57][1] ),
    .B(net238),
    .C(net220),
    .X(\u_usb_host.u_core.u_fifo_rx._0620_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1056_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[48][1] ),
    .B(net230),
    .C(net227),
    .X(\u_usb_host.u_core.u_fifo_rx._0621_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1057_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[18][1] ),
    .B(net247),
    .C(net198),
    .X(\u_usb_host.u_core.u_fifo_rx._0622_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1058_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[32][1] ),
    .B(net229),
    .C(net206),
    .X(\u_usb_host.u_core.u_fifo_rx._0623_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1059_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[58][1] ),
    .B(net236),
    .C(net192),
    .X(\u_usb_host.u_core.u_fifo_rx._0624_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1060_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[51][1] ),
    .B(net234),
    .C(net189),
    .X(\u_usb_host.u_core.u_fifo_rx._0625_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1061_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[49][1] ),
    .B(net230),
    .C(net193),
    .X(\u_usb_host.u_core.u_fifo_rx._0626_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1062_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[8][1] ),
    .B(net225),
    .C(net217),
    .X(\u_usb_host.u_core.u_fifo_rx._0627_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1063_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[41][1] ),
    .B(net219),
    .C(net204),
    .X(\u_usb_host.u_core.u_fifo_rx._0628_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1064_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[34][1] ),
    .B(net210),
    .C(net200),
    .X(\u_usb_host.u_core.u_fifo_rx._0629_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1065_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[42][1] ),
    .B(net204),
    .C(net191),
    .X(\u_usb_host.u_core.u_fifo_rx._0630_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1066_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[63][1] ),
    .B(net258),
    .C(net242),
    .X(\u_usb_host.u_core.u_fifo_rx._0631_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1067_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[44][1] ),
    .B(net204),
    .C(net180),
    .X(\u_usb_host.u_core.u_fifo_rx._0632_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1068_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[36][1] ),
    .B(net211),
    .C(net177),
    .X(\u_usb_host.u_core.u_fifo_rx._0633_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1069_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[20][1] ),
    .B(net247),
    .C(net179),
    .X(\u_usb_host.u_core.u_fifo_rx._0634_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1070_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[38][1] ),
    .B(net212),
    .C(net172),
    .X(\u_usb_host.u_core.u_fifo_rx._0635_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1071_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[14][1] ),
    .B(net221),
    .C(net184),
    .X(\u_usb_host.u_core.u_fifo_rx._0636_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1072_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[15][1] ),
    .B(net255),
    .C(net223),
    .X(\u_usb_host.u_core.u_fifo_rx._0637_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1073_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[60][1] ),
    .B(net232),
    .C(net182),
    .X(\u_usb_host.u_core.u_fifo_rx._0638_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1074_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[47][1] ),
    .B(net255),
    .C(net203),
    .X(\u_usb_host.u_core.u_fifo_rx._0639_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1075_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[31][1] ),
    .B(net256),
    .C(net246),
    .X(\u_usb_host.u_core.u_fifo_rx._0640_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1076_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[39][1] ),
    .B(net259),
    .C(net209),
    .X(\u_usb_host.u_core.u_fifo_rx._0641_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1077_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[46][1] ),
    .B(net203),
    .C(net184),
    .X(\u_usb_host.u_core.u_fifo_rx._0642_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1078_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[61][1] ),
    .B(net233),
    .C(net175),
    .X(\u_usb_host.u_core.u_fifo_rx._0643_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1079_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[45][1] ),
    .B(net201),
    .C(net173),
    .X(\u_usb_host.u_core.u_fifo_rx._0644_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1080_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[52][1] ),
    .B(net241),
    .C(net177),
    .X(\u_usb_host.u_core.u_fifo_rx._0645_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1081_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[21][1] ),
    .B(net253),
    .C(net170),
    .X(\u_usb_host.u_core.u_fifo_rx._0646_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1082_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[28][1] ),
    .B(net250),
    .C(net182),
    .X(\u_usb_host.u_core.u_fifo_rx._0647_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1083_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[62][1] ),
    .B(net239),
    .C(net187),
    .X(\u_usb_host.u_core.u_fifo_rx._0648_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1084_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[37][1] ),
    .B(net212),
    .C(net171),
    .X(\u_usb_host.u_core.u_fifo_rx._0649_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1085_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[19][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0538_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0550_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[26][1] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0650_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1086_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[13][1] ),
    .A2(net221),
    .A3(net173),
    .B1(\u_usb_host.u_core.u_fifo_rx._0626_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0636_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0651_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1087_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[5][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0564_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0567_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[6][1] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0652_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1088_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[1][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0543_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[3][1] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0653_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1089_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[27][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0536_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0568_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[4][1] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0652_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0654_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1090_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[2][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0542_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0569_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[7][1] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0653_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0655_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1091_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[25][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0513_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0517_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[24][1] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0650_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0656_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_rx._1092_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[29][1] ),
    .A2(net250),
    .A3(net176),
    .B1(\u_usb_host.u_core.u_fifo_rx._0647_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0657_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1093_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[30][1] ),
    .A2(net250),
    .A3(net187),
    .B1(\u_usb_host.u_core.u_fifo_rx._0623_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0657_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0658_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1094_  (.A(\u_usb_host.u_core.u_fifo_rx._0654_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0655_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0656_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0658_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0659_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1095_  (.A(\u_usb_host.u_core.u_fifo_rx._0621_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0639_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0642_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0644_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0660_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1096_  (.A(\u_usb_host.u_core.u_fifo_rx._0614_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0628_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0630_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0632_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0661_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1097_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[23][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0552_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0615_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0619_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0622_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0662_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1098_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[22][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0583_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0634_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0640_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0646_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0663_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1099_  (.A(\u_usb_host.u_core.u_fifo_rx._0660_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0661_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0662_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0663_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0664_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1100_  (.A(\u_usb_host.u_core.u_fifo_rx._0620_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0627_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0631_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0648_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0665_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1101_  (.A(\u_usb_host.u_core.u_fifo_rx._0616_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0624_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0638_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0643_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0666_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1102_  (.A(\u_usb_host.u_core.u_fifo_rx._0613_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0617_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0629_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0633_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0667_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1103_  (.A(\u_usb_host.u_core.u_fifo_rx._0612_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0635_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0641_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0649_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0668_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1104_  (.A(\u_usb_host.u_core.u_fifo_rx._0665_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0666_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0667_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0668_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0669_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1105_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[55][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0562_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[54][1] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0670_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1106_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[53][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0578_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0618_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0625_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0645_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0671_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1107_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[56][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0530_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0670_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0671_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0510_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0672_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1108_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[9][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0547_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[10][1] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0673_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._1109_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[12][1] ),
    .A2(net223),
    .A3(net180),
    .B1(\u_usb_host.u_core.u_fifo_rx._0529_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[11][1] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0674_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_rx._1110_  (.A(\u_usb_host.u_core.u_fifo_rx._0637_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0651_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0673_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0674_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0675_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1111_  (.A(\u_usb_host.u_core.u_fifo_rx._0664_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0669_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0672_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0675_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0676_ ));
 sky130_fd_sc_hd__o22a_1 \u_usb_host.u_core.u_fifo_rx._1112_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[0][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0511_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0659_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0676_ ),
    .X(\u_usb_host.u_core.u_fifo_rx.data_o[1] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1113_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[40][2] ),
    .B(net217),
    .C(net213),
    .X(\u_usb_host.u_core.u_fifo_rx._0677_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1114_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[34][2] ),
    .B(net210),
    .C(net200),
    .X(\u_usb_host.u_core.u_fifo_rx._0678_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1115_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[17][2] ),
    .B(net244),
    .C(net194),
    .X(\u_usb_host.u_core.u_fifo_rx._0679_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1116_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[59][2] ),
    .B(net237),
    .C(net197),
    .X(\u_usb_host.u_core.u_fifo_rx._0680_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1117_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[35][2] ),
    .B(net214),
    .C(net190),
    .X(\u_usb_host.u_core.u_fifo_rx._0681_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1118_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[50][2] ),
    .B(net234),
    .C(net199),
    .X(\u_usb_host.u_core.u_fifo_rx._0682_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1119_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[16][2] ),
    .B(net254),
    .C(net228),
    .X(\u_usb_host.u_core.u_fifo_rx._0683_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1120_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[57][2] ),
    .B(net238),
    .C(net220),
    .X(\u_usb_host.u_core.u_fifo_rx._0684_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1121_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[48][2] ),
    .B(net231),
    .C(net227),
    .X(\u_usb_host.u_core.u_fifo_rx._0685_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1122_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[18][2] ),
    .B(net246),
    .C(net198),
    .X(\u_usb_host.u_core.u_fifo_rx._0686_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1123_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[32][2] ),
    .B(net229),
    .C(net206),
    .X(\u_usb_host.u_core.u_fifo_rx._0687_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1124_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[41][2] ),
    .B(net219),
    .C(net206),
    .X(\u_usb_host.u_core.u_fifo_rx._0688_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1125_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[58][2] ),
    .B(net237),
    .C(net192),
    .X(\u_usb_host.u_core.u_fifo_rx._0689_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1126_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[51][2] ),
    .B(net235),
    .C(net189),
    .X(\u_usb_host.u_core.u_fifo_rx._0690_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1127_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[43][2] ),
    .B(net206),
    .C(net196),
    .X(\u_usb_host.u_core.u_fifo_rx._0691_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1128_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[8][2] ),
    .B(net225),
    .C(net217),
    .X(\u_usb_host.u_core.u_fifo_rx._0692_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1129_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[33][2] ),
    .B(net211),
    .C(net195),
    .X(\u_usb_host.u_core.u_fifo_rx._0693_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1130_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[42][2] ),
    .B(net202),
    .C(net191),
    .X(\u_usb_host.u_core.u_fifo_rx._0694_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1131_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[49][2] ),
    .B(net230),
    .C(net193),
    .X(\u_usb_host.u_core.u_fifo_rx._0695_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1132_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[63][2] ),
    .B(net258),
    .C(net242),
    .X(\u_usb_host.u_core.u_fifo_rx._0696_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1133_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[44][2] ),
    .B(net202),
    .C(net180),
    .X(\u_usb_host.u_core.u_fifo_rx._0697_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1134_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[62][2] ),
    .B(net238),
    .C(net187),
    .X(\u_usb_host.u_core.u_fifo_rx._0698_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1135_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[20][2] ),
    .B(net254),
    .C(net179),
    .X(\u_usb_host.u_core.u_fifo_rx._0699_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1136_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[38][2] ),
    .B(net209),
    .C(net172),
    .X(\u_usb_host.u_core.u_fifo_rx._0700_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1137_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[14][2] ),
    .B(net221),
    .C(net184),
    .X(\u_usb_host.u_core.u_fifo_rx._0701_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1138_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[15][2] ),
    .B(net255),
    .C(net223),
    .X(\u_usb_host.u_core.u_fifo_rx._0702_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1139_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[28][2] ),
    .B(net249),
    .C(net182),
    .X(\u_usb_host.u_core.u_fifo_rx._0703_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1140_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[60][2] ),
    .B(net233),
    .C(net183),
    .X(\u_usb_host.u_core.u_fifo_rx._0704_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1141_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[47][2] ),
    .B(net255),
    .C(net201),
    .X(\u_usb_host.u_core.u_fifo_rx._0705_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1142_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[31][2] ),
    .B(net256),
    .C(net248),
    .X(\u_usb_host.u_core.u_fifo_rx._0706_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1143_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[37][2] ),
    .B(net213),
    .C(net171),
    .X(\u_usb_host.u_core.u_fifo_rx._0707_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1144_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[46][2] ),
    .B(net201),
    .C(net185),
    .X(\u_usb_host.u_core.u_fifo_rx._0708_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1145_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[61][2] ),
    .B(net236),
    .C(net175),
    .X(\u_usb_host.u_core.u_fifo_rx._0709_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1146_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[45][2] ),
    .B(net201),
    .C(net174),
    .X(\u_usb_host.u_core.u_fifo_rx._0710_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1147_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[21][2] ),
    .B(net253),
    .C(net170),
    .X(\u_usb_host.u_core.u_fifo_rx._0711_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1148_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[36][2] ),
    .B(net210),
    .C(net178),
    .X(\u_usb_host.u_core.u_fifo_rx._0712_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1149_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[52][2] ),
    .B(net241),
    .C(net177),
    .X(\u_usb_host.u_core.u_fifo_rx._0713_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1150_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[39][2] ),
    .B(net259),
    .C(net209),
    .X(\u_usb_host.u_core.u_fifo_rx._0714_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1151_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[19][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0538_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0550_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[26][2] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0715_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1152_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[13][2] ),
    .A2(net221),
    .A3(net173),
    .B1(\u_usb_host.u_core.u_fifo_rx._0695_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0701_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0086_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1153_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[5][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0564_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0567_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[6][2] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0087_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1154_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[1][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0543_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[3][2] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0088_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1155_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[27][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0536_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0568_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[4][2] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0087_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0089_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1156_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[2][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0542_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0569_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[7][2] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0088_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0090_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1157_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[25][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0513_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0517_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[24][2] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0715_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0091_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_rx._1158_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[29][2] ),
    .A2(net249),
    .A3(net176),
    .B1(\u_usb_host.u_core.u_fifo_rx._0703_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0092_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1159_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[30][2] ),
    .A2(net249),
    .A3(net186),
    .B1(\u_usb_host.u_core.u_fifo_rx._0687_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0092_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0093_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1160_  (.A(\u_usb_host.u_core.u_fifo_rx._0089_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0090_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0091_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0093_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0094_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1161_  (.A(\u_usb_host.u_core.u_fifo_rx._0685_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0705_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0708_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0710_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0095_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1162_  (.A(\u_usb_host.u_core.u_fifo_rx._0688_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0691_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0694_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0697_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0096_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1163_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[23][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0552_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0679_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0683_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0686_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0097_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1164_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[22][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0583_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0699_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0706_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0711_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0098_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1165_  (.A(\u_usb_host.u_core.u_fifo_rx._0095_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0096_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0097_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0098_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0099_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1166_  (.A(\u_usb_host.u_core.u_fifo_rx._0684_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0692_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0696_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0698_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0100_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1167_  (.A(\u_usb_host.u_core.u_fifo_rx._0680_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0689_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0704_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0709_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0101_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1168_  (.A(\u_usb_host.u_core.u_fifo_rx._0678_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0681_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0693_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0712_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0102_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1169_  (.A(\u_usb_host.u_core.u_fifo_rx._0677_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0700_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0707_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0714_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0103_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1170_  (.A(\u_usb_host.u_core.u_fifo_rx._0100_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0101_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0102_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0103_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0104_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1171_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[55][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0562_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[54][2] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0105_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1172_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[53][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0578_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0682_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0690_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0713_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0106_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1173_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[56][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0530_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0105_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0106_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0510_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0107_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1174_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[9][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0547_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[10][2] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0108_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._1175_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[12][2] ),
    .A2(net223),
    .A3(net181),
    .B1(\u_usb_host.u_core.u_fifo_rx._0529_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[11][2] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0109_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_rx._1176_  (.A(\u_usb_host.u_core.u_fifo_rx._0702_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0086_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0108_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0109_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0110_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1177_  (.A(\u_usb_host.u_core.u_fifo_rx._0099_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0104_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0107_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0110_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0111_ ));
 sky130_fd_sc_hd__o22a_1 \u_usb_host.u_core.u_fifo_rx._1178_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[0][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0511_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0094_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0111_ ),
    .X(\u_usb_host.u_core.u_fifo_rx.data_o[2] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1179_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[40][3] ),
    .B(net218),
    .C(net213),
    .X(\u_usb_host.u_core.u_fifo_rx._0112_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1180_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[33][3] ),
    .B(net211),
    .C(net195),
    .X(\u_usb_host.u_core.u_fifo_rx._0113_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1181_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[43][3] ),
    .B(net208),
    .C(net196),
    .X(\u_usb_host.u_core.u_fifo_rx._0114_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1182_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[17][3] ),
    .B(net244),
    .C(net194),
    .X(\u_usb_host.u_core.u_fifo_rx._0115_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1183_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[59][3] ),
    .B(net237),
    .C(net197),
    .X(\u_usb_host.u_core.u_fifo_rx._0116_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1184_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[35][3] ),
    .B(net214),
    .C(net190),
    .X(\u_usb_host.u_core.u_fifo_rx._0117_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1185_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[50][3] ),
    .B(net234),
    .C(net199),
    .X(\u_usb_host.u_core.u_fifo_rx._0118_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1186_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[16][3] ),
    .B(net245),
    .C(net228),
    .X(\u_usb_host.u_core.u_fifo_rx._0119_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1187_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[57][3] ),
    .B(net238),
    .C(net220),
    .X(\u_usb_host.u_core.u_fifo_rx._0120_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1188_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[48][3] ),
    .B(net231),
    .C(net227),
    .X(\u_usb_host.u_core.u_fifo_rx._0121_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1189_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[18][3] ),
    .B(net246),
    .C(net198),
    .X(\u_usb_host.u_core.u_fifo_rx._0122_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1190_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[32][3] ),
    .B(net229),
    .C(net206),
    .X(\u_usb_host.u_core.u_fifo_rx._0123_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1191_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[58][3] ),
    .B(net236),
    .C(net192),
    .X(\u_usb_host.u_core.u_fifo_rx._0124_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1192_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[51][3] ),
    .B(net235),
    .C(net189),
    .X(\u_usb_host.u_core.u_fifo_rx._0125_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1193_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[49][3] ),
    .B(net230),
    .C(net193),
    .X(\u_usb_host.u_core.u_fifo_rx._0126_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1194_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[8][3] ),
    .B(net225),
    .C(net217),
    .X(\u_usb_host.u_core.u_fifo_rx._0127_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1195_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[41][3] ),
    .B(net219),
    .C(net204),
    .X(\u_usb_host.u_core.u_fifo_rx._0128_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1196_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[34][3] ),
    .B(net216),
    .C(net200),
    .X(\u_usb_host.u_core.u_fifo_rx._0129_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1197_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[42][3] ),
    .B(net204),
    .C(net191),
    .X(\u_usb_host.u_core.u_fifo_rx._0130_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1198_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[63][3] ),
    .B(net258),
    .C(net238),
    .X(\u_usb_host.u_core.u_fifo_rx._0131_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1199_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[44][3] ),
    .B(net205),
    .C(net180),
    .X(\u_usb_host.u_core.u_fifo_rx._0132_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1200_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[36][3] ),
    .B(net216),
    .C(net178),
    .X(\u_usb_host.u_core.u_fifo_rx._0133_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1201_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[20][3] ),
    .B(net247),
    .C(net179),
    .X(\u_usb_host.u_core.u_fifo_rx._0134_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1202_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[38][3] ),
    .B(net213),
    .C(net172),
    .X(\u_usb_host.u_core.u_fifo_rx._0135_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1203_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[14][3] ),
    .B(net221),
    .C(net184),
    .X(\u_usb_host.u_core.u_fifo_rx._0136_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1204_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[15][3] ),
    .B(net255),
    .C(net223),
    .X(\u_usb_host.u_core.u_fifo_rx._0137_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1205_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[60][3] ),
    .B(net232),
    .C(net183),
    .X(\u_usb_host.u_core.u_fifo_rx._0138_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1206_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[47][3] ),
    .B(net255),
    .C(net203),
    .X(\u_usb_host.u_core.u_fifo_rx._0139_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1207_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[31][3] ),
    .B(net257),
    .C(net246),
    .X(\u_usb_host.u_core.u_fifo_rx._0140_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1208_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[39][3] ),
    .B(net259),
    .C(net209),
    .X(\u_usb_host.u_core.u_fifo_rx._0141_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1209_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[46][3] ),
    .B(net203),
    .C(net185),
    .X(\u_usb_host.u_core.u_fifo_rx._0142_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1210_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[61][3] ),
    .B(net236),
    .C(net175),
    .X(\u_usb_host.u_core.u_fifo_rx._0143_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1211_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[45][3] ),
    .B(net201),
    .C(net174),
    .X(\u_usb_host.u_core.u_fifo_rx._0144_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1212_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[52][3] ),
    .B(net241),
    .C(net177),
    .X(\u_usb_host.u_core.u_fifo_rx._0145_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1213_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[21][3] ),
    .B(net253),
    .C(net170),
    .X(\u_usb_host.u_core.u_fifo_rx._0146_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1214_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[28][3] ),
    .B(net249),
    .C(net182),
    .X(\u_usb_host.u_core.u_fifo_rx._0147_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1215_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[62][3] ),
    .B(net238),
    .C(net187),
    .X(\u_usb_host.u_core.u_fifo_rx._0148_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1216_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[37][3] ),
    .B(net213),
    .C(net171),
    .X(\u_usb_host.u_core.u_fifo_rx._0149_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1217_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[19][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0538_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0550_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[26][3] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0150_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1218_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[13][3] ),
    .A2(net221),
    .A3(net173),
    .B1(\u_usb_host.u_core.u_fifo_rx._0126_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0136_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0151_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1219_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[5][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0564_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0567_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[6][3] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0152_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1220_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[1][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0543_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[3][3] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0153_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1221_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[27][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0536_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0568_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[4][3] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0152_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0154_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1222_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[2][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0542_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0569_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[7][3] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0153_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0155_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1223_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[25][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0513_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0517_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[24][3] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0150_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0156_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_rx._1224_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[29][3] ),
    .A2(net249),
    .A3(net176),
    .B1(\u_usb_host.u_core.u_fifo_rx._0147_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0157_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1225_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[30][3] ),
    .A2(net249),
    .A3(net186),
    .B1(\u_usb_host.u_core.u_fifo_rx._0123_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0157_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0158_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1226_  (.A(\u_usb_host.u_core.u_fifo_rx._0154_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0155_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0156_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0158_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0159_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1227_  (.A(\u_usb_host.u_core.u_fifo_rx._0121_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0139_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0142_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0144_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0160_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1228_  (.A(\u_usb_host.u_core.u_fifo_rx._0114_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0128_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0130_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0132_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0161_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1229_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[23][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0552_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0115_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0119_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0122_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0162_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1230_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[22][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0583_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0134_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0140_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0146_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0163_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_rx._1231_  (.A(\u_usb_host.u_core.u_fifo_rx._0160_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0161_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0162_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0163_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0164_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1232_  (.A(\u_usb_host.u_core.u_fifo_rx._0120_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0127_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0131_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0148_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0165_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1233_  (.A(\u_usb_host.u_core.u_fifo_rx._0116_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0124_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0138_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0143_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0166_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1234_  (.A(\u_usb_host.u_core.u_fifo_rx._0113_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0117_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0129_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0133_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0167_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1235_  (.A(\u_usb_host.u_core.u_fifo_rx._0112_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0135_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0141_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0149_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0168_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1236_  (.A(\u_usb_host.u_core.u_fifo_rx._0165_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0166_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0167_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0168_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0169_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1237_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[55][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0562_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[54][3] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0170_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1238_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[53][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0578_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0118_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0125_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0145_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0171_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1239_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[56][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0530_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0170_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0171_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0510_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0172_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1240_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[9][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0547_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[10][3] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0173_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._1241_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[12][3] ),
    .A2(net224),
    .A3(net181),
    .B1(\u_usb_host.u_core.u_fifo_rx._0529_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[11][3] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0174_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_rx._1242_  (.A(\u_usb_host.u_core.u_fifo_rx._0137_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0151_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0173_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0174_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0175_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1243_  (.A(\u_usb_host.u_core.u_fifo_rx._0164_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0169_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0172_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0175_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0176_ ));
 sky130_fd_sc_hd__o22a_1 \u_usb_host.u_core.u_fifo_rx._1244_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[0][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0511_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0159_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0176_ ),
    .X(\u_usb_host.u_core.u_fifo_rx.data_o[3] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1245_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[40][4] ),
    .B(net218),
    .C(net213),
    .X(\u_usb_host.u_core.u_fifo_rx._0177_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1246_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[33][4] ),
    .B(net211),
    .C(net195),
    .X(\u_usb_host.u_core.u_fifo_rx._0178_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1247_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[43][4] ),
    .B(net207),
    .C(net196),
    .X(\u_usb_host.u_core.u_fifo_rx._0179_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1248_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[17][4] ),
    .B(net244),
    .C(net194),
    .X(\u_usb_host.u_core.u_fifo_rx._0180_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1249_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[59][4] ),
    .B(net233),
    .C(net197),
    .X(\u_usb_host.u_core.u_fifo_rx._0181_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1250_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[35][4] ),
    .B(net214),
    .C(net190),
    .X(\u_usb_host.u_core.u_fifo_rx._0182_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1251_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[50][4] ),
    .B(net234),
    .C(net199),
    .X(\u_usb_host.u_core.u_fifo_rx._0183_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1252_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[16][4] ),
    .B(net245),
    .C(net228),
    .X(\u_usb_host.u_core.u_fifo_rx._0184_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1253_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[57][4] ),
    .B(net238),
    .C(net220),
    .X(\u_usb_host.u_core.u_fifo_rx._0185_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1254_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[48][4] ),
    .B(net231),
    .C(net227),
    .X(\u_usb_host.u_core.u_fifo_rx._0186_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1255_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[18][4] ),
    .B(net247),
    .C(net198),
    .X(\u_usb_host.u_core.u_fifo_rx._0187_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1256_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[32][4] ),
    .B(net229),
    .C(net206),
    .X(\u_usb_host.u_core.u_fifo_rx._0188_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1257_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[58][4] ),
    .B(net237),
    .C(net192),
    .X(\u_usb_host.u_core.u_fifo_rx._0189_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1258_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[51][4] ),
    .B(net234),
    .C(net189),
    .X(\u_usb_host.u_core.u_fifo_rx._0190_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1259_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[49][4] ),
    .B(net230),
    .C(net193),
    .X(\u_usb_host.u_core.u_fifo_rx._0191_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1260_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[8][4] ),
    .B(net225),
    .C(net217),
    .X(\u_usb_host.u_core.u_fifo_rx._0192_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1261_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[41][4] ),
    .B(net219),
    .C(net207),
    .X(\u_usb_host.u_core.u_fifo_rx._0193_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1262_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[34][4] ),
    .B(net216),
    .C(net200),
    .X(\u_usb_host.u_core.u_fifo_rx._0194_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1263_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[42][4] ),
    .B(net208),
    .C(net191),
    .X(\u_usb_host.u_core.u_fifo_rx._0195_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1264_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[63][4] ),
    .B(net258),
    .C(net238),
    .X(\u_usb_host.u_core.u_fifo_rx._0196_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1265_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[44][4] ),
    .B(net204),
    .C(net180),
    .X(\u_usb_host.u_core.u_fifo_rx._0197_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1266_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[36][4] ),
    .B(net216),
    .C(net178),
    .X(\u_usb_host.u_core.u_fifo_rx._0198_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1267_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[20][4] ),
    .B(net247),
    .C(net179),
    .X(\u_usb_host.u_core.u_fifo_rx._0199_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1268_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[38][4] ),
    .B(net215),
    .C(net172),
    .X(\u_usb_host.u_core.u_fifo_rx._0200_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1269_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[14][4] ),
    .B(net221),
    .C(net184),
    .X(\u_usb_host.u_core.u_fifo_rx._0201_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1270_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[15][4] ),
    .B(net255),
    .C(net223),
    .X(\u_usb_host.u_core.u_fifo_rx._0202_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1271_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[60][4] ),
    .B(net232),
    .C(net183),
    .X(\u_usb_host.u_core.u_fifo_rx._0203_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1272_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[47][4] ),
    .B(net257),
    .C(net205),
    .X(\u_usb_host.u_core.u_fifo_rx._0204_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1273_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[31][4] ),
    .B(net257),
    .C(net246),
    .X(\u_usb_host.u_core.u_fifo_rx._0205_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1274_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[39][4] ),
    .B(net259),
    .C(net209),
    .X(\u_usb_host.u_core.u_fifo_rx._0206_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1275_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[46][4] ),
    .B(net205),
    .C(net185),
    .X(\u_usb_host.u_core.u_fifo_rx._0207_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1276_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[61][4] ),
    .B(net233),
    .C(net175),
    .X(\u_usb_host.u_core.u_fifo_rx._0208_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1277_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[45][4] ),
    .B(net202),
    .C(net174),
    .X(\u_usb_host.u_core.u_fifo_rx._0209_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1278_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[52][4] ),
    .B(net241),
    .C(net177),
    .X(\u_usb_host.u_core.u_fifo_rx._0210_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1279_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[21][4] ),
    .B(net253),
    .C(net170),
    .X(\u_usb_host.u_core.u_fifo_rx._0211_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1280_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[28][4] ),
    .B(net249),
    .C(net182),
    .X(\u_usb_host.u_core.u_fifo_rx._0212_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1281_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[62][4] ),
    .B(net238),
    .C(net187),
    .X(\u_usb_host.u_core.u_fifo_rx._0213_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1282_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[37][4] ),
    .B(net213),
    .C(net171),
    .X(\u_usb_host.u_core.u_fifo_rx._0214_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1283_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[19][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0538_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0550_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[26][4] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0215_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1284_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[13][4] ),
    .A2(net221),
    .A3(net173),
    .B1(\u_usb_host.u_core.u_fifo_rx._0191_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0201_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0216_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1285_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[5][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0564_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0567_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[6][4] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0217_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1286_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[1][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0543_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[3][4] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0218_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1287_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[27][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0536_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0568_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[4][4] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0217_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0219_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1288_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[2][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0542_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0569_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[7][4] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0218_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0220_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1289_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[25][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0513_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0517_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[24][4] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0215_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0221_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_rx._1290_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[29][4] ),
    .A2(net249),
    .A3(net176),
    .B1(\u_usb_host.u_core.u_fifo_rx._0212_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0222_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1291_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[30][4] ),
    .A2(net249),
    .A3(net186),
    .B1(\u_usb_host.u_core.u_fifo_rx._0188_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0222_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0223_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1292_  (.A(\u_usb_host.u_core.u_fifo_rx._0219_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0220_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0221_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0223_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0224_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1293_  (.A(\u_usb_host.u_core.u_fifo_rx._0186_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0204_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0207_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0209_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0225_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1294_  (.A(\u_usb_host.u_core.u_fifo_rx._0179_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0193_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0195_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0197_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0226_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1295_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[23][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0552_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0180_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0184_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0187_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0227_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1296_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[22][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0583_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0199_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0205_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0211_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0228_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1297_  (.A(\u_usb_host.u_core.u_fifo_rx._0225_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0226_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0227_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0228_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0229_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1298_  (.A(\u_usb_host.u_core.u_fifo_rx._0185_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0192_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0196_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0213_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0230_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1299_  (.A(\u_usb_host.u_core.u_fifo_rx._0181_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0189_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0203_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0208_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0231_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1300_  (.A(\u_usb_host.u_core.u_fifo_rx._0178_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0182_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0194_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0198_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0232_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1301_  (.A(\u_usb_host.u_core.u_fifo_rx._0177_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0200_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0206_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0214_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0233_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1302_  (.A(\u_usb_host.u_core.u_fifo_rx._0230_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0231_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0232_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0233_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0234_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1303_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[55][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0562_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[54][4] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0235_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1304_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[53][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0578_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0183_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0190_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0210_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0236_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1305_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[56][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0530_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0235_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0236_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0510_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0237_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1306_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[9][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0547_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[10][4] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0238_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._1307_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[12][4] ),
    .A2(net223),
    .A3(net180),
    .B1(\u_usb_host.u_core.u_fifo_rx._0529_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[11][4] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0239_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_rx._1308_  (.A(\u_usb_host.u_core.u_fifo_rx._0202_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0216_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0238_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0239_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0240_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1309_  (.A(\u_usb_host.u_core.u_fifo_rx._0229_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0234_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0237_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0240_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0241_ ));
 sky130_fd_sc_hd__o22a_1 \u_usb_host.u_core.u_fifo_rx._1310_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[0][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0511_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0224_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0241_ ),
    .X(\u_usb_host.u_core.u_fifo_rx.data_o[4] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1311_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[34][5] ),
    .B(net210),
    .C(net200),
    .X(\u_usb_host.u_core.u_fifo_rx._0242_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1312_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[58][5] ),
    .B(net237),
    .C(net192),
    .X(\u_usb_host.u_core.u_fifo_rx._0243_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1313_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[43][5] ),
    .B(net207),
    .C(net196),
    .X(\u_usb_host.u_core.u_fifo_rx._0244_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1314_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[8][5] ),
    .B(net225),
    .C(net217),
    .X(\u_usb_host.u_core.u_fifo_rx._0245_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1315_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[17][5] ),
    .B(net245),
    .C(net194),
    .X(\u_usb_host.u_core.u_fifo_rx._0246_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1316_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[40][5] ),
    .B(net218),
    .C(net212),
    .X(\u_usb_host.u_core.u_fifo_rx._0247_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1317_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[50][5] ),
    .B(net234),
    .C(net199),
    .X(\u_usb_host.u_core.u_fifo_rx._0248_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1318_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[16][5] ),
    .B(net245),
    .C(net228),
    .X(\u_usb_host.u_core.u_fifo_rx._0249_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1319_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[57][5] ),
    .B(net239),
    .C(net220),
    .X(\u_usb_host.u_core.u_fifo_rx._0250_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1320_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[48][5] ),
    .B(net231),
    .C(net227),
    .X(\u_usb_host.u_core.u_fifo_rx._0251_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1321_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[18][5] ),
    .B(net246),
    .C(net198),
    .X(\u_usb_host.u_core.u_fifo_rx._0252_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1322_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[41][5] ),
    .B(net219),
    .C(net207),
    .X(\u_usb_host.u_core.u_fifo_rx._0253_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1323_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[35][5] ),
    .B(net214),
    .C(net190),
    .X(\u_usb_host.u_core.u_fifo_rx._0254_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1324_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[59][5] ),
    .B(net236),
    .C(net197),
    .X(\u_usb_host.u_core.u_fifo_rx._0255_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1325_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[46][5] ),
    .B(net203),
    .C(net185),
    .X(\u_usb_host.u_core.u_fifo_rx._0256_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1326_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[51][5] ),
    .B(net235),
    .C(net189),
    .X(\u_usb_host.u_core.u_fifo_rx._0257_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1327_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[42][5] ),
    .B(net208),
    .C(net191),
    .X(\u_usb_host.u_core.u_fifo_rx._0258_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1328_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[33][5] ),
    .B(net211),
    .C(net195),
    .X(\u_usb_host.u_core.u_fifo_rx._0259_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1329_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[32][5] ),
    .B(net229),
    .C(net207),
    .X(\u_usb_host.u_core.u_fifo_rx._0260_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1330_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[49][5] ),
    .B(net230),
    .C(net193),
    .X(\u_usb_host.u_core.u_fifo_rx._0261_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1331_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[36][5] ),
    .B(net210),
    .C(net178),
    .X(\u_usb_host.u_core.u_fifo_rx._0262_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1332_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[63][5] ),
    .B(net258),
    .C(net240),
    .X(\u_usb_host.u_core.u_fifo_rx._0263_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1333_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[20][5] ),
    .B(net247),
    .C(net179),
    .X(\u_usb_host.u_core.u_fifo_rx._0264_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1334_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[31][5] ),
    .B(net256),
    .C(net247),
    .X(\u_usb_host.u_core.u_fifo_rx._0265_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1335_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[44][5] ),
    .B(net204),
    .C(net180),
    .X(\u_usb_host.u_core.u_fifo_rx._0266_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1336_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[14][5] ),
    .B(net222),
    .C(net184),
    .X(\u_usb_host.u_core.u_fifo_rx._0267_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1337_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[15][5] ),
    .B(net256),
    .C(net224),
    .X(\u_usb_host.u_core.u_fifo_rx._0268_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1338_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[5][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0564_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0567_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[6][5] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0269_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1339_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[60][5] ),
    .B(net232),
    .C(net183),
    .X(\u_usb_host.u_core.u_fifo_rx._0270_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1340_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[47][5] ),
    .B(net257),
    .C(net203),
    .X(\u_usb_host.u_core.u_fifo_rx._0271_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1341_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[39][5] ),
    .B(net259),
    .C(net209),
    .X(\u_usb_host.u_core.u_fifo_rx._0272_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1342_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[61][5] ),
    .B(net236),
    .C(net175),
    .X(\u_usb_host.u_core.u_fifo_rx._0273_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1343_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[45][5] ),
    .B(net201),
    .C(net174),
    .X(\u_usb_host.u_core.u_fifo_rx._0274_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1344_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[38][5] ),
    .B(net212),
    .C(net172),
    .X(\u_usb_host.u_core.u_fifo_rx._0275_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1345_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[62][5] ),
    .B(net240),
    .C(net188),
    .X(\u_usb_host.u_core.u_fifo_rx._0276_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1346_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[52][5] ),
    .B(net241),
    .C(net177),
    .X(\u_usb_host.u_core.u_fifo_rx._0277_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1347_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[28][5] ),
    .B(net250),
    .C(net182),
    .X(\u_usb_host.u_core.u_fifo_rx._0278_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1348_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[21][5] ),
    .B(net253),
    .C(net170),
    .X(\u_usb_host.u_core.u_fifo_rx._0279_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1349_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[37][5] ),
    .B(net212),
    .C(net171),
    .X(\u_usb_host.u_core.u_fifo_rx._0280_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1350_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[19][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0538_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0550_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[26][5] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0281_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1351_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[13][5] ),
    .A2(net222),
    .A3(net173),
    .B1(\u_usb_host.u_core.u_fifo_rx._0261_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0267_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0282_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1352_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[1][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0543_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[3][5] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0283_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1353_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[27][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0536_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0568_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[4][5] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0269_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0284_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1354_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[2][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0542_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0569_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[7][5] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0283_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0285_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1355_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[25][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0513_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0517_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[24][5] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0281_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0286_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_rx._1356_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[29][5] ),
    .A2(net250),
    .A3(net176),
    .B1(\u_usb_host.u_core.u_fifo_rx._0278_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0287_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1357_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[30][5] ),
    .A2(net250),
    .A3(net187),
    .B1(\u_usb_host.u_core.u_fifo_rx._0260_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0287_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0288_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1358_  (.A(\u_usb_host.u_core.u_fifo_rx._0284_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0285_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0286_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0288_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0289_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1359_  (.A(\u_usb_host.u_core.u_fifo_rx._0251_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0256_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0271_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0274_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0290_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1360_  (.A(\u_usb_host.u_core.u_fifo_rx._0244_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0253_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0258_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0266_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0291_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1361_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[23][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0552_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0246_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0249_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0252_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0292_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1362_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[22][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0583_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0264_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0265_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0279_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0293_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1363_  (.A(\u_usb_host.u_core.u_fifo_rx._0290_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0291_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0292_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0293_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0294_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1364_  (.A(\u_usb_host.u_core.u_fifo_rx._0245_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0250_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0263_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0276_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0295_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1365_  (.A(\u_usb_host.u_core.u_fifo_rx._0243_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0255_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0270_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0273_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0296_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1366_  (.A(\u_usb_host.u_core.u_fifo_rx._0242_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0254_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0259_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0262_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0297_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1367_  (.A(\u_usb_host.u_core.u_fifo_rx._0247_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0272_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0275_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0280_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0298_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1368_  (.A(\u_usb_host.u_core.u_fifo_rx._0295_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0296_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0297_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0298_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0299_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1369_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[55][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0562_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[54][5] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0300_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1370_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[53][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0578_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0248_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0257_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0277_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0301_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1371_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[56][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0530_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0300_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0301_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0510_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0302_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1372_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[9][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0547_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[10][5] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0303_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._1373_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[12][5] ),
    .A2(net224),
    .A3(net181),
    .B1(\u_usb_host.u_core.u_fifo_rx._0529_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[11][5] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0304_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_rx._1374_  (.A(\u_usb_host.u_core.u_fifo_rx._0268_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0282_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0303_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0304_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0305_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1375_  (.A(\u_usb_host.u_core.u_fifo_rx._0294_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0299_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0302_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0305_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0306_ ));
 sky130_fd_sc_hd__o22a_1 \u_usb_host.u_core.u_fifo_rx._1376_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[0][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0511_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0289_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0306_ ),
    .X(\u_usb_host.u_core.u_fifo_rx.data_o[5] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1377_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[40][6] ),
    .B(net218),
    .C(net213),
    .X(\u_usb_host.u_core.u_fifo_rx._0307_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1378_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[34][6] ),
    .B(net210),
    .C(net200),
    .X(\u_usb_host.u_core.u_fifo_rx._0308_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1379_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[43][6] ),
    .B(net207),
    .C(net196),
    .X(\u_usb_host.u_core.u_fifo_rx._0309_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1380_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[17][6] ),
    .B(net244),
    .C(net194),
    .X(\u_usb_host.u_core.u_fifo_rx._0310_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1381_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[58][6] ),
    .B(net237),
    .C(net192),
    .X(\u_usb_host.u_core.u_fifo_rx._0311_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1382_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[35][6] ),
    .B(net214),
    .C(net190),
    .X(\u_usb_host.u_core.u_fifo_rx._0312_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1383_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[50][6] ),
    .B(net234),
    .C(net199),
    .X(\u_usb_host.u_core.u_fifo_rx._0313_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1384_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[16][6] ),
    .B(net244),
    .C(net228),
    .X(\u_usb_host.u_core.u_fifo_rx._0314_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1385_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[57][6] ),
    .B(net238),
    .C(net220),
    .X(\u_usb_host.u_core.u_fifo_rx._0315_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1386_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[48][6] ),
    .B(net231),
    .C(net227),
    .X(\u_usb_host.u_core.u_fifo_rx._0316_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1387_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[18][6] ),
    .B(net246),
    .C(net198),
    .X(\u_usb_host.u_core.u_fifo_rx._0317_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1388_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[32][6] ),
    .B(\u_usb_host.u_core.u_fifo_rx._0508_ ),
    .C(net207),
    .X(\u_usb_host.u_core.u_fifo_rx._0318_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1389_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[59][6] ),
    .B(net232),
    .C(net197),
    .X(\u_usb_host.u_core.u_fifo_rx._0319_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1390_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[51][6] ),
    .B(net235),
    .C(net189),
    .X(\u_usb_host.u_core.u_fifo_rx._0320_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1391_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[49][6] ),
    .B(net230),
    .C(net193),
    .X(\u_usb_host.u_core.u_fifo_rx._0321_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1392_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[8][6] ),
    .B(net225),
    .C(net217),
    .X(\u_usb_host.u_core.u_fifo_rx._0322_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1393_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[41][6] ),
    .B(net219),
    .C(net204),
    .X(\u_usb_host.u_core.u_fifo_rx._0323_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1394_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[33][6] ),
    .B(net211),
    .C(net195),
    .X(\u_usb_host.u_core.u_fifo_rx._0324_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1395_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[42][6] ),
    .B(net204),
    .C(net191),
    .X(\u_usb_host.u_core.u_fifo_rx._0325_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1396_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[63][6] ),
    .B(net258),
    .C(net242),
    .X(\u_usb_host.u_core.u_fifo_rx._0326_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1397_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[44][6] ),
    .B(net204),
    .C(net180),
    .X(\u_usb_host.u_core.u_fifo_rx._0327_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1398_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[62][6] ),
    .B(net239),
    .C(net188),
    .X(\u_usb_host.u_core.u_fifo_rx._0328_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1399_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[20][6] ),
    .B(net247),
    .C(net179),
    .X(\u_usb_host.u_core.u_fifo_rx._0329_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1400_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[38][6] ),
    .B(net213),
    .C(net172),
    .X(\u_usb_host.u_core.u_fifo_rx._0330_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1401_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[14][6] ),
    .B(net221),
    .C(net184),
    .X(\u_usb_host.u_core.u_fifo_rx._0331_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1402_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[15][6] ),
    .B(net256),
    .C(net224),
    .X(\u_usb_host.u_core.u_fifo_rx._0332_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1403_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[28][6] ),
    .B(net251),
    .C(net182),
    .X(\u_usb_host.u_core.u_fifo_rx._0333_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1404_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[60][6] ),
    .B(net232),
    .C(net183),
    .X(\u_usb_host.u_core.u_fifo_rx._0334_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1405_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[47][6] ),
    .B(net257),
    .C(net203),
    .X(\u_usb_host.u_core.u_fifo_rx._0335_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1406_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[31][6] ),
    .B(net256),
    .C(net247),
    .X(\u_usb_host.u_core.u_fifo_rx._0336_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1407_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[37][6] ),
    .B(net213),
    .C(net171),
    .X(\u_usb_host.u_core.u_fifo_rx._0337_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1408_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[46][6] ),
    .B(net203),
    .C(net185),
    .X(\u_usb_host.u_core.u_fifo_rx._0338_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1409_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[61][6] ),
    .B(net232),
    .C(net175),
    .X(\u_usb_host.u_core.u_fifo_rx._0339_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1410_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[45][6] ),
    .B(net201),
    .C(net174),
    .X(\u_usb_host.u_core.u_fifo_rx._0340_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1411_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[21][6] ),
    .B(net253),
    .C(net170),
    .X(\u_usb_host.u_core.u_fifo_rx._0341_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1412_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[36][6] ),
    .B(net211),
    .C(net178),
    .X(\u_usb_host.u_core.u_fifo_rx._0342_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1413_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[52][6] ),
    .B(net241),
    .C(net177),
    .X(\u_usb_host.u_core.u_fifo_rx._0343_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1414_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[39][6] ),
    .B(\u_usb_host.u_core.u_fifo_rx._0497_ ),
    .C(net215),
    .X(\u_usb_host.u_core.u_fifo_rx._0344_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1415_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[19][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0538_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0550_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[26][6] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0345_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1416_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[13][6] ),
    .A2(net221),
    .A3(net173),
    .B1(\u_usb_host.u_core.u_fifo_rx._0321_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0331_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0346_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1417_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[5][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0564_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0567_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[6][6] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0347_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1418_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[1][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0543_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[3][6] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0348_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1419_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[27][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0536_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0568_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[4][6] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0347_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0349_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1420_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[2][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0542_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0569_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[7][6] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0348_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0350_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1421_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[25][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0513_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0517_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[24][6] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0345_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0351_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_rx._1422_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[29][6] ),
    .A2(net251),
    .A3(net175),
    .B1(\u_usb_host.u_core.u_fifo_rx._0333_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0352_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1423_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[30][6] ),
    .A2(net251),
    .A3(net187),
    .B1(\u_usb_host.u_core.u_fifo_rx._0318_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0352_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0353_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1424_  (.A(\u_usb_host.u_core.u_fifo_rx._0349_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0350_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0351_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0353_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0354_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1425_  (.A(\u_usb_host.u_core.u_fifo_rx._0316_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0335_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0338_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0340_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0355_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1426_  (.A(\u_usb_host.u_core.u_fifo_rx._0309_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0323_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0325_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0327_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0356_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1427_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[23][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0552_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0310_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0314_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0317_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0357_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1428_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[22][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0583_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0329_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0336_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0341_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0358_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1429_  (.A(\u_usb_host.u_core.u_fifo_rx._0355_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0356_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0357_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0358_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0359_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1430_  (.A(\u_usb_host.u_core.u_fifo_rx._0315_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0322_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0326_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0328_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0360_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1431_  (.A(\u_usb_host.u_core.u_fifo_rx._0311_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0319_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0334_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0339_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0361_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1432_  (.A(\u_usb_host.u_core.u_fifo_rx._0308_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0312_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0324_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0342_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0362_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1433_  (.A(\u_usb_host.u_core.u_fifo_rx._0307_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0330_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0337_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0344_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0363_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1434_  (.A(\u_usb_host.u_core.u_fifo_rx._0360_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0361_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0362_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0363_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0364_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1435_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[55][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0562_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[54][6] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0365_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1436_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[53][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0578_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0313_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0320_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0343_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0366_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1437_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[56][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0530_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0365_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0366_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0510_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0367_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1438_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[9][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0547_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[10][6] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0368_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._1439_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[12][6] ),
    .A2(net224),
    .A3(net181),
    .B1(\u_usb_host.u_core.u_fifo_rx._0529_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[11][6] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0369_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_rx._1440_  (.A(\u_usb_host.u_core.u_fifo_rx._0332_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0346_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0368_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0369_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0370_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1441_  (.A(\u_usb_host.u_core.u_fifo_rx._0359_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0364_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0367_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0370_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0371_ ));
 sky130_fd_sc_hd__o22a_1 \u_usb_host.u_core.u_fifo_rx._1442_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[0][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0511_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0354_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0371_ ),
    .X(\u_usb_host.u_core.u_fifo_rx.data_o[6] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1443_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[34][7] ),
    .B(net210),
    .C(net200),
    .X(\u_usb_host.u_core.u_fifo_rx._0372_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1444_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[58][7] ),
    .B(net237),
    .C(net192),
    .X(\u_usb_host.u_core.u_fifo_rx._0373_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1445_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[42][7] ),
    .B(net202),
    .C(net191),
    .X(\u_usb_host.u_core.u_fifo_rx._0374_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1446_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[43][7] ),
    .B(net206),
    .C(net196),
    .X(\u_usb_host.u_core.u_fifo_rx._0375_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1447_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[8][7] ),
    .B(net226),
    .C(net217),
    .X(\u_usb_host.u_core.u_fifo_rx._0376_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1448_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[40][7] ),
    .B(net218),
    .C(net212),
    .X(\u_usb_host.u_core.u_fifo_rx._0377_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1449_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[50][7] ),
    .B(net234),
    .C(net199),
    .X(\u_usb_host.u_core.u_fifo_rx._0378_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1450_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[16][7] ),
    .B(net244),
    .C(net228),
    .X(\u_usb_host.u_core.u_fifo_rx._0379_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1451_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[57][7] ),
    .B(net239),
    .C(net220),
    .X(\u_usb_host.u_core.u_fifo_rx._0380_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1452_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[48][7] ),
    .B(net231),
    .C(net227),
    .X(\u_usb_host.u_core.u_fifo_rx._0381_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1453_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[18][7] ),
    .B(net246),
    .C(net198),
    .X(\u_usb_host.u_core.u_fifo_rx._0382_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1454_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[17][7] ),
    .B(net244),
    .C(net194),
    .X(\u_usb_host.u_core.u_fifo_rx._0383_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1455_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[35][7] ),
    .B(net214),
    .C(net190),
    .X(\u_usb_host.u_core.u_fifo_rx._0384_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1456_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[59][7] ),
    .B(net236),
    .C(net197),
    .X(\u_usb_host.u_core.u_fifo_rx._0385_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1457_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[46][7] ),
    .B(net203),
    .C(net185),
    .X(\u_usb_host.u_core.u_fifo_rx._0386_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1458_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[51][7] ),
    .B(net235),
    .C(net189),
    .X(\u_usb_host.u_core.u_fifo_rx._0387_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1459_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[49][7] ),
    .B(net230),
    .C(net193),
    .X(\u_usb_host.u_core.u_fifo_rx._0388_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1460_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[41][7] ),
    .B(net219),
    .C(net206),
    .X(\u_usb_host.u_core.u_fifo_rx._0389_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1461_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[33][7] ),
    .B(net211),
    .C(net195),
    .X(\u_usb_host.u_core.u_fifo_rx._0390_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1462_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[32][7] ),
    .B(\u_usb_host.u_core.u_fifo_rx._0508_ ),
    .C(net207),
    .X(\u_usb_host.u_core.u_fifo_rx._0391_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1463_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[36][7] ),
    .B(net210),
    .C(net178),
    .X(\u_usb_host.u_core.u_fifo_rx._0392_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1464_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[63][7] ),
    .B(net258),
    .C(net242),
    .X(\u_usb_host.u_core.u_fifo_rx._0393_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1465_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[20][7] ),
    .B(net248),
    .C(net179),
    .X(\u_usb_host.u_core.u_fifo_rx._0394_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1466_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[13][7] ),
    .B(net222),
    .C(net173),
    .X(\u_usb_host.u_core.u_fifo_rx._0395_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1467_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[31][7] ),
    .B(net257),
    .C(net248),
    .X(\u_usb_host.u_core.u_fifo_rx._0396_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1468_  (.A(\u_usb_host.u_core.u_fifo_rx._0716_ ),
    .B(net202),
    .C(net180),
    .X(\u_usb_host.u_core.u_fifo_rx._0397_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1469_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[14][7] ),
    .B(net222),
    .C(net184),
    .X(\u_usb_host.u_core.u_fifo_rx._0398_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1470_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[15][7] ),
    .B(net255),
    .C(net222),
    .X(\u_usb_host.u_core.u_fifo_rx._0399_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1471_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[5][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0564_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0567_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[6][7] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0400_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1472_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[60][7] ),
    .B(net232),
    .C(net183),
    .X(\u_usb_host.u_core.u_fifo_rx._0401_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1473_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[47][7] ),
    .B(net257),
    .C(net203),
    .X(\u_usb_host.u_core.u_fifo_rx._0402_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1474_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[39][7] ),
    .B(\u_usb_host.u_core.u_fifo_rx._0497_ ),
    .C(net209),
    .X(\u_usb_host.u_core.u_fifo_rx._0403_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1475_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[61][7] ),
    .B(net236),
    .C(net176),
    .X(\u_usb_host.u_core.u_fifo_rx._0404_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1476_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[45][7] ),
    .B(net201),
    .C(net174),
    .X(\u_usb_host.u_core.u_fifo_rx._0405_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1477_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[38][7] ),
    .B(net209),
    .C(\u_usb_host.u_core.u_fifo_rx._0560_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0406_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1478_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[62][7] ),
    .B(net239),
    .C(net188),
    .X(\u_usb_host.u_core.u_fifo_rx._0407_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1479_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[52][7] ),
    .B(net241),
    .C(net177),
    .X(\u_usb_host.u_core.u_fifo_rx._0408_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1480_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[28][7] ),
    .B(net251),
    .C(net182),
    .X(\u_usb_host.u_core.u_fifo_rx._0409_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1481_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[21][7] ),
    .B(net253),
    .C(net170),
    .X(\u_usb_host.u_core.u_fifo_rx._0410_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1482_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[37][7] ),
    .B(net212),
    .C(net171),
    .X(\u_usb_host.u_core.u_fifo_rx._0411_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1483_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[19][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0538_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0550_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[26][7] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0412_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1484_  (.A(\u_usb_host.u_core.u_fifo_rx._0388_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0395_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0398_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0399_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0413_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1485_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[1][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0543_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[3][7] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0414_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1486_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[27][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0536_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0568_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[4][7] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0400_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0415_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1487_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[2][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0542_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0569_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[7][7] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0414_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0416_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1488_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[25][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0513_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0517_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[24][7] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0412_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0417_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_rx._1489_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[29][7] ),
    .A2(net250),
    .A3(net175),
    .B1(\u_usb_host.u_core.u_fifo_rx._0409_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0418_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1490_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[30][7] ),
    .A2(net251),
    .A3(net187),
    .B1(\u_usb_host.u_core.u_fifo_rx._0391_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0418_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0419_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1491_  (.A(\u_usb_host.u_core.u_fifo_rx._0415_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0416_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0417_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0419_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0420_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1492_  (.A(\u_usb_host.u_core.u_fifo_rx._0381_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0386_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0402_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0405_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0421_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1493_  (.A(\u_usb_host.u_core.u_fifo_rx._0374_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0375_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0389_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0397_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0422_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1494_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[23][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0552_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0379_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0382_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0383_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0423_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1495_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[22][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0583_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0394_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0396_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0410_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0424_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1496_  (.A(\u_usb_host.u_core.u_fifo_rx._0421_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0422_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0423_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0424_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0425_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1497_  (.A(\u_usb_host.u_core.u_fifo_rx._0376_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0380_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0393_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0407_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0426_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1498_  (.A(\u_usb_host.u_core.u_fifo_rx._0373_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0385_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0401_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0404_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0427_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1499_  (.A(\u_usb_host.u_core.u_fifo_rx._0372_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0384_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0390_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0392_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0428_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1500_  (.A(\u_usb_host.u_core.u_fifo_rx._0377_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0403_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0406_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0411_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0429_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1501_  (.A(\u_usb_host.u_core.u_fifo_rx._0426_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0427_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0428_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0429_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0430_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1502_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[55][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0562_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[54][7] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0431_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1503_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[53][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0578_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0378_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0387_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0408_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0432_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1504_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[56][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0530_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0431_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0432_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0510_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0433_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1505_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[9][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0547_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[10][7] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0434_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._1506_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[12][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0509_ ),
    .A3(net181),
    .B1(\u_usb_host.u_core.u_fifo_rx._0529_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[11][7] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0435_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_core.u_fifo_rx._1507_  (.A(\u_usb_host.u_core.u_fifo_rx._0413_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0434_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0435_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0436_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1508_  (.A(\u_usb_host.u_core.u_fifo_rx._0425_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0430_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0433_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0436_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0437_ ));
 sky130_fd_sc_hd__o22a_1 \u_usb_host.u_core.u_fifo_rx._1509_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[0][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0511_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0420_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0437_ ),
    .X(\u_usb_host.u_core.u_fifo_rx.data_o[7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1510_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ),
    .D(net165),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1511_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ),
    .D(net156),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1512_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ),
    .D(net150),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1513_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ),
    .D(net142),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1514_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ),
    .D(net133),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1515_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ),
    .D(net125),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1516_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ),
    .D(net116),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1517_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ),
    .D(net107),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1518_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ),
    .D(net166),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[58][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1519_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ),
    .D(net157),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[58][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1520_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ),
    .D(net149),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[58][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1521_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ),
    .D(net142),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[58][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1522_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ),
    .D(net133),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[58][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1523_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ),
    .D(net126),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[58][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1524_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ),
    .D(net117),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[58][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1525_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ),
    .D(net108),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[58][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1526_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ),
    .D(net165),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1527_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ),
    .D(net159),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1528_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ),
    .D(net151),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1529_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ),
    .D(net143),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1530_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ),
    .D(net135),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1531_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ),
    .D(net125),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1532_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ),
    .D(net116),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1533_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ),
    .D(net110),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1534_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ),
    .D(net165),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1535_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ),
    .D(net159),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1536_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ),
    .D(net151),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1537_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ),
    .D(net143),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1538_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ),
    .D(net133),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1539_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ),
    .D(net125),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1540_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ),
    .D(net116),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1541_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ),
    .D(net110),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1542_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ),
    .D(net167),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[57][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1543_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ),
    .D(net158),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[57][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1544_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ),
    .D(net149),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[57][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1545_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ),
    .D(net141),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[57][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1546_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ),
    .D(net134),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[57][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1547_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ),
    .D(net127),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[57][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1548_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ),
    .D(net118),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[57][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1549_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ),
    .D(net109),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[57][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1550_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ),
    .D(net165),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1551_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ),
    .D(net159),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1552_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ),
    .D(net151),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1553_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ),
    .D(net143),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1554_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ),
    .D(net133),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1555_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ),
    .D(net125),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1556_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ),
    .D(net116),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1557_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ),
    .D(net110),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1558_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ),
    .D(net166),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[56][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1559_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ),
    .D(net156),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[56][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1560_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ),
    .D(net149),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[56][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1561_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ),
    .D(net141),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[56][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1562_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ),
    .D(net134),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[56][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1563_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ),
    .D(net126),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[56][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1564_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ),
    .D(net117),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[56][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1565_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ),
    .D(net108),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[56][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1566_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ),
    .D(net163),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1567_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ),
    .D(net155),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1568_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ),
    .D(net147),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1569_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ),
    .D(net137),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1570_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ),
    .D(net129),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1571_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ),
    .D(net121),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1572_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ),
    .D(net112),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1573_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ),
    .D(net105),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1574_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ),
    .D(net164),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1575_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ),
    .D(net155),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1576_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ),
    .D(net147),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1577_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ),
    .D(net139),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1578_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ),
    .D(net131),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1579_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ),
    .D(net123),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1580_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ),
    .D(net114),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1581_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ),
    .D(net106),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1582_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ),
    .D(net166),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[55][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1583_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ),
    .D(net158),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[55][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1584_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ),
    .D(net149),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[55][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1585_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ),
    .D(net141),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[55][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1586_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ),
    .D(net134),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[55][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1587_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ),
    .D(net128),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[55][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1588_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ),
    .D(net117),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[55][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1589_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ),
    .D(net109),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[55][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1590_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ),
    .D(net164),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1591_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ),
    .D(net156),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1592_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ),
    .D(net147),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1593_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ),
    .D(net139),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1594_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ),
    .D(net131),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1595_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ),
    .D(net123),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1596_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ),
    .D(net115),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1597_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ),
    .D(net106),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1598_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ),
    .D(net166),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[54][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1599_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ),
    .D(net157),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[54][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1600_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ),
    .D(net149),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[54][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1601_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ),
    .D(net141),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[54][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1602_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ),
    .D(net134),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[54][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1603_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ),
    .D(net126),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[54][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1604_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ),
    .D(net117),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[54][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1605_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ),
    .D(net108),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[54][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1606_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ),
    .D(net164),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1607_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ),
    .D(net155),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1608_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ),
    .D(net147),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1609_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ),
    .D(net139),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1610_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ),
    .D(net131),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1611_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ),
    .D(net123),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1612_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ),
    .D(net115),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1613_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ),
    .D(net106),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1614_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ),
    .D(net165),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1615_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ),
    .D(net159),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1616_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ),
    .D(net151),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1617_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ),
    .D(net143),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1618_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ),
    .D(net135),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1619_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ),
    .D(net125),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1620_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ),
    .D(net116),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1621_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ),
    .D(net110),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1622_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ),
    .D(net166),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[53][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1623_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ),
    .D(net156),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[53][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1624_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ),
    .D(net149),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[53][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1625_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ),
    .D(net141),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[53][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1626_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ),
    .D(net134),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[53][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1627_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ),
    .D(net126),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[53][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1628_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ),
    .D(net117),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[53][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1629_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ),
    .D(net108),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[53][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1630_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ),
    .D(net164),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1631_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ),
    .D(net155),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1632_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ),
    .D(net148),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1633_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ),
    .D(net140),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1634_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ),
    .D(net132),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1635_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ),
    .D(net124),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1636_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ),
    .D(net115),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1637_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ),
    .D(net106),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1638_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ),
    .D(net166),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[52][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1639_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ),
    .D(net156),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[52][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1640_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ),
    .D(net149),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[52][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1641_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ),
    .D(net142),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[52][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1642_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ),
    .D(net136),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[52][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1643_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ),
    .D(net126),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[52][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1644_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ),
    .D(net117),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[52][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1645_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ),
    .D(net108),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[52][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1646_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ),
    .D(net163),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1647_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ),
    .D(net153),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1648_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ),
    .D(net145),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1649_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ),
    .D(net138),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1650_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ),
    .D(net130),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1651_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ),
    .D(net122),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1652_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ),
    .D(net112),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1653_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ),
    .D(net105),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1654_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ),
    .D(net163),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1655_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ),
    .D(net154),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1656_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ),
    .D(net146),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1657_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ),
    .D(net138),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1658_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ),
    .D(net130),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1659_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ),
    .D(net122),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1660_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ),
    .D(net112),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1661_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ),
    .D(net105),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1662_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ),
    .D(net166),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[51][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1663_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ),
    .D(net157),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[51][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1664_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ),
    .D(net149),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[51][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1665_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ),
    .D(net141),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[51][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1666_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ),
    .D(net134),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[51][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1667_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ),
    .D(net126),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[51][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1668_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ),
    .D(net117),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[51][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1669_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ),
    .D(net108),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[51][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1670_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ),
    .D(net162),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1671_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ),
    .D(net153),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1672_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ),
    .D(net145),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1673_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ),
    .D(net137),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1674_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ),
    .D(net129),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1675_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ),
    .D(net121),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1676_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ),
    .D(net112),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1677_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ),
    .D(net104),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1678_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ),
    .D(net164),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[50][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1679_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ),
    .D(net157),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[50][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1680_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ),
    .D(net148),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[50][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1681_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ),
    .D(net140),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[50][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1682_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ),
    .D(net132),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[50][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1683_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ),
    .D(net124),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[50][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1684_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ),
    .D(net114),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[50][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1685_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ),
    .D(net106),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[50][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1686_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ),
    .D(net162),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1687_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ),
    .D(net153),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1688_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ),
    .D(net145),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1689_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ),
    .D(net137),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1690_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ),
    .D(net129),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1691_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ),
    .D(net121),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1692_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ),
    .D(net112),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1693_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ),
    .D(net104),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1694_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ),
    .D(net162),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1695_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ),
    .D(net153),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1696_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ),
    .D(net145),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1697_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ),
    .D(net137),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1698_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ),
    .D(net129),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1699_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ),
    .D(net121),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1700_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ),
    .D(net112),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1701_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ),
    .D(net104),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1702_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ),
    .D(net162),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[49][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1703_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ),
    .D(net153),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[49][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1704_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ),
    .D(net145),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[49][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1705_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ),
    .D(net137),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[49][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1706_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ),
    .D(net129),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[49][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1707_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ),
    .D(net121),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[49][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1708_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ),
    .D(net112),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[49][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1709_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ),
    .D(net104),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[49][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1710_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ),
    .D(net162),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1711_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ),
    .D(net153),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1712_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ),
    .D(net145),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1713_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ),
    .D(net137),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1714_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ),
    .D(net129),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1715_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ),
    .D(net121),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1716_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ),
    .D(net114),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1717_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ),
    .D(net104),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1718_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ),
    .D(net162),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[48][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1719_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ),
    .D(net154),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[48][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1720_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ),
    .D(net146),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[48][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1721_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ),
    .D(net138),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[48][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1722_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ),
    .D(net130),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[48][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1723_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ),
    .D(net122),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[48][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1724_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ),
    .D(net112),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[48][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1725_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ),
    .D(net104),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[48][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1726_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ),
    .D(net162),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1727_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ),
    .D(net153),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1728_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ),
    .D(net145),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1729_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ),
    .D(net137),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1730_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ),
    .D(net129),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1731_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ),
    .D(net121),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1732_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ),
    .D(net114),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1733_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ),
    .D(net104),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1734_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ),
    .D(net162),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1735_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ),
    .D(net153),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1736_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ),
    .D(net145),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1737_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ),
    .D(net137),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1738_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ),
    .D(net129),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1739_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ),
    .D(net121),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1740_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ),
    .D(net112),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1741_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ),
    .D(net104),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1742_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ),
    .D(net162),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[47][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1743_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ),
    .D(net154),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[47][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1744_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ),
    .D(net146),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[47][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1745_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ),
    .D(net138),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[47][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1746_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ),
    .D(net130),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[47][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1747_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ),
    .D(net122),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[47][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1748_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ),
    .D(net113),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[47][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1749_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ),
    .D(net104),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[47][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1750_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ),
    .D(net162),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1751_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ),
    .D(net153),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1752_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ),
    .D(net145),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1753_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ),
    .D(net137),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1754_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ),
    .D(net129),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1755_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ),
    .D(net121),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1756_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ),
    .D(net114),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1757_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ),
    .D(net104),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1758_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ),
    .D(net163),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[46][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1759_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ),
    .D(net154),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[46][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1760_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ),
    .D(net146),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[46][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1761_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ),
    .D(net138),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[46][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1762_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ),
    .D(net130),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[46][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1763_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ),
    .D(net122),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[46][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1764_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ),
    .D(net113),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[46][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1765_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ),
    .D(net105),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[46][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1766_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ),
    .D(net168),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1767_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ),
    .D(net158),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1768_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ),
    .D(net152),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1769_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ),
    .D(net144),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1770_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ),
    .D(net135),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1771_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ),
    .D(net127),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1772_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ),
    .D(net118),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1773_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ),
    .D(net111),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1774_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ),
    .D(net167),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1775_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ),
    .D(net159),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1776_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ),
    .D(net151),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1777_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ),
    .D(net143),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1778_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ),
    .D(net135),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1779_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ),
    .D(net127),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1780_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ),
    .D(net119),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1781_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ),
    .D(net110),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1782_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ),
    .D(net163),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[45][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1783_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ),
    .D(net153),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[45][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1784_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ),
    .D(net146),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[45][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1785_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ),
    .D(net137),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[45][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1786_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ),
    .D(net129),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[45][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1787_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ),
    .D(net121),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[45][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1788_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ),
    .D(net113),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[45][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1789_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ),
    .D(net105),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[45][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1790_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ),
    .D(net165),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1791_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ),
    .D(net156),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1792_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ),
    .D(net150),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1793_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ),
    .D(net142),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1794_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ),
    .D(net133),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1795_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ),
    .D(net125),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1796_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ),
    .D(net116),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1797_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ),
    .D(net107),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1798_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ),
    .D(net163),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[44][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1799_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ),
    .D(net154),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[44][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1800_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ),
    .D(net146),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[44][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1801_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ),
    .D(net138),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[44][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1802_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ),
    .D(net130),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[44][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1803_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ),
    .D(net122),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[44][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1804_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ),
    .D(net113),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[44][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1805_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ),
    .D(net105),
    .Q(\u_usb_host.u_core.u_fifo_rx._0716_ ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1806_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ),
    .D(net165),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1807_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ),
    .D(net156),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1808_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ),
    .D(net150),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1809_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ),
    .D(net142),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1810_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ),
    .D(net133),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1811_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ),
    .D(net125),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1812_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ),
    .D(net116),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1813_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ),
    .D(net107),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1814_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ),
    .D(net165),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1815_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ),
    .D(net156),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1816_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ),
    .D(net150),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1817_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ),
    .D(net142),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1818_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ),
    .D(net133),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1819_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ),
    .D(net125),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1820_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ),
    .D(net116),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1821_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ),
    .D(net107),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1822_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ),
    .D(net169),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[43][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1823_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ),
    .D(net155),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[43][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1824_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ),
    .D(net148),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[43][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1825_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ),
    .D(net139),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[43][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1826_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ),
    .D(net131),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[43][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1827_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ),
    .D(net123),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[43][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1828_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ),
    .D(net114),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[43][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1829_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ),
    .D(net106),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[43][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1830_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ),
    .D(net167),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1831_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ),
    .D(net159),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1832_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ),
    .D(net151),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1833_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ),
    .D(net143),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1834_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ),
    .D(net135),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1835_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ),
    .D(net127),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1836_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ),
    .D(net119),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1837_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ),
    .D(net110),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1838_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ),
    .D(net163),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[42][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1839_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ),
    .D(net154),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[42][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1840_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ),
    .D(net145),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[42][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1841_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ),
    .D(net138),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[42][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1842_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ),
    .D(net130),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[42][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1843_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ),
    .D(net122),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[42][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1844_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ),
    .D(net113),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[42][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1845_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ),
    .D(net105),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[42][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1846_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ),
    .D(net167),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1847_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ),
    .D(net159),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1848_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ),
    .D(net151),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1849_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ),
    .D(net143),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1850_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ),
    .D(net135),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1851_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ),
    .D(net127),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1852_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ),
    .D(net119),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1853_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ),
    .D(net110),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1854_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ),
    .D(net163),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[41][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1855_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ),
    .D(net161),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[41][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1856_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ),
    .D(net148),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[41][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1857_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ),
    .D(net138),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[41][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1858_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ),
    .D(net130),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[41][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1859_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ),
    .D(net122),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[41][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1860_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ),
    .D(net112),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[41][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1861_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ),
    .D(net105),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[41][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1862_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ),
    .D(net167),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1863_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ),
    .D(net159),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1864_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ),
    .D(net151),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1865_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ),
    .D(net143),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1866_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ),
    .D(net135),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1867_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ),
    .D(net127),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1868_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ),
    .D(net119),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1869_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ),
    .D(net110),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1870_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ),
    .D(net167),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[40][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1871_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ),
    .D(net158),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[40][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1872_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ),
    .D(net151),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[40][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1873_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ),
    .D(net143),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[40][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1874_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ),
    .D(net135),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[40][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1875_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ),
    .D(net127),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[40][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1876_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ),
    .D(net118),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[40][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1877_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ),
    .D(net109),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[40][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1878_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ),
    .D(net165),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1879_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ),
    .D(net156),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1880_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ),
    .D(net150),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1881_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ),
    .D(net142),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1882_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ),
    .D(net133),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1883_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ),
    .D(net125),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1884_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ),
    .D(net116),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1885_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ),
    .D(net107),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1886_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ),
    .D(net168),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[39][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1887_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ),
    .D(net159),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[39][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1888_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ),
    .D(net151),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[39][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1889_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ),
    .D(net143),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[39][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1890_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ),
    .D(net135),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[39][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1891_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ),
    .D(net127),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[39][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1892_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ),
    .D(net119),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[39][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1893_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ),
    .D(net111),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[39][7] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_fifo_rx._1894_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0000_ ),
    .RESET_B(net267),
    .Q(\u_usb_host.u_core.u_fifo_rx.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_fifo_rx._1895_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0001_ ),
    .RESET_B(net267),
    .Q(\u_usb_host.u_core.u_fifo_rx.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1896_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0002_ ),
    .RESET_B(net267),
    .Q(\u_usb_host.u_core.u_fifo_rx.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1897_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0003_ ),
    .RESET_B(net268),
    .Q(\u_usb_host.u_core.u_fifo_rx.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1898_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0004_ ),
    .RESET_B(net270),
    .Q(\u_usb_host.u_core.u_fifo_rx.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1899_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0005_ ),
    .RESET_B(net270),
    .Q(\u_usb_host.u_core.u_fifo_rx.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1900_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0006_ ),
    .RESET_B(net270),
    .Q(\u_usb_host.u_core.u_fifo_rx.count[6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1901_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ),
    .D(net167),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[38][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1902_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ),
    .D(net158),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[38][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1903_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ),
    .D(net152),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[38][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1904_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ),
    .D(net144),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[38][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1905_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ),
    .D(net136),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[38][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1906_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ),
    .D(net128),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[38][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1907_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ),
    .D(net119),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[38][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1908_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ),
    .D(net110),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[38][7] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1909_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0007_ ),
    .RESET_B(net269),
    .Q(\u_usb_host.u_core.u_fifo_rx.rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1910_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0008_ ),
    .RESET_B(net269),
    .Q(\u_usb_host.u_core.u_fifo_rx.rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1911_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0009_ ),
    .RESET_B(net269),
    .Q(\u_usb_host.u_core.u_fifo_rx.rd_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1912_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0010_ ),
    .RESET_B(net269),
    .Q(\u_usb_host.u_core.u_fifo_rx.rd_ptr[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1913_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0011_ ),
    .RESET_B(net269),
    .Q(\u_usb_host.u_core.u_fifo_rx.rd_ptr[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1914_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0012_ ),
    .RESET_B(net269),
    .Q(\u_usb_host.u_core.u_fifo_rx.rd_ptr[5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1915_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ),
    .D(net168),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[37][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1916_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ),
    .D(net158),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[37][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1917_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ),
    .D(net152),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[37][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1918_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ),
    .D(net144),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[37][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1919_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ),
    .D(net136),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[37][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1920_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ),
    .D(net128),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[37][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1921_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ),
    .D(net118),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[37][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1922_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ),
    .D(net109),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[37][7] ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1923_  (.CLK(clknet_4_15_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0019_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0717_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1924_  (.CLK(clknet_4_12_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0020_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0718_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1925_  (.CLK(clknet_4_14_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0021_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0719_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1926_  (.CLK(clknet_4_12_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0022_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0720_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1927_  (.CLK(clknet_4_7_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0023_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0721_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1928_  (.CLK(clknet_4_7_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0024_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0722_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1929_  (.CLK(clknet_4_7_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0025_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0723_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1930_  (.CLK(clknet_4_12_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0026_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0724_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1931_  (.CLK(clknet_4_14_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0027_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0725_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1932_  (.CLK(clknet_4_14_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0028_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0726_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1933_  (.CLK(clknet_4_14_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0029_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0727_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1934_  (.CLK(clknet_4_12_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0030_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0728_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1935_  (.CLK(clknet_4_9_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0031_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0729_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1936_  (.CLK(clknet_4_9_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0032_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0730_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1937_  (.CLK(clknet_4_14_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0033_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0731_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1938_  (.CLK(clknet_4_14_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0034_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0732_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1939_  (.CLK(clknet_4_7_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0035_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0733_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1940_  (.CLK(clknet_4_4_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0036_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0734_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1941_  (.CLK(clknet_4_7_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0037_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0735_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1942_  (.CLK(clknet_4_5_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0038_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0736_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1943_  (.CLK(clknet_4_4_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0039_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0737_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1944_  (.CLK(clknet_4_4_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0040_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0738_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1945_  (.CLK(clknet_4_4_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0041_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0739_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1946_  (.CLK(clknet_4_5_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0042_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0740_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1947_  (.CLK(clknet_4_5_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0043_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0741_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1948_  (.CLK(clknet_4_5_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0044_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0742_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1949_  (.CLK(clknet_4_14_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0045_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0743_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1950_  (.CLK(clknet_4_13_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0046_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0744_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1951_  (.CLK(clknet_4_13_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0047_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0745_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1952_  (.CLK(clknet_4_13_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0048_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0746_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1953_  (.CLK(clknet_4_5_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0049_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0747_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1954_  (.CLK(clknet_4_14_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0050_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0748_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1955_  (.CLK(clknet_4_14_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0051_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0749_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1956_  (.CLK(clknet_4_9_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0052_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0750_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1957_  (.CLK(clknet_4_12_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0053_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0751_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1958_  (.CLK(clknet_4_6_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0054_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0752_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1959_  (.CLK(clknet_4_6_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0055_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0753_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1960_  (.CLK(clknet_4_7_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0056_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0754_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1961_  (.CLK(clknet_4_5_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0057_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0755_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1962_  (.CLK(clknet_4_12_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0058_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0756_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1963_  (.CLK(clknet_4_15_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0059_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0757_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1964_  (.CLK(clknet_4_15_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0060_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0758_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1965_  (.CLK(clknet_4_15_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0061_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0759_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1966_  (.CLK(clknet_4_15_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0062_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0760_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1967_  (.CLK(clknet_4_15_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0063_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0761_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1968_  (.CLK(clknet_4_15_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0064_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0762_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1969_  (.CLK(clknet_4_14_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0065_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0763_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1970_  (.CLK(clknet_4_15_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0066_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0764_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1971_  (.CLK(clknet_4_5_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0067_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0765_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1972_  (.CLK(clknet_4_5_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0068_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0766_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1973_  (.CLK(clknet_4_5_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0069_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0767_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1974_  (.CLK(clknet_4_5_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0070_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0768_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1975_  (.CLK(clknet_4_4_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0071_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0769_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1976_  (.CLK(clknet_4_4_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0072_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0770_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1977_  (.CLK(clknet_4_4_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0073_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0771_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1978_  (.CLK(clknet_4_5_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0074_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0772_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1979_  (.CLK(clknet_4_4_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0075_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0773_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1980_  (.CLK(clknet_4_13_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0076_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0774_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1981_  (.CLK(clknet_4_13_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0077_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0775_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1982_  (.CLK(clknet_4_15_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0078_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0776_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1983_  (.CLK(clknet_4_13_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0079_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0777_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1984_  (.CLK(clknet_4_13_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0080_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0778_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1985_  (.CLK(clknet_4_15_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0081_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0779_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1986_  (.CLK(clknet_4_13_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0082_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0780_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1987_  (.CLK(clknet_4_15_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0083_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0781_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1988_  (.CLK(clknet_4_12_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0084_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0782_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1989_  (.CLK(clknet_4_12_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0085_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0783_ ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1990_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0717_ ),
    .D(net167),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[63][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1991_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0717_ ),
    .D(net160),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[63][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1992_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0717_ ),
    .D(net149),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[63][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1993_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0717_ ),
    .D(net141),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[63][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1994_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0717_ ),
    .D(net133),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[63][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1995_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0717_ ),
    .D(net127),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[63][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1996_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0717_ ),
    .D(net118),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[63][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1997_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0717_ ),
    .D(net109),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[63][7] ));
 sky130_fd_sc_hd__dfrtp_4 \u_usb_host.u_core.u_fifo_rx._1998_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0013_ ),
    .RESET_B(net269),
    .Q(\u_usb_host.u_core.u_fifo_rx.wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_4 \u_usb_host.u_core.u_fifo_rx._1999_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0014_ ),
    .RESET_B(net279),
    .Q(\u_usb_host.u_core.u_fifo_rx.wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._2000_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0015_ ),
    .RESET_B(net269),
    .Q(\u_usb_host.u_core.u_fifo_rx.wr_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._2001_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0016_ ),
    .RESET_B(net269),
    .Q(\u_usb_host.u_core.u_fifo_rx.wr_ptr[3] ));
 sky130_fd_sc_hd__dfrtp_4 \u_usb_host.u_core.u_fifo_rx._2002_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0017_ ),
    .RESET_B(net279),
    .Q(\u_usb_host.u_core.u_fifo_rx.wr_ptr[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._2003_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0018_ ),
    .RESET_B(net271),
    .Q(\u_usb_host.u_core.u_fifo_rx.wr_ptr[5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2004_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0719_ ),
    .D(net167),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[62][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2005_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0719_ ),
    .D(net158),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[62][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2006_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0719_ ),
    .D(net150),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[62][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2007_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0719_ ),
    .D(net141),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[62][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2008_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0719_ ),
    .D(net134),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[62][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2009_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0719_ ),
    .D(net127),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[62][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2010_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0719_ ),
    .D(net118),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[62][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2011_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0719_ ),
    .D(net109),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[62][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2012_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0720_ ),
    .D(net166),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[60][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2013_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0720_ ),
    .D(net157),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[60][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2014_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0720_ ),
    .D(net147),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[60][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2015_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0720_ ),
    .D(net139),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[60][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2016_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0720_ ),
    .D(net131),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[60][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2017_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0720_ ),
    .D(net123),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[60][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2018_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0720_ ),
    .D(net115),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[60][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2019_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0720_ ),
    .D(net108),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[60][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2020_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ),
    .D(net166),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[59][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2021_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ),
    .D(net157),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[59][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2022_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ),
    .D(net149),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[59][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2023_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ),
    .D(net141),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[59][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2024_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ),
    .D(net136),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[59][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2025_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ),
    .D(net126),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[59][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2026_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ),
    .D(net117),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[59][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2027_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ),
    .D(net108),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[59][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2028_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ),
    .D(net168),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[36][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2029_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ),
    .D(net160),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[36][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2030_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ),
    .D(net152),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[36][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2031_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ),
    .D(net142),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[36][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2032_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ),
    .D(net134),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[36][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2033_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ),
    .D(net128),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[36][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2034_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ),
    .D(net118),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[36][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2035_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ),
    .D(net109),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[36][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2036_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ),
    .D(net164),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2037_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ),
    .D(net155),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2038_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ),
    .D(net147),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2039_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ),
    .D(net139),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2040_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ),
    .D(net131),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2041_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ),
    .D(net123),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2042_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ),
    .D(net114),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2043_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ),
    .D(net107),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2044_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ),
    .D(net164),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2045_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ),
    .D(net155),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2046_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ),
    .D(net147),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2047_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ),
    .D(net139),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2048_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ),
    .D(net131),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2049_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ),
    .D(net123),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2050_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ),
    .D(net114),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2051_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ),
    .D(net107),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2052_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ),
    .D(net164),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2053_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ),
    .D(net155),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2054_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ),
    .D(net147),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2055_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ),
    .D(net139),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2056_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ),
    .D(net131),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2057_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ),
    .D(net123),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2058_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ),
    .D(net114),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2059_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ),
    .D(net107),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2060_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ),
    .D(net164),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2061_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ),
    .D(net155),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2062_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ),
    .D(net147),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2063_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ),
    .D(net139),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2064_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ),
    .D(net131),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2065_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ),
    .D(net123),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2066_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ),
    .D(net115),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2067_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ),
    .D(net106),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2068_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ),
    .D(net164),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[32][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2069_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ),
    .D(net155),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[32][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2070_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ),
    .D(net147),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[32][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2071_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ),
    .D(net139),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[32][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2072_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ),
    .D(net131),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[32][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2073_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ),
    .D(net123),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[32][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2074_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ),
    .D(net114),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[32][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2075_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ),
    .D(net107),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[32][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2076_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ),
    .D(net168),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[33][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2077_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ),
    .D(net158),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[33][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2078_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ),
    .D(net152),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[33][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2079_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ),
    .D(net144),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[33][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2080_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ),
    .D(net135),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[33][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2081_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ),
    .D(net128),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[33][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2082_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ),
    .D(net118),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[33][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2083_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ),
    .D(net109),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[33][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2084_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ),
    .D(net167),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[34][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2085_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ),
    .D(net158),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[34][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2086_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ),
    .D(net152),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[34][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2087_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ),
    .D(net141),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[34][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2088_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ),
    .D(net134),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[34][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2089_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ),
    .D(net128),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[34][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2090_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ),
    .D(net118),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[34][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2091_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ),
    .D(net109),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[34][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2092_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ),
    .D(net168),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[35][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2093_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ),
    .D(net158),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[35][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2094_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ),
    .D(net152),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[35][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2095_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ),
    .D(net144),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[35][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2096_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ),
    .D(net136),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[35][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2097_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ),
    .D(net128),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[35][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2098_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ),
    .D(net118),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[35][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2099_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ),
    .D(net109),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[35][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2100_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0718_ ),
    .D(net165),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[61][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2101_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0718_ ),
    .D(net156),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[61][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2102_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0718_ ),
    .D(net150),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[61][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2103_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0718_ ),
    .D(net142),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[61][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2104_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0718_ ),
    .D(net133),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[61][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2105_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0718_ ),
    .D(net125),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[61][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2106_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0718_ ),
    .D(net116),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[61][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2107_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0718_ ),
    .D(net107),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[61][7] ));
 sky130_fd_sc_hd__nand2b_1 \u_usb_host.u_core.u_sie._01_  (.A_N(\u_usb_host.u_core.u_sie.utmi_rxvalid_i ),
    .B(\u_usb_host.u_core.u_sie.utmi_rxactive_i ),
    .Y(\u_usb_host.u_core.u_sie.shift_en_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._02_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net483),
    .RESET_B(net287),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._03_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net471),
    .RESET_B(net288),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._04_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net463),
    .RESET_B(net289),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._05_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net465),
    .RESET_B(net290),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._06_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net464),
    .RESET_B(net290),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._07_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net472),
    .RESET_B(net288),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._08_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net470),
    .RESET_B(net288),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._09_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net475),
    .RESET_B(net287),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._10_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net460),
    .RESET_B(net287),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._11_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net458),
    .RESET_B(net286),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._12_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net452),
    .RESET_B(net289),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._13_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net456),
    .RESET_B(net290),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._14_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net454),
    .RESET_B(net290),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._15_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net455),
    .RESET_B(net288),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._16_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net457),
    .RESET_B(net286),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._17_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net459),
    .RESET_B(net287),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._18_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net478),
    .RESET_B(net287),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._19_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net474),
    .RESET_B(net286),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._20_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net473),
    .RESET_B(net289),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._21_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net466),
    .RESET_B(net289),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._22_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net462),
    .RESET_B(net289),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._23_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net476),
    .RESET_B(net286),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._24_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net480),
    .RESET_B(net286),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._25_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net469),
    .RESET_B(net287),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._26_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net490),
    .RESET_B(net287),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._27_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net444),
    .RESET_B(net286),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._28_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net442),
    .RESET_B(net289),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._29_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net445),
    .RESET_B(net289),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._30_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net441),
    .RESET_B(net289),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._31_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net446),
    .RESET_B(net286),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._32_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net440),
    .RESET_B(net286),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._33_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core.u_sie._00_ ),
    .D(net443),
    .RESET_B(net287),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[31] ));
 sky130_fd_sc_hd__dlclkp_4 \u_usb_host.u_core.u_sie._34_  (.CLK(clknet_4_11_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_sie.shift_en_w ),
    .GCLK(\u_usb_host.u_core.u_sie._00_ ));
 sky130_fd_sc_hd__clkbuf_1 \u_usb_host.u_core.u_sie._76_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[0] ),
    .X(\u_usb_host.u_core.fifo_rx_data_w[0] ));
 sky130_fd_sc_hd__clkbuf_1 \u_usb_host.u_core.u_sie._77_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[1] ),
    .X(\u_usb_host.u_core.fifo_rx_data_w[1] ));
 sky130_fd_sc_hd__buf_2 \u_usb_host.u_core.u_sie._78_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[2] ),
    .X(\u_usb_host.u_core.fifo_rx_data_w[2] ));
 sky130_fd_sc_hd__buf_2 \u_usb_host.u_core.u_sie._79_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[3] ),
    .X(\u_usb_host.u_core.fifo_rx_data_w[3] ));
 sky130_fd_sc_hd__clkbuf_2 \u_usb_host.u_core.u_sie._80_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[4] ),
    .X(\u_usb_host.u_core.fifo_rx_data_w[4] ));
 sky130_fd_sc_hd__buf_2 \u_usb_host.u_core.u_sie._81_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[5] ),
    .X(\u_usb_host.u_core.fifo_rx_data_w[5] ));
 sky130_fd_sc_hd__clkbuf_1 \u_usb_host.u_core.u_sie._82_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[6] ),
    .X(\u_usb_host.u_core.fifo_rx_data_w[6] ));
 sky130_fd_sc_hd__clkbuf_2 \u_usb_host.u_core.u_sie._83_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[7] ),
    .X(\u_usb_host.u_core.fifo_rx_data_w[7] ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_phy._194_  (.A(net293),
    .Y(\u_usb_host.u_phy._039_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_phy._195_  (.A(\u_usb_host.u_phy.ones_count_q[0] ),
    .Y(\u_usb_host.u_phy._040_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_phy._196_  (.A(net295),
    .Y(\u_usb_host.u_phy._041_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_phy._197_  (.A(net363),
    .Y(\u_usb_host.u_phy._042_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_phy._197__363  (.LO(net363));
 sky130_fd_sc_hd__and2b_2 \u_usb_host.u_phy._198_  (.A_N(\u_usb_host.u_phy.state_q[2] ),
    .B(net293),
    .X(\u_usb_host.u_phy._043_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._199_  (.A(net294),
    .B(net295),
    .Y(\u_usb_host.u_phy._044_ ));
 sky130_fd_sc_hd__or2_2 \u_usb_host.u_phy._200_  (.A(\u_usb_host.u_phy.state_q[1] ),
    .B(net295),
    .X(\u_usb_host.u_phy._045_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_phy._201_  (.A(\u_usb_host.u_phy.state_q[2] ),
    .B(\u_usb_host.u_phy._039_ ),
    .C(net294),
    .X(\u_usb_host.u_phy._046_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._202_  (.A(net295),
    .B(\u_usb_host.u_phy._046_ ),
    .X(\u_usb_host.u_phy._047_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_phy._203_  (.A(\u_usb_host.u_phy._047_ ),
    .Y(\u_usb_host.u_phy._159_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._204_  (.A(\u_usb_host.u_phy.sample_cnt_q[1] ),
    .B(\u_usb_host.u_phy.sample_cnt_q[0] ),
    .X(\u_usb_host.u_phy._048_ ));
 sky130_fd_sc_hd__nor3_4 \u_usb_host.u_phy._205_  (.A(\u_usb_host.u_phy.sample_cnt_q[2] ),
    .B(\u_usb_host.u_phy.sample_cnt_q[1] ),
    .C(\u_usb_host.u_phy.sample_cnt_q[0] ),
    .Y(\u_usb_host.u_phy._049_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_phy._206_  (.A(\u_usb_host.u_phy.sample_cnt_q[2] ),
    .B(\u_usb_host.u_phy.sample_cnt_q[1] ),
    .C(\u_usb_host.u_phy.sample_cnt_q[0] ),
    .X(\u_usb_host.u_phy._050_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_phy._207_  (.A_N(\u_usb_host.u_phy.ones_count_q[0] ),
    .B(\u_usb_host.u_phy.ones_count_q[1] ),
    .X(\u_usb_host.u_phy._051_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_phy._208_  (.A(\u_usb_host.u_phy.ones_count_q[2] ),
    .B(\u_usb_host.u_phy._051_ ),
    .X(\u_usb_host.u_phy._052_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_phy._209_  (.A(\u_usb_host.u_phy.ones_count_q[2] ),
    .B(\u_usb_host.u_phy._051_ ),
    .Y(\u_usb_host.u_phy._053_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_phy._210_  (.A(net294),
    .B(net295),
    .Y(\u_usb_host.u_phy._054_ ));
 sky130_fd_sc_hd__nand2b_1 \u_usb_host.u_phy._211_  (.A_N(net293),
    .B(\u_usb_host.u_phy.state_q[2] ),
    .Y(\u_usb_host.u_phy._055_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_phy._212_  (.A(\u_usb_host.u_phy.state_q[2] ),
    .B(\u_usb_host.u_phy.state_q[1] ),
    .Y(\u_usb_host.u_phy._056_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_phy._213_  (.A(\u_usb_host.u_phy._054_ ),
    .B(\u_usb_host.u_phy._055_ ),
    .Y(\u_usb_host.u_phy._057_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_phy._214_  (.A(\u_usb_host.u_phy.state_q[2] ),
    .B(net293),
    .X(\u_usb_host.u_phy._058_ ));
 sky130_fd_sc_hd__nand2_2 \u_usb_host.u_phy._215_  (.A(\u_usb_host.u_phy.state_q[2] ),
    .B(net293),
    .Y(\u_usb_host.u_phy._059_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._216_  (.A(\u_usb_host.u_phy.state_q[2] ),
    .B(net293),
    .Y(\u_usb_host.u_phy._060_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._217_  (.A(\u_usb_host.u_phy.state_q[2] ),
    .B(net293),
    .X(\u_usb_host.u_phy._061_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._218_  (.A(\u_usb_host.u_phy._043_ ),
    .B(\u_usb_host.u_phy._057_ ),
    .Y(\u_usb_host.u_phy._062_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._219_  (.A(net293),
    .B(net295),
    .Y(\u_usb_host.u_phy._063_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._220_  (.A(\u_usb_host.u_phy.state_q[0] ),
    .B(\u_usb_host.u_phy._061_ ),
    .Y(\u_usb_host.u_phy._030_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._221_  (.A(\u_usb_host.u_phy._045_ ),
    .B(\u_usb_host.u_phy._061_ ),
    .Y(\u_usb_host.u_phy._064_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_phy._222_  (.A(\u_usb_host.u_phy.state_q[2] ),
    .B(net293),
    .C(net294),
    .D(net295),
    .X(\u_usb_host.u_phy._065_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._223_  (.A(net294),
    .B(\u_usb_host.u_phy._059_ ),
    .Y(\u_usb_host.u_phy._066_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_phy._224_  (.A(net294),
    .B(\u_usb_host.u_phy._043_ ),
    .Y(\u_usb_host.u_phy._067_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_phy._225_  (.A(\u_usb_host.u_phy._043_ ),
    .B(\u_usb_host.u_phy._057_ ),
    .C(\u_usb_host.u_phy._064_ ),
    .D(\u_usb_host.u_phy._066_ ),
    .X(\u_usb_host.u_phy._068_ ));
 sky130_fd_sc_hd__or3_2 \u_usb_host.u_phy._226_  (.A(\u_usb_host.u_phy._045_ ),
    .B(\u_usb_host.u_phy._049_ ),
    .C(\u_usb_host.u_phy._059_ ),
    .X(\u_usb_host.u_phy._069_ ));
 sky130_fd_sc_hd__or4b_1 \u_usb_host.u_phy._227_  (.A(\u_usb_host.u_phy._046_ ),
    .B(\u_usb_host.u_phy._052_ ),
    .C(net102),
    .D_N(\u_usb_host.u_core.u_sie.utmi_data_i[0] ),
    .X(\u_usb_host.u_phy._070_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_phy._228_  (.A1(net294),
    .A2(\u_usb_host.u_phy._043_ ),
    .B1(net102),
    .Y(\u_usb_host.u_phy._071_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_phy._229_  (.A(\u_usb_host.u_phy._068_ ),
    .B(\u_usb_host.u_phy._069_ ),
    .C(\u_usb_host.u_phy._070_ ),
    .D(\u_usb_host.u_phy._071_ ),
    .X(\u_usb_host.u_phy._037_ ));
 sky130_fd_sc_hd__o211a_1 \u_usb_host.u_phy._230_  (.A1(\u_usb_host.u_phy._058_ ),
    .A2(\u_usb_host.u_phy._060_ ),
    .B1(\u_usb_host.u_phy._069_ ),
    .C1(\u_usb_host.u_phy._044_ ),
    .X(\u_usb_host.u_phy._024_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_phy._231_  (.A(\u_usb_host.u_phy._045_ ),
    .B(\u_usb_host.u_phy._055_ ),
    .Y(\u_usb_host.u_core.u_sie.utmi_rxactive_i ));
 sky130_fd_sc_hd__nor2_4 \u_usb_host.u_phy._232_  (.A(\u_usb_host.u_phy._039_ ),
    .B(\u_usb_host.u_phy._056_ ),
    .Y(\u_usb_host.u_phy._072_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_phy._233_  (.A(\u_usb_host.u_phy._072_ ),
    .Y(\u_usb_host.u_phy._031_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_phy._234_  (.A(\u_usb_host.u_phy._065_ ),
    .B(\u_usb_host.u_phy._031_ ),
    .X(\u_usb_host.u_phy._073_ ));
 sky130_fd_sc_hd__o211a_1 \u_usb_host.u_phy._235_  (.A1(\u_usb_host.u_phy._049_ ),
    .A2(\u_usb_host.u_phy._060_ ),
    .B1(\u_usb_host.u_phy._059_ ),
    .C1(\u_usb_host.u_phy._044_ ),
    .X(\u_usb_host.u_phy._026_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_phy._236_  (.A(\u_usb_host.u_phy._044_ ),
    .B(\u_usb_host.u_phy._059_ ),
    .C(\u_usb_host.u_phy._061_ ),
    .X(\u_usb_host.u_phy._074_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_phy._237_  (.A(\u_usb_host.u_phy._057_ ),
    .B(\u_usb_host.u_phy._074_ ),
    .Y(\u_usb_host.u_phy._075_ ));
 sky130_fd_sc_hd__a2bb2o_1 \u_usb_host.u_phy._238_  (.A1_N(\u_usb_host.u_phy._049_ ),
    .A2_N(\u_usb_host.u_phy._075_ ),
    .B1(\u_usb_host.u_phy._074_ ),
    .B2(\u_usb_host.u_phy._052_ ),
    .X(\u_usb_host.u_phy._076_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_phy._239_  (.A1(\u_usb_host.u_phy._065_ ),
    .A2(\u_usb_host.u_phy._075_ ),
    .B1(\u_usb_host.u_phy._076_ ),
    .Y(\u_usb_host.u_phy._028_ ));
 sky130_fd_sc_hd__o211a_1 \u_usb_host.u_phy._240_  (.A1(net294),
    .A2(\u_usb_host.u_phy._042_ ),
    .B1(\u_usb_host.u_phy._043_ ),
    .C1(\u_usb_host.u_phy._041_ ),
    .X(\u_usb_host.u_phy._029_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_phy._241_  (.A(net294),
    .B(\u_usb_host.u_phy._030_ ),
    .Y(\u_usb_host.u_phy._077_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_phy._242_  (.A(\u_usb_host.u_phy._077_ ),
    .Y(\u_usb_host.u_phy._160_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._243_  (.A(\u_usb_host.u_phy.rx_dn_q ),
    .B(\u_usb_host.u_phy.rx_dp_q ),
    .Y(\u_usb_host.u_phy._078_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._244_  (.A(\u_usb_host.u_phy.rx_dn_q ),
    .B(\u_usb_host.u_phy.rx_dp_q ),
    .X(\u_usb_host.u_phy._079_ ));
 sky130_fd_sc_hd__o21a_2 \u_usb_host.u_phy._245_  (.A1(\u_usb_host.u_phy.rx_dn_q ),
    .A2(\u_usb_host.u_phy.rx_dp_q ),
    .B1(\u_usb_host.u_phy.rxd_q ),
    .X(\u_usb_host.u_phy.in_j_w ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_phy._246_  (.A(\u_usb_host.u_phy.bit_count_q[1] ),
    .B(\u_usb_host.u_phy.bit_count_q[0] ),
    .Y(\u_usb_host.u_phy._080_ ));
 sky130_fd_sc_hd__nand3_2 \u_usb_host.u_phy._247_  (.A(\u_usb_host.u_phy.bit_count_q[2] ),
    .B(\u_usb_host.u_phy.bit_count_q[1] ),
    .C(\u_usb_host.u_phy.bit_count_q[0] ),
    .Y(\u_usb_host.u_phy._081_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._248_  (.A(net102),
    .B(\u_usb_host.u_phy._081_ ),
    .Y(\u_usb_host.u_phy._082_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._249_  (.A(net102),
    .B(\u_usb_host.u_phy._081_ ),
    .X(\u_usb_host.u_phy._083_ ));
 sky130_fd_sc_hd__o211a_1 \u_usb_host.u_phy._250_  (.A1(\u_usb_host.u_phy._042_ ),
    .A2(\u_usb_host.u_phy.send_eop_q ),
    .B1(\u_usb_host.u_phy._053_ ),
    .C1(\u_usb_host.u_phy._082_ ),
    .X(\u_usb_host.u_phy._084_ ));
 sky130_fd_sc_hd__nor4_1 \u_usb_host.u_phy._251_  (.A(\u_usb_host.u_core.utmi_xcvrselect_o[1] ),
    .B(\u_usb_host.u_core.utmi_xcvrselect_o[0] ),
    .C(\u_usb_host.u_core.utmi_termselect_o ),
    .D(\u_usb_host.u_core.utmi_op_mode_o[0] ),
    .Y(\u_usb_host.u_phy._085_ ));
 sky130_fd_sc_hd__a41o_1 \u_usb_host.u_phy._252_  (.A1(\u_usb_host.u_core.utmi_op_mode_o[1] ),
    .A2(\u_usb_host.u_core.utmi_dppulldown_o ),
    .A3(\u_usb_host.u_core.utmi_dmpulldown_o ),
    .A4(\u_usb_host.u_phy._085_ ),
    .B1(net322),
    .X(\u_usb_host.u_phy._086_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_phy._252__322  (.LO(net322));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._253_  (.A(net364),
    .B(\u_usb_host.u_phy._086_ ),
    .X(\u_usb_host.u_phy._087_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_phy._253__364  (.LO(net364));
 sky130_fd_sc_hd__o21ba_1 \u_usb_host.u_phy._254_  (.A1(\u_usb_host.u_phy.rx_dn_q ),
    .A2(\u_usb_host.u_phy.rx_dp_q ),
    .B1_N(\u_usb_host.u_phy.rxd_q ),
    .X(\u_usb_host.u_phy._088_ ));
 sky130_fd_sc_hd__o32a_1 \u_usb_host.u_phy._255_  (.A1(\u_usb_host.u_phy._065_ ),
    .A2(\u_usb_host.u_phy._087_ ),
    .A3(\u_usb_host.u_phy._088_ ),
    .B1(\u_usb_host.u_phy._084_ ),
    .B2(\u_usb_host.u_phy._047_ ),
    .X(\u_usb_host.u_phy._089_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_phy._256_  (.A(\u_usb_host.u_phy._049_ ),
    .B(\u_usb_host.u_phy._088_ ),
    .X(\u_usb_host.u_phy._090_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_phy._257_  (.A(\u_usb_host.u_phy._049_ ),
    .B(\u_usb_host.u_phy._088_ ),
    .Y(\u_usb_host.u_phy._091_ ));
 sky130_fd_sc_hd__or4b_1 \u_usb_host.u_phy._258_  (.A(\u_usb_host.u_phy.bit_count_q[2] ),
    .B(net103),
    .C(\u_usb_host.u_phy.bit_count_q[1] ),
    .D_N(\u_usb_host.u_phy.bit_count_q[0] ),
    .X(\u_usb_host.u_phy._092_ ));
 sky130_fd_sc_hd__or3b_1 \u_usb_host.u_phy._259_  (.A(\u_usb_host.u_phy._077_ ),
    .B(\u_usb_host.u_phy._090_ ),
    .C_N(\u_usb_host.u_phy._092_ ),
    .X(\u_usb_host.u_phy._093_ ));
 sky130_fd_sc_hd__and4bb_1 \u_usb_host.u_phy._260_  (.A_N(\u_usb_host.u_phy.state_q[2] ),
    .B_N(\u_usb_host.u_phy.state_q[3] ),
    .C(\u_usb_host.u_phy.state_q[1] ),
    .D(\u_usb_host.u_phy.state_q[0] ),
    .X(\u_usb_host.u_phy._094_ ));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_phy._261_  (.A1(net103),
    .A2(\u_usb_host.u_phy._078_ ),
    .B1(\u_usb_host.u_phy._094_ ),
    .X(\u_usb_host.u_phy._095_ ));
 sky130_fd_sc_hd__nand2b_1 \u_usb_host.u_phy._262_  (.A_N(net294),
    .B(net295),
    .Y(\u_usb_host.u_phy._096_ ));
 sky130_fd_sc_hd__or3b_1 \u_usb_host.u_phy._263_  (.A(\u_usb_host.u_phy._059_ ),
    .B(\u_usb_host.u_phy._096_ ),
    .C_N(\u_usb_host.u_phy._086_ ),
    .X(\u_usb_host.u_phy._097_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_phy._264_  (.A(\u_usb_host.u_phy.rx_dn_q ),
    .B(\u_usb_host.u_phy.rx_dp_q ),
    .Y(\u_usb_host.u_phy._098_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_phy._265_  (.A1(\u_usb_host.u_phy._079_ ),
    .A2(\u_usb_host.u_phy._098_ ),
    .B1(net102),
    .X(\u_usb_host.u_phy._099_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_phy._266_  (.A1(\u_usb_host.u_phy._057_ ),
    .A2(\u_usb_host.u_phy._083_ ),
    .B1(\u_usb_host.u_phy._099_ ),
    .B2(\u_usb_host.u_core.u_sie.utmi_rxactive_i ),
    .X(\u_usb_host.u_phy._100_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_phy._267_  (.A1(\u_usb_host.u_phy._043_ ),
    .A2(\u_usb_host.u_phy._045_ ),
    .A3(net102),
    .B1(\u_usb_host.u_phy._072_ ),
    .C1(\u_usb_host.u_phy._095_ ),
    .X(\u_usb_host.u_phy._101_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._268_  (.A(\u_usb_host.u_phy._100_ ),
    .B(\u_usb_host.u_phy._101_ ),
    .Y(\u_usb_host.u_phy._102_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_phy._269_  (.A(\u_usb_host.u_phy._089_ ),
    .B(\u_usb_host.u_phy._093_ ),
    .C(\u_usb_host.u_phy._097_ ),
    .D(\u_usb_host.u_phy._102_ ),
    .X(\u_usb_host.u_phy._023_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_phy._270_  (.A(\u_usb_host.u_phy.rx_dn1_q ),
    .B(\u_usb_host.u_phy.rx_dn0_q ),
    .X(\u_usb_host.u_phy._004_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._271_  (.A(\u_usb_host.u_phy.rx_dn1_q ),
    .B(\u_usb_host.u_phy.rx_dn0_q ),
    .Y(\u_usb_host.u_phy._103_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._272_  (.A(\u_usb_host.u_phy._004_ ),
    .B(\u_usb_host.u_phy._103_ ),
    .X(\u_usb_host.u_phy._027_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_phy._273_  (.A(\u_usb_host.u_phy.rx_dp1_q ),
    .B(\u_usb_host.u_phy.rx_dp0_q ),
    .X(\u_usb_host.u_phy._005_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._274_  (.A(\u_usb_host.u_phy.rx_dp1_q ),
    .B(\u_usb_host.u_phy.rx_dp0_q ),
    .Y(\u_usb_host.u_phy._104_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._275_  (.A(\u_usb_host.u_phy._005_ ),
    .B(\u_usb_host.u_phy._104_ ),
    .X(\u_usb_host.u_phy._025_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_phy._276_  (.A1(net102),
    .A2(\u_usb_host.u_phy._065_ ),
    .B1(\u_usb_host.u_phy._072_ ),
    .Y(\u_usb_host.u_phy._034_ ));
 sky130_fd_sc_hd__a21boi_1 \u_usb_host.u_phy._281_  (.A1(\u_usb_host.u_phy._060_ ),
    .A2(\u_usb_host.u_phy._096_ ),
    .B1_N(\u_usb_host.u_phy._075_ ),
    .Y(\u_usb_host.u_phy._107_ ));
 sky130_fd_sc_hd__a211oi_1 \u_usb_host.u_phy._282_  (.A1(net103),
    .A2(\u_usb_host.u_phy._160_ ),
    .B1(\u_usb_host.u_phy._107_ ),
    .C1(\u_usb_host.u_phy._076_ ),
    .Y(\u_usb_host.u_phy._036_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._283_  (.A(\u_usb_host.u_phy.adjust_delayed_q ),
    .B(\u_usb_host.u_phy._072_ ),
    .Y(\u_usb_host.u_phy._035_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_phy._284_  (.A(\u_usb_host.u_phy.rxd1_q ),
    .B(\u_usb_host.u_phy.rxd0_q ),
    .X(\u_usb_host.u_phy._009_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._285_  (.A(\u_usb_host.u_phy.rxd1_q ),
    .B(\u_usb_host.u_phy.rxd0_q ),
    .Y(\u_usb_host.u_phy._108_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._286_  (.A(\u_usb_host.u_phy._009_ ),
    .B(\u_usb_host.u_phy._108_ ),
    .X(\u_usb_host.u_phy._021_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_phy._301_  (.A(net438),
    .B(\u_usb_host.u_phy.in_j_w ),
    .X(\u_usb_host.u_phy._116_ ));
 sky130_fd_sc_hd__o211a_1 \u_usb_host.u_phy._302_  (.A1(\u_usb_host.u_phy._041_ ),
    .A2(\u_usb_host.u_phy._056_ ),
    .B1(\u_usb_host.u_phy._116_ ),
    .C1(\u_usb_host.u_phy._039_ ),
    .X(\u_usb_host.u_phy._117_ ));
 sky130_fd_sc_hd__or3b_1 \u_usb_host.u_phy._303_  (.A(\u_usb_host.u_phy.sample_cnt_q[0] ),
    .B(\u_usb_host.u_phy._117_ ),
    .C_N(\u_usb_host.u_phy.sample_cnt_q[1] ),
    .X(\u_usb_host.u_phy._118_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_phy._304_  (.A(net103),
    .B(\u_usb_host.u_phy._118_ ),
    .Y(\u_usb_host.u_phy._010_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_phy._305_  (.A(\u_usb_host.u_phy.sample_cnt_q[1] ),
    .B(\u_usb_host.u_phy.sample_cnt_q[0] ),
    .Y(\u_usb_host.u_phy._119_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_phy._306_  (.A(\u_usb_host.u_phy._048_ ),
    .B(\u_usb_host.u_phy._119_ ),
    .Y(\u_usb_host.u_phy._120_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._307_  (.A(\u_usb_host.u_phy._117_ ),
    .B(\u_usb_host.u_phy._120_ ),
    .Y(\u_usb_host.u_phy._011_ ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_phy._308_  (.A0(\u_usb_host.u_phy._119_ ),
    .A1(\u_usb_host.u_phy._120_ ),
    .S(\u_usb_host.u_phy.sample_cnt_q[2] ),
    .X(\u_usb_host.u_phy._121_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._309_  (.A(\u_usb_host.u_phy._117_ ),
    .B(\u_usb_host.u_phy._121_ ),
    .Y(\u_usb_host.u_phy._012_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._310_  (.A(\u_usb_host.u_phy._064_ ),
    .B(\u_usb_host.u_phy._094_ ),
    .Y(\u_usb_host.u_phy._122_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_phy._311_  (.A_N(\u_usb_host.u_phy.bit_count_q[0] ),
    .B(\u_usb_host.u_phy._122_ ),
    .X(\u_usb_host.u_phy._001_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._312_  (.A(\u_usb_host.u_phy.bit_count_q[1] ),
    .B(\u_usb_host.u_phy.bit_count_q[0] ),
    .X(\u_usb_host.u_phy._123_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_phy._313_  (.A(\u_usb_host.u_phy._080_ ),
    .B(\u_usb_host.u_phy._122_ ),
    .C(\u_usb_host.u_phy._123_ ),
    .X(\u_usb_host.u_phy._002_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_phy._314_  (.A1(\u_usb_host.u_phy.bit_count_q[1] ),
    .A2(\u_usb_host.u_phy.bit_count_q[0] ),
    .B1(\u_usb_host.u_phy.bit_count_q[2] ),
    .X(\u_usb_host.u_phy._124_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_phy._315_  (.A(\u_usb_host.u_phy._081_ ),
    .B(\u_usb_host.u_phy._122_ ),
    .C(\u_usb_host.u_phy._124_ ),
    .X(\u_usb_host.u_phy._003_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_phy._316_  (.A(\u_usb_host.u_phy.ones_count_q[1] ),
    .B(\u_usb_host.u_phy.ones_count_q[2] ),
    .Y(\u_usb_host.u_phy._125_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_phy._317_  (.A1(net295),
    .A2(\u_usb_host.u_phy._060_ ),
    .B1(\u_usb_host.u_phy._058_ ),
    .Y(\u_usb_host.u_phy._126_ ));
 sky130_fd_sc_hd__or4b_1 \u_usb_host.u_phy._318_  (.A(\u_usb_host.u_phy.rxd_q ),
    .B(\u_usb_host.u_phy.sync_j_detected_q ),
    .C(\u_usb_host.u_phy._078_ ),
    .D_N(\u_usb_host.u_phy.state_q[1] ),
    .X(\u_usb_host.u_phy._127_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_phy._319_  (.A1(\u_usb_host.u_phy._126_ ),
    .A2(\u_usb_host.u_phy._127_ ),
    .B1(\u_usb_host.u_phy._098_ ),
    .Y(\u_usb_host.u_phy._128_ ));
 sky130_fd_sc_hd__a2bb2o_1 \u_usb_host.u_phy._320_  (.A1_N(\u_usb_host.u_phy._040_ ),
    .A2_N(\u_usb_host.u_phy._125_ ),
    .B1(\u_usb_host.u_phy._128_ ),
    .B2(\u_usb_host.u_phy._049_ ),
    .X(\u_usb_host.u_phy._007_ ));
 sky130_fd_sc_hd__mux2_2 \u_usb_host.u_phy._321_  (.A0(\u_usb_host.u_phy.usb_tx_dp_o ),
    .A1(\u_usb_host.u_phy.rx_dp_q ),
    .S(\u_usb_host.u_phy.usb_tx_oen_o ),
    .X(\u_usb_host.u_core.u_sie.utmi_linestate_i[0] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_phy._322_  (.A0(\u_usb_host.u_phy.usb_tx_dn_o ),
    .A1(\u_usb_host.u_phy.rx_dn_q ),
    .S(\u_usb_host.u_phy.usb_tx_oen_o ),
    .X(\u_usb_host.u_core.u_sie.utmi_linestate_i[1] ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_phy._323_  (.A1(net461),
    .A2(\u_usb_host.u_phy.in_j_w ),
    .B1(net102),
    .Y(\u_usb_host.u_phy._129_ ));
 sky130_fd_sc_hd__o21ai_2 \u_usb_host.u_phy._324_  (.A1(net461),
    .A2(\u_usb_host.u_phy.in_j_w ),
    .B1(\u_usb_host.u_phy._129_ ),
    .Y(\u_usb_host.u_phy._130_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._325_  (.A(\u_usb_host.u_phy._040_ ),
    .B(\u_usb_host.u_phy.ones_count_q[1] ),
    .Y(\u_usb_host.u_phy._131_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_phy._326_  (.A(\u_usb_host.u_phy.ones_count_q[2] ),
    .B(\u_usb_host.u_phy._159_ ),
    .C(\u_usb_host.u_phy._130_ ),
    .D(\u_usb_host.u_phy._131_ ),
    .X(\u_usb_host.u_phy._132_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_phy._327_  (.A(\u_usb_host.u_phy._045_ ),
    .B(\u_usb_host.u_phy._054_ ),
    .C(\u_usb_host.u_phy._060_ ),
    .D(\u_usb_host.u_phy._090_ ),
    .X(\u_usb_host.u_phy._133_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_phy._328_  (.A(\u_usb_host.u_phy._045_ ),
    .B(net102),
    .C(\u_usb_host.u_phy._055_ ),
    .D(\u_usb_host.u_phy._079_ ),
    .X(\u_usb_host.u_phy._134_ ));
 sky130_fd_sc_hd__o311a_1 \u_usb_host.u_phy._329_  (.A1(net293),
    .A2(\u_usb_host.u_phy._049_ ),
    .A3(\u_usb_host.u_phy._096_ ),
    .B1(\u_usb_host.u_phy._134_ ),
    .C1(\u_usb_host.u_phy._073_ ),
    .X(\u_usb_host.u_phy._135_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_phy._330_  (.A1(net295),
    .A2(\u_usb_host.u_phy._067_ ),
    .B1(\u_usb_host.u_phy._135_ ),
    .Y(\u_usb_host.u_phy._136_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_phy._331_  (.A(\u_usb_host.u_phy._132_ ),
    .B(\u_usb_host.u_phy._133_ ),
    .C(\u_usb_host.u_phy._136_ ),
    .X(\u_usb_host.u_phy.next_state_r[0] ));
 sky130_fd_sc_hd__a31oi_1 \u_usb_host.u_phy._332_  (.A1(\u_usb_host.u_phy.ones_count_q[2] ),
    .A2(\u_usb_host.u_phy._130_ ),
    .A3(\u_usb_host.u_phy._131_ ),
    .B1(\u_usb_host.u_phy._047_ ),
    .Y(\u_usb_host.u_phy._137_ ));
 sky130_fd_sc_hd__and3b_1 \u_usb_host.u_phy._333_  (.A_N(\u_usb_host.u_phy._056_ ),
    .B(\u_usb_host.u_phy._063_ ),
    .C(net102),
    .X(\u_usb_host.u_phy._138_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_phy._334_  (.A(\u_usb_host.u_phy._043_ ),
    .B(\u_usb_host.u_phy._045_ ),
    .C(\u_usb_host.u_phy._054_ ),
    .X(\u_usb_host.u_phy._139_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._335_  (.A(\u_usb_host.u_phy._055_ ),
    .B(\u_usb_host.u_phy._096_ ),
    .Y(\u_usb_host.u_phy._140_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_phy._336_  (.A(\u_usb_host.u_phy._049_ ),
    .B(\u_usb_host.u_phy._078_ ),
    .C(\u_usb_host.u_phy._140_ ),
    .X(\u_usb_host.u_phy._141_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_phy._337_  (.A1(\u_usb_host.u_phy._091_ ),
    .A2(\u_usb_host.u_phy._094_ ),
    .B1(\u_usb_host.u_phy._138_ ),
    .Y(\u_usb_host.u_phy._142_ ));
 sky130_fd_sc_hd__or4b_1 \u_usb_host.u_phy._338_  (.A(\u_usb_host.u_phy._133_ ),
    .B(\u_usb_host.u_phy._139_ ),
    .C(\u_usb_host.u_phy._141_ ),
    .D_N(\u_usb_host.u_phy._142_ ),
    .X(\u_usb_host.u_phy._143_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._339_  (.A(\u_usb_host.u_phy._073_ ),
    .B(\u_usb_host.u_phy._088_ ),
    .X(\u_usb_host.u_phy._144_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_phy._340_  (.A(\u_usb_host.u_phy._144_ ),
    .Y(\u_usb_host.u_phy._145_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_phy._341_  (.A1(net365),
    .A2(\u_usb_host.u_phy._145_ ),
    .B1(\u_usb_host.u_phy._143_ ),
    .C1(\u_usb_host.u_phy._137_ ),
    .X(\u_usb_host.u_phy.next_state_r[1] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_phy._341__365  (.LO(net365));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_phy._342_  (.A1(net103),
    .A2(\u_usb_host.u_phy._078_ ),
    .B1(\u_usb_host.u_phy._140_ ),
    .X(\u_usb_host.u_phy._146_ ));
 sky130_fd_sc_hd__o211ai_1 \u_usb_host.u_phy._343_  (.A1(\u_usb_host.u_phy._041_ ),
    .A2(\u_usb_host.u_phy._067_ ),
    .B1(\u_usb_host.u_phy._069_ ),
    .C1(\u_usb_host.u_phy._134_ ),
    .Y(\u_usb_host.u_phy._147_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_phy._344_  (.A1(net436),
    .A2(\u_usb_host.u_phy._090_ ),
    .A3(\u_usb_host.u_phy._094_ ),
    .B1(\u_usb_host.u_phy._147_ ),
    .X(\u_usb_host.u_phy._148_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_phy._345_  (.A(\u_usb_host.u_phy._138_ ),
    .B(\u_usb_host.u_phy._145_ ),
    .C(\u_usb_host.u_phy._146_ ),
    .D(\u_usb_host.u_phy._148_ ),
    .X(\u_usb_host.u_phy.next_state_r[2] ));
 sky130_fd_sc_hd__o211ai_1 \u_usb_host.u_phy._346_  (.A1(net366),
    .A2(\u_usb_host.u_phy._144_ ),
    .B1(\u_usb_host.u_phy._069_ ),
    .C1(\u_usb_host.u_phy._062_ ),
    .Y(\u_usb_host.u_phy.next_state_r[3] ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_phy._346__366  (.LO(net366));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_phy._349_  (.A1(\u_usb_host.u_core.u_sie.utmi_data_i[0] ),
    .A2(\u_usb_host.u_phy._159_ ),
    .A3(\u_usb_host.u_phy._053_ ),
    .B1(\u_usb_host.u_core.u_sie.utmi_rxactive_i ),
    .B2(\u_usb_host.u_phy._130_ ),
    .X(\u_usb_host.u_phy._150_ ));
 sky130_fd_sc_hd__a21bo_1 \u_usb_host.u_phy._350_  (.A1(\u_usb_host.u_phy._040_ ),
    .A2(\u_usb_host.u_phy._150_ ),
    .B1_N(\u_usb_host.u_phy._074_ ),
    .X(\u_usb_host.u_phy._169_ ));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_phy._351_  (.A1(\u_usb_host.u_phy._051_ ),
    .A2(\u_usb_host.u_phy._131_ ),
    .B1(\u_usb_host.u_phy._150_ ),
    .X(\u_usb_host.u_phy._170_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_phy._352_  (.A1(\u_usb_host.u_phy.ones_count_q[0] ),
    .A2(\u_usb_host.u_phy.ones_count_q[1] ),
    .B1(\u_usb_host.u_phy.ones_count_q[2] ),
    .X(\u_usb_host.u_phy._151_ ));
 sky130_fd_sc_hd__o211a_1 \u_usb_host.u_phy._353_  (.A1(\u_usb_host.u_phy._040_ ),
    .A2(\u_usb_host.u_phy._125_ ),
    .B1(\u_usb_host.u_phy._150_ ),
    .C1(\u_usb_host.u_phy._151_ ),
    .X(\u_usb_host.u_phy._171_ ));
 sky130_fd_sc_hd__o21ba_2 \u_usb_host.u_phy._354_  (.A1(\u_usb_host.u_phy._159_ ),
    .A2(\u_usb_host.u_phy._057_ ),
    .B1_N(\u_usb_host.u_phy._081_ ),
    .X(\u_usb_host.u_phy._152_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._355_  (.A(\u_usb_host.u_core.u_sie.utmi_rxactive_i ),
    .B(\u_usb_host.u_phy._081_ ),
    .X(\u_usb_host.u_phy._153_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_phy._356_  (.A_N(\u_usb_host.u_phy._075_ ),
    .B(\u_usb_host.u_phy._153_ ),
    .X(\u_usb_host.u_phy._154_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_phy._357_  (.A1(net355),
    .A2(\u_usb_host.u_phy._152_ ),
    .B1(\u_usb_host.u_phy._154_ ),
    .B2(\u_usb_host.u_core.u_sie.utmi_data_i[1] ),
    .X(\u_usb_host.u_phy._161_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_phy._357__355  (.LO(net355));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_phy._358_  (.A1(net356),
    .A2(\u_usb_host.u_phy._152_ ),
    .B1(\u_usb_host.u_phy._153_ ),
    .B2(\u_usb_host.u_core.u_sie.utmi_data_i[2] ),
    .C1(\u_usb_host.u_phy._075_ ),
    .X(\u_usb_host.u_phy._162_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_phy._358__356  (.LO(net356));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_phy._359_  (.A1(net357),
    .A2(\u_usb_host.u_phy._152_ ),
    .B1(\u_usb_host.u_phy._154_ ),
    .B2(\u_usb_host.u_core.u_sie.utmi_data_i[3] ),
    .X(\u_usb_host.u_phy._163_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_phy._359__357  (.LO(net357));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_phy._360_  (.A1(net358),
    .A2(\u_usb_host.u_phy._152_ ),
    .B1(\u_usb_host.u_phy._153_ ),
    .B2(\u_usb_host.u_core.u_sie.utmi_data_i[4] ),
    .C1(\u_usb_host.u_phy._075_ ),
    .X(\u_usb_host.u_phy._164_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_phy._360__358  (.LO(net358));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_phy._361_  (.A1(net359),
    .A2(\u_usb_host.u_phy._152_ ),
    .B1(\u_usb_host.u_phy._154_ ),
    .B2(\u_usb_host.u_core.u_sie.utmi_data_i[5] ),
    .X(\u_usb_host.u_phy._165_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_phy._361__359  (.LO(net359));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_phy._362_  (.A1(net360),
    .A2(\u_usb_host.u_phy._152_ ),
    .B1(\u_usb_host.u_phy._153_ ),
    .B2(\u_usb_host.u_core.u_sie.utmi_data_i[6] ),
    .C1(\u_usb_host.u_phy._075_ ),
    .X(\u_usb_host.u_phy._166_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_phy._362__360  (.LO(net360));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_phy._363_  (.A1(net361),
    .A2(\u_usb_host.u_phy._152_ ),
    .B1(\u_usb_host.u_phy._154_ ),
    .B2(\u_usb_host.u_core.u_sie.utmi_data_i[7] ),
    .X(\u_usb_host.u_phy._167_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_phy._363__361  (.LO(net361));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_phy._364_  (.A1(net362),
    .A2(\u_usb_host.u_phy._152_ ),
    .B1(\u_usb_host.u_phy._154_ ),
    .B2(\u_usb_host.u_phy._130_ ),
    .X(\u_usb_host.u_phy._168_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_phy._364__362  (.LO(net362));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_phy._365_  (.A1(\u_usb_host.u_phy._059_ ),
    .A2(\u_usb_host.u_phy._096_ ),
    .B1(\u_usb_host.u_phy._062_ ),
    .X(\u_usb_host.u_phy._155_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._366_  (.A(\u_usb_host.u_phy.usb_tx_dp_o ),
    .B(\u_usb_host.u_phy._046_ ),
    .Y(\u_usb_host.u_phy._156_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_phy._367_  (.A1(\u_usb_host.u_core.u_sie.utmi_data_i[0] ),
    .A2(\u_usb_host.u_phy._057_ ),
    .B1(\u_usb_host.u_phy._155_ ),
    .C1(\u_usb_host.u_phy._156_ ),
    .X(\u_usb_host.u_phy._193_ ));
 sky130_fd_sc_hd__or4b_1 \u_usb_host.u_phy._368_  (.A(\u_usb_host.u_phy.usb_tx_dn_o ),
    .B(\u_usb_host.u_phy._064_ ),
    .C(\u_usb_host.u_phy._066_ ),
    .D_N(\u_usb_host.u_phy._067_ ),
    .X(\u_usb_host.u_phy._157_ ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_phy._369_  (.A0(\u_usb_host.u_phy._157_ ),
    .A1(\u_usb_host.u_core.u_sie.utmi_data_i[0] ),
    .S(\u_usb_host.u_phy._057_ ),
    .X(\u_usb_host.u_phy._158_ ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_phy._370_  (.A(\u_usb_host.u_phy._158_ ),
    .Y(\u_usb_host.u_phy._192_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_phy._371_  (.A(\u_usb_host.u_phy._053_ ),
    .B(\u_usb_host.u_core.u_sie.utmi_rxactive_i ),
    .C(\u_usb_host.u_phy._082_ ),
    .X(\u_usb_host.u_phy._008_ ));
 sky130_fd_sc_hd__and3b_1 \u_usb_host.u_phy._372_  (.A_N(\u_usb_host.u_phy.adjust_delayed_q ),
    .B(\u_usb_host.u_phy._049_ ),
    .C(\u_usb_host.u_phy._117_ ),
    .X(\u_usb_host.u_phy._000_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_phy._373_  (.A1(\u_usb_host.u_phy._045_ ),
    .A2(\u_usb_host.u_phy._059_ ),
    .B1(\u_usb_host.u_phy._087_ ),
    .Y(\u_usb_host.u_phy._006_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_phy._374_  (.A(\u_usb_host.u_phy._068_ ),
    .B(\u_usb_host.u_phy._069_ ),
    .C(\u_usb_host.u_phy._070_ ),
    .D(\u_usb_host.u_phy._071_ ),
    .X(\u_usb_host.u_phy._038_ ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_phy._375_  (.A(\u_usb_host.u_phy._072_ ),
    .Y(\u_usb_host.u_phy._033_ ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_phy._376_  (.A(\u_usb_host.u_phy._072_ ),
    .Y(\u_usb_host.u_phy._032_ ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._378_  (.CLK(\u_usb_host.u_phy._179_ ),
    .D(\u_usb_host.u_phy._004_ ),
    .RESET_B(net283),
    .Q(\u_usb_host.u_phy.rx_dn_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._379_  (.CLK(\u_usb_host.u_phy._181_ ),
    .D(\u_usb_host.u_phy._159_ ),
    .RESET_B(net282),
    .Q(\u_usb_host.u_phy.send_eop_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._380_  (.CLK(\u_usb_host.u_phy._182_ ),
    .D(\u_usb_host.u_phy._160_ ),
    .RESET_B(net285),
    .Q(\u_usb_host.u_phy.sync_j_detected_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._381_  (.CLK(\u_usb_host.u_phy._183_ ),
    .D(\u_usb_host.u_phy._007_ ),
    .RESET_B(net280),
    .Q(\u_usb_host.u_core.utmi_rxerror_i ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._382_  (.CLK(\u_usb_host.u_phy._189_ ),
    .D(\u_usb_host.u_phy._192_ ),
    .RESET_B(net283),
    .Q(\u_usb_host.u_phy.usb_tx_dn_o ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._383_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_phy._188_ ),
    .D(\u_usb_host.u_phy._001_ ),
    .RESET_B(net284),
    .Q(\u_usb_host.u_phy.bit_count_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._384_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._188_ ),
    .D(\u_usb_host.u_phy._002_ ),
    .RESET_B(net284),
    .Q(\u_usb_host.u_phy.bit_count_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._385_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._188_ ),
    .D(\u_usb_host.u_phy._003_ ),
    .RESET_B(net285),
    .Q(\u_usb_host.u_phy.bit_count_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._386_  (.CLK(\u_usb_host.u_phy._184_ ),
    .D(\u_usb_host.u_phy._000_ ),
    .RESET_B(net284),
    .Q(\u_usb_host.u_phy.adjust_delayed_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._387_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_phy._187_ ),
    .D(\u_usb_host.u_phy._010_ ),
    .RESET_B(net290),
    .Q(\u_usb_host.u_phy.sample_cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._388_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._187_ ),
    .D(\u_usb_host.u_phy._011_ ),
    .RESET_B(net290),
    .Q(\u_usb_host.u_phy.sample_cnt_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._389_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._187_ ),
    .D(\u_usb_host.u_phy._012_ ),
    .RESET_B(net290),
    .Q(\u_usb_host.u_phy.sample_cnt_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._390_  (.CLK(\u_usb_host.u_phy._185_ ),
    .D(\u_usb_host.u_phy._008_ ),
    .RESET_B(net280),
    .Q(\u_usb_host.u_core.u_sie.utmi_rxvalid_i ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._391_  (.CLK(\u_usb_host.u_phy._173_ ),
    .D(\u_usb_host.u_phy._009_ ),
    .RESET_B(net283),
    .Q(\u_usb_host.u_phy.rxd_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._392_  (.CLK(\u_usb_host.u_phy._177_ ),
    .D(\u_usb_host.u_phy._005_ ),
    .RESET_B(net283),
    .Q(\u_usb_host.u_phy.rx_dp_q ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_phy._393_  (.CLK(\u_usb_host.u_phy._190_ ),
    .D(\u_usb_host.u_phy._193_ ),
    .RESET_B(net281),
    .Q(\u_usb_host.u_phy.usb_tx_dp_o ));
 sky130_fd_sc_hd__dfstp_1 \u_usb_host.u_phy._394_  (.CLK(\u_usb_host.u_phy._176_ ),
    .D(\u_usb_host.u_phy._006_ ),
    .SET_B(net283),
    .Q(\u_usb_host.u_phy.usb_tx_oen_o ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._395_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_phy._175_ ),
    .D(\u_usb_host.u_phy.next_state_r[0] ),
    .RESET_B(net285),
    .Q(\u_usb_host.u_phy.state_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._396_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._175_ ),
    .D(\u_usb_host.u_phy.next_state_r[1] ),
    .RESET_B(net282),
    .Q(\u_usb_host.u_phy.state_q[1] ));
 sky130_fd_sc_hd__dfrtp_4 \u_usb_host.u_phy._397_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_phy._175_ ),
    .D(\u_usb_host.u_phy.next_state_r[2] ),
    .RESET_B(net284),
    .Q(\u_usb_host.u_phy.state_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._398_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._175_ ),
    .D(\u_usb_host.u_phy.next_state_r[3] ),
    .RESET_B(net282),
    .Q(\u_usb_host.u_phy.state_q[3] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_phy._406_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._180_ ),
    .D(\u_usb_host.u_phy._161_ ),
    .RESET_B(net286),
    .Q(\u_usb_host.u_core.u_sie.utmi_data_i[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._407_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._180_ ),
    .D(\u_usb_host.u_phy._162_ ),
    .RESET_B(net280),
    .Q(\u_usb_host.u_core.u_sie.utmi_data_i[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._408_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_phy._180_ ),
    .D(\u_usb_host.u_phy._163_ ),
    .RESET_B(net289),
    .Q(\u_usb_host.u_core.u_sie.utmi_data_i[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._409_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_phy._180_ ),
    .D(\u_usb_host.u_phy._164_ ),
    .RESET_B(net284),
    .Q(\u_usb_host.u_core.u_sie.utmi_data_i[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._410_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_phy._180_ ),
    .D(\u_usb_host.u_phy._165_ ),
    .RESET_B(net289),
    .Q(\u_usb_host.u_core.u_sie.utmi_data_i[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._411_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_phy._180_ ),
    .D(\u_usb_host.u_phy._166_ ),
    .RESET_B(net280),
    .Q(\u_usb_host.u_core.u_sie.utmi_data_i[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._412_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._180_ ),
    .D(\u_usb_host.u_phy._167_ ),
    .RESET_B(net286),
    .Q(\u_usb_host.u_core.u_sie.utmi_data_i[6] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._413_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._180_ ),
    .D(\u_usb_host.u_phy._168_ ),
    .RESET_B(net282),
    .Q(\u_usb_host.u_core.u_sie.utmi_data_i[7] ));
 sky130_fd_sc_hd__dfstp_1 \u_usb_host.u_phy._414_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._178_ ),
    .D(\u_usb_host.u_phy._169_ ),
    .SET_B(net280),
    .Q(\u_usb_host.u_phy.ones_count_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._415_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._178_ ),
    .D(\u_usb_host.u_phy._170_ ),
    .RESET_B(net280),
    .Q(\u_usb_host.u_phy.ones_count_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._416_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_phy._178_ ),
    .D(\u_usb_host.u_phy._171_ ),
    .RESET_B(net280),
    .Q(\u_usb_host.u_phy.ones_count_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._418_  (.CLK(\u_usb_host.u_phy._186_ ),
    .D(\u_usb_host.u_phy.in_j_w ),
    .RESET_B(net281),
    .Q(\u_usb_host.u_phy.rxd_last_j_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._419_  (.CLK(clknet_4_10_0_usb_clk),
    .D(\u_usb_host.u_phy.usb_rx_dp_i ),
    .RESET_B(net284),
    .Q(\u_usb_host.u_phy.rx_dp_ms ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._420_  (.CLK(clknet_4_10_0_usb_clk),
    .D(\u_usb_host.u_phy.usb_rx_dn_i ),
    .RESET_B(net284),
    .Q(\u_usb_host.u_phy.rx_dn_ms ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._421_  (.CLK(clknet_4_10_0_usb_clk),
    .D(\u_usb_host.u_phy.usb_rx_rcv_i ),
    .RESET_B(net284),
    .Q(\u_usb_host.u_phy.rxd_ms ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._422_  (.CLK(clknet_4_10_0_usb_clk),
    .D(net492),
    .RESET_B(net283),
    .Q(\u_usb_host.u_phy.rx_dp0_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._423_  (.CLK(clknet_4_10_0_usb_clk),
    .D(\u_usb_host.u_phy.rx_dn_ms ),
    .RESET_B(net283),
    .Q(\u_usb_host.u_phy.rx_dn0_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._424_  (.CLK(clknet_4_10_0_usb_clk),
    .D(\u_usb_host.u_phy.rx_dp0_q ),
    .RESET_B(net283),
    .Q(\u_usb_host.u_phy.rx_dp1_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._425_  (.CLK(clknet_4_10_0_usb_clk),
    .D(\u_usb_host.u_phy.rx_dn0_q ),
    .RESET_B(net283),
    .Q(\u_usb_host.u_phy.rx_dn1_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._426_  (.CLK(clknet_4_10_0_usb_clk),
    .D(net491),
    .RESET_B(net284),
    .Q(\u_usb_host.u_phy.rxd0_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._427_  (.CLK(clknet_4_10_0_usb_clk),
    .D(\u_usb_host.u_phy.rxd0_q ),
    .RESET_B(net283),
    .Q(\u_usb_host.u_phy.rxd1_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._428_  (.CLK(clknet_4_10_0_usb_clk),
    .D(\u_usb_host.u_phy.in_j_w ),
    .RESET_B(net281),
    .Q(\u_usb_host.u_phy.rxd_last_q ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._430_  (.CLK(clknet_4_10_0_usb_clk),
    .GATE(\u_usb_host.u_phy._021_ ),
    .GCLK(\u_usb_host.u_phy._173_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._432_  (.CLK(clknet_4_11_0_usb_clk),
    .GATE(\u_usb_host.u_phy._023_ ),
    .GCLK(\u_usb_host.u_phy._175_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._433_  (.CLK(clknet_4_10_0_usb_clk),
    .GATE(\u_usb_host.u_phy._024_ ),
    .GCLK(\u_usb_host.u_phy._176_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._434_  (.CLK(clknet_4_10_0_usb_clk),
    .GATE(\u_usb_host.u_phy._025_ ),
    .GCLK(\u_usb_host.u_phy._177_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._435_  (.CLK(clknet_4_10_0_usb_clk),
    .GATE(\u_usb_host.u_phy._026_ ),
    .GCLK(\u_usb_host.u_phy._178_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._436_  (.CLK(clknet_4_10_0_usb_clk),
    .GATE(\u_usb_host.u_phy._027_ ),
    .GCLK(\u_usb_host.u_phy._179_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_phy._437_  (.CLK(clknet_4_11_0_usb_clk),
    .GATE(\u_usb_host.u_phy._028_ ),
    .GCLK(\u_usb_host.u_phy._180_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._438_  (.CLK(clknet_4_11_0_usb_clk),
    .GATE(\u_usb_host.u_phy._029_ ),
    .GCLK(\u_usb_host.u_phy._181_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._439_  (.CLK(clknet_4_10_0_usb_clk),
    .GATE(\u_usb_host.u_phy._030_ ),
    .GCLK(\u_usb_host.u_phy._182_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._440_  (.CLK(clknet_4_11_0_usb_clk),
    .GATE(\u_usb_host.u_phy._031_ ),
    .GCLK(\u_usb_host.u_phy._183_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._441_  (.CLK(clknet_4_11_0_usb_clk),
    .GATE(\u_usb_host.u_phy._032_ ),
    .GCLK(\u_usb_host.u_phy._184_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._442_  (.CLK(clknet_4_11_0_usb_clk),
    .GATE(\u_usb_host.u_phy._033_ ),
    .GCLK(\u_usb_host.u_phy._185_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._443_  (.CLK(clknet_4_11_0_usb_clk),
    .GATE(\u_usb_host.u_phy._034_ ),
    .GCLK(\u_usb_host.u_phy._186_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._444_  (.CLK(clknet_4_11_0_usb_clk),
    .GATE(\u_usb_host.u_phy._035_ ),
    .GCLK(\u_usb_host.u_phy._187_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._445_  (.CLK(clknet_4_11_0_usb_clk),
    .GATE(\u_usb_host.u_phy._036_ ),
    .GCLK(\u_usb_host.u_phy._188_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._446_  (.CLK(clknet_4_10_0_usb_clk),
    .GATE(\u_usb_host.u_phy._037_ ),
    .GCLK(\u_usb_host.u_phy._189_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._447_  (.CLK(clknet_4_10_0_usb_clk),
    .GATE(\u_usb_host.u_phy._038_ ),
    .GCLK(\u_usb_host.u_phy._190_ ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_usb_rst._1_  (.CLK(clknet_4_0_0_usb_clk),
    .D(net378),
    .RESET_B(net46),
    .Q(\u_usb_host.u_usb_rst.in_data_s ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_usb_rst._1__378  (.HI(net378));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_usb_rst._2_  (.CLK(clknet_4_0_0_usb_clk),
    .D(net482),
    .RESET_B(net46),
    .Q(\u_usb_host.u_usb_rst.in_data_2s ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_usb_rst.u_buf.genblk1.u_mux  (.A0(net391),
    .A1(net46),
    .S(net323),
    .X(\u_usb_host.u_async_wb.u_cmd_if.rd_reset_n ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_usb_rst.u_buf.genblk1.u_mux_323  (.LO(net323));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_usb_xcvr._2_  (.A(\u_usb_host.u_phy.usb_tx_dn_o ),
    .Y(\u_usb_host.u_usb_xcvr._1_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_usb_xcvr._3_  (.A_N(net44),
    .B(net45),
    .X(\u_usb_host.u_phy.usb_rx_rcv_i ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_usb_xcvr._4_  (.A(\u_usb_host.u_phy.usb_tx_dp_o ),
    .B(net369),
    .Y(\u_usb_host.u_usb_xcvr._0_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_usb_xcvr._4__369  (.HI(net369));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_usb_xcvr._5_  (.A0(net370),
    .A1(\u_usb_host.u_usb_xcvr._0_ ),
    .S(\u_usb_host.u_usb_xcvr._1_ ),
    .X(net82));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_usb_xcvr._5__370  (.HI(net370));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_usb_xcvr._6_  (.A1(\u_usb_host.u_usb_xcvr._1_ ),
    .A2(net371),
    .B1(\u_usb_host.u_phy.usb_tx_dp_o ),
    .X(net83));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_usb_xcvr._6__371  (.HI(net371));
 sky130_fd_sc_hd__clkbuf_1 \u_usb_host.u_usb_xcvr._7_  (.A(\u_usb_host.u_phy.usb_tx_oen_o ),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 \u_usb_host.u_usb_xcvr._8_  (.A(net44),
    .X(\u_usb_host.u_phy.usb_rx_dn_i ));
 sky130_fd_sc_hd__clkbuf_1 \u_usb_host.u_usb_xcvr._9_  (.A(net45),
    .X(\u_usb_host.u_phy.usb_rx_dp_i ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_wb_rst._1_  (.CLK(clknet_1_0__leaf_app_clk),
    .D(net379),
    .RESET_B(net46),
    .Q(\u_usb_host.u_wb_rst.in_data_s ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_wb_rst._1__379  (.HI(net379));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_wb_rst._2_  (.CLK(clknet_1_0__leaf_app_clk),
    .D(net489),
    .RESET_B(net46),
    .Q(\u_usb_host.u_wb_rst.in_data_2s ));
 sky130_fd_sc_hd__mux2_2 \u_usb_host.u_wb_rst.u_buf.genblk1.u_mux  (.A0(net389),
    .A1(net46),
    .S(net324),
    .X(\u_usb_host.u_async_wb.u_cmd_if.wr_reset_n ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_wb_rst.u_buf.genblk1.u_mux_324  (.LO(net324));
 sky130_fd_sc_hd__buf_4 wire1 (.A(net381),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_2 wire2 (.A(usb_clk),
    .X(net381));
endmodule

