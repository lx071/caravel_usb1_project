// This is the unpowered netlist.
module wb_interconnect (clk_i,
    m0_wbd_ack_o,
    m0_wbd_cyc_i,
    m0_wbd_err_o,
    m0_wbd_lack_o,
    m0_wbd_stb_i,
    m0_wbd_we_i,
    m1_wbd_ack_o,
    m1_wbd_bry_i,
    m1_wbd_cyc_i,
    m1_wbd_err_o,
    m1_wbd_lack_o,
    m1_wbd_stb_i,
    m1_wbd_we_i,
    m2_wbd_ack_o,
    m2_wbd_bry_i,
    m2_wbd_cyc_i,
    m2_wbd_err_o,
    m2_wbd_lack_o,
    m2_wbd_stb_i,
    m2_wbd_we_i,
    m3_wbd_ack_o,
    m3_wbd_bry_i,
    m3_wbd_cyc_i,
    m3_wbd_err_o,
    m3_wbd_lack_o,
    m3_wbd_stb_i,
    m3_wbd_we_i,
    mclk_raw,
    peri_wbclk,
    riscv_wbclk,
    rst_n,
    s0_idle,
    s0_mclk,
    s0_wbd_ack_i,
    s0_wbd_bry_o,
    s0_wbd_cyc_o,
    s0_wbd_lack_i,
    s0_wbd_stb_o,
    s0_wbd_we_o,
    s1_mclk,
    s1_wbd_ack_i,
    s1_wbd_cyc_o,
    s1_wbd_stb_o,
    s1_wbd_we_o,
    s2_mclk,
    s2_wbd_ack_i,
    s2_wbd_cyc_o,
    s2_wbd_stb_o,
    s2_wbd_we_o,
    wbd_clk_int,
    wbd_clk_wi,
    cfg_cska_wi,
    ch_clk_in,
    ch_clk_out,
    ch_data_in,
    ch_data_out,
    m0_wbd_adr_i,
    m0_wbd_dat_i,
    m0_wbd_dat_o,
    m0_wbd_sel_i,
    m1_wbd_adr_i,
    m1_wbd_bl_i,
    m1_wbd_dat_i,
    m1_wbd_dat_o,
    m1_wbd_sel_i,
    m2_wbd_adr_i,
    m2_wbd_bl_i,
    m2_wbd_dat_i,
    m2_wbd_dat_o,
    m2_wbd_sel_i,
    m3_wbd_adr_i,
    m3_wbd_bl_i,
    m3_wbd_dat_o,
    m3_wbd_sel_i,
    s0_wbd_adr_o,
    s0_wbd_bl_o,
    s0_wbd_dat_i,
    s0_wbd_dat_o,
    s0_wbd_sel_o,
    s1_wbd_adr_o,
    s1_wbd_dat_i,
    s1_wbd_dat_o,
    s1_wbd_sel_o,
    s2_wbd_adr_o,
    s2_wbd_dat_i,
    s2_wbd_dat_o,
    s2_wbd_sel_o);
 input clk_i;
 output m0_wbd_ack_o;
 input m0_wbd_cyc_i;
 output m0_wbd_err_o;
 output m0_wbd_lack_o;
 input m0_wbd_stb_i;
 input m0_wbd_we_i;
 output m1_wbd_ack_o;
 input m1_wbd_bry_i;
 input m1_wbd_cyc_i;
 output m1_wbd_err_o;
 output m1_wbd_lack_o;
 input m1_wbd_stb_i;
 input m1_wbd_we_i;
 output m2_wbd_ack_o;
 input m2_wbd_bry_i;
 input m2_wbd_cyc_i;
 output m2_wbd_err_o;
 output m2_wbd_lack_o;
 input m2_wbd_stb_i;
 input m2_wbd_we_i;
 output m3_wbd_ack_o;
 input m3_wbd_bry_i;
 input m3_wbd_cyc_i;
 output m3_wbd_err_o;
 output m3_wbd_lack_o;
 input m3_wbd_stb_i;
 input m3_wbd_we_i;
 input mclk_raw;
 output peri_wbclk;
 output riscv_wbclk;
 input rst_n;
 input s0_idle;
 output s0_mclk;
 input s0_wbd_ack_i;
 output s0_wbd_bry_o;
 output s0_wbd_cyc_o;
 input s0_wbd_lack_i;
 output s0_wbd_stb_o;
 output s0_wbd_we_o;
 output s1_mclk;
 input s1_wbd_ack_i;
 output s1_wbd_cyc_o;
 output s1_wbd_stb_o;
 output s1_wbd_we_o;
 output s2_mclk;
 input s2_wbd_ack_i;
 output s2_wbd_cyc_o;
 output s2_wbd_stb_o;
 output s2_wbd_we_o;
 input wbd_clk_int;
 output wbd_clk_wi;
 input [3:0] cfg_cska_wi;
 input [2:0] ch_clk_in;
 output [2:0] ch_clk_out;
 input [157:0] ch_data_in;
 output [157:0] ch_data_out;
 input [31:0] m0_wbd_adr_i;
 input [31:0] m0_wbd_dat_i;
 output [31:0] m0_wbd_dat_o;
 input [3:0] m0_wbd_sel_i;
 input [31:0] m1_wbd_adr_i;
 input [2:0] m1_wbd_bl_i;
 input [31:0] m1_wbd_dat_i;
 output [31:0] m1_wbd_dat_o;
 input [3:0] m1_wbd_sel_i;
 input [31:0] m2_wbd_adr_i;
 input [9:0] m2_wbd_bl_i;
 input [31:0] m2_wbd_dat_i;
 output [31:0] m2_wbd_dat_o;
 input [3:0] m2_wbd_sel_i;
 input [31:0] m3_wbd_adr_i;
 input [9:0] m3_wbd_bl_i;
 output [31:0] m3_wbd_dat_o;
 input [3:0] m3_wbd_sel_i;
 output [31:0] s0_wbd_adr_o;
 output [9:0] s0_wbd_bl_o;
 input [31:0] s0_wbd_dat_i;
 output [31:0] s0_wbd_dat_o;
 output [3:0] s0_wbd_sel_o;
 output [8:0] s1_wbd_adr_o;
 input [31:0] s1_wbd_dat_i;
 output [31:0] s1_wbd_dat_o;
 output [3:0] s1_wbd_sel_o;
 output [10:0] s2_wbd_adr_o;
 input [31:0] s2_wbd_dat_i;
 output [31:0] s2_wbd_dat_o;
 output [3:0] s2_wbd_sel_o;

 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire clknet_0_mclk_raw;
 wire \clknet_0_u_dsync.out_clk ;
 wire clknet_1_0_0_mclk_raw;
 wire \clknet_1_0_0_u_dsync.out_clk ;
 wire clknet_1_1_0_mclk_raw;
 wire \clknet_1_1_0_u_dsync.out_clk ;
 wire clknet_2_0__leaf_mclk_raw;
 wire clknet_2_1__leaf_mclk_raw;
 wire clknet_2_2__leaf_mclk_raw;
 wire clknet_2_3__leaf_mclk_raw;
 wire \clknet_3_0__leaf_u_dsync.out_clk ;
 wire \clknet_3_1__leaf_u_dsync.out_clk ;
 wire \clknet_3_2__leaf_u_dsync.out_clk ;
 wire \clknet_3_3__leaf_u_dsync.out_clk ;
 wire \clknet_3_4__leaf_u_dsync.out_clk ;
 wire \clknet_3_5__leaf_u_dsync.out_clk ;
 wire \clknet_3_6__leaf_u_dsync.out_clk ;
 wire \clknet_3_7__leaf_u_dsync.out_clk ;
 wire \clknet_leaf_0_u_dsync.out_clk ;
 wire \clknet_leaf_100_u_dsync.out_clk ;
 wire \clknet_leaf_101_u_dsync.out_clk ;
 wire \clknet_leaf_102_u_dsync.out_clk ;
 wire \clknet_leaf_103_u_dsync.out_clk ;
 wire \clknet_leaf_104_u_dsync.out_clk ;
 wire \clknet_leaf_105_u_dsync.out_clk ;
 wire \clknet_leaf_106_u_dsync.out_clk ;
 wire \clknet_leaf_107_u_dsync.out_clk ;
 wire \clknet_leaf_108_u_dsync.out_clk ;
 wire \clknet_leaf_109_u_dsync.out_clk ;
 wire \clknet_leaf_10_u_dsync.out_clk ;
 wire \clknet_leaf_11_u_dsync.out_clk ;
 wire \clknet_leaf_12_u_dsync.out_clk ;
 wire \clknet_leaf_13_u_dsync.out_clk ;
 wire \clknet_leaf_14_u_dsync.out_clk ;
 wire \clknet_leaf_15_u_dsync.out_clk ;
 wire \clknet_leaf_16_u_dsync.out_clk ;
 wire \clknet_leaf_17_u_dsync.out_clk ;
 wire \clknet_leaf_18_u_dsync.out_clk ;
 wire \clknet_leaf_19_u_dsync.out_clk ;
 wire \clknet_leaf_1_u_dsync.out_clk ;
 wire \clknet_leaf_20_u_dsync.out_clk ;
 wire \clknet_leaf_21_u_dsync.out_clk ;
 wire \clknet_leaf_22_u_dsync.out_clk ;
 wire \clknet_leaf_23_u_dsync.out_clk ;
 wire \clknet_leaf_24_u_dsync.out_clk ;
 wire \clknet_leaf_25_u_dsync.out_clk ;
 wire \clknet_leaf_26_u_dsync.out_clk ;
 wire \clknet_leaf_27_u_dsync.out_clk ;
 wire \clknet_leaf_28_u_dsync.out_clk ;
 wire \clknet_leaf_29_u_dsync.out_clk ;
 wire \clknet_leaf_2_u_dsync.out_clk ;
 wire \clknet_leaf_30_u_dsync.out_clk ;
 wire \clknet_leaf_31_u_dsync.out_clk ;
 wire \clknet_leaf_32_u_dsync.out_clk ;
 wire \clknet_leaf_33_u_dsync.out_clk ;
 wire \clknet_leaf_34_u_dsync.out_clk ;
 wire \clknet_leaf_35_u_dsync.out_clk ;
 wire \clknet_leaf_36_u_dsync.out_clk ;
 wire \clknet_leaf_37_u_dsync.out_clk ;
 wire \clknet_leaf_38_u_dsync.out_clk ;
 wire \clknet_leaf_39_u_dsync.out_clk ;
 wire \clknet_leaf_3_u_dsync.out_clk ;
 wire \clknet_leaf_40_u_dsync.out_clk ;
 wire \clknet_leaf_41_u_dsync.out_clk ;
 wire \clknet_leaf_42_u_dsync.out_clk ;
 wire \clknet_leaf_43_u_dsync.out_clk ;
 wire \clknet_leaf_44_u_dsync.out_clk ;
 wire \clknet_leaf_45_u_dsync.out_clk ;
 wire \clknet_leaf_46_u_dsync.out_clk ;
 wire \clknet_leaf_47_u_dsync.out_clk ;
 wire \clknet_leaf_48_u_dsync.out_clk ;
 wire \clknet_leaf_49_u_dsync.out_clk ;
 wire \clknet_leaf_4_u_dsync.out_clk ;
 wire \clknet_leaf_50_u_dsync.out_clk ;
 wire \clknet_leaf_51_u_dsync.out_clk ;
 wire \clknet_leaf_52_u_dsync.out_clk ;
 wire \clknet_leaf_53_u_dsync.out_clk ;
 wire \clknet_leaf_54_u_dsync.out_clk ;
 wire \clknet_leaf_55_u_dsync.out_clk ;
 wire \clknet_leaf_56_u_dsync.out_clk ;
 wire \clknet_leaf_57_u_dsync.out_clk ;
 wire \clknet_leaf_58_u_dsync.out_clk ;
 wire \clknet_leaf_59_u_dsync.out_clk ;
 wire \clknet_leaf_5_u_dsync.out_clk ;
 wire \clknet_leaf_60_u_dsync.out_clk ;
 wire \clknet_leaf_61_u_dsync.out_clk ;
 wire \clknet_leaf_62_u_dsync.out_clk ;
 wire \clknet_leaf_63_u_dsync.out_clk ;
 wire \clknet_leaf_64_u_dsync.out_clk ;
 wire \clknet_leaf_65_u_dsync.out_clk ;
 wire \clknet_leaf_66_u_dsync.out_clk ;
 wire \clknet_leaf_67_u_dsync.out_clk ;
 wire \clknet_leaf_68_u_dsync.out_clk ;
 wire \clknet_leaf_69_u_dsync.out_clk ;
 wire \clknet_leaf_6_u_dsync.out_clk ;
 wire \clknet_leaf_70_u_dsync.out_clk ;
 wire \clknet_leaf_71_u_dsync.out_clk ;
 wire \clknet_leaf_72_u_dsync.out_clk ;
 wire \clknet_leaf_73_u_dsync.out_clk ;
 wire \clknet_leaf_74_u_dsync.out_clk ;
 wire \clknet_leaf_75_u_dsync.out_clk ;
 wire \clknet_leaf_76_u_dsync.out_clk ;
 wire \clknet_leaf_77_u_dsync.out_clk ;
 wire \clknet_leaf_78_u_dsync.out_clk ;
 wire \clknet_leaf_79_u_dsync.out_clk ;
 wire \clknet_leaf_7_u_dsync.out_clk ;
 wire \clknet_leaf_80_u_dsync.out_clk ;
 wire \clknet_leaf_81_u_dsync.out_clk ;
 wire \clknet_leaf_82_u_dsync.out_clk ;
 wire \clknet_leaf_83_u_dsync.out_clk ;
 wire \clknet_leaf_84_u_dsync.out_clk ;
 wire \clknet_leaf_85_u_dsync.out_clk ;
 wire \clknet_leaf_86_u_dsync.out_clk ;
 wire \clknet_leaf_87_u_dsync.out_clk ;
 wire \clknet_leaf_88_u_dsync.out_clk ;
 wire \clknet_leaf_89_u_dsync.out_clk ;
 wire \clknet_leaf_8_u_dsync.out_clk ;
 wire \clknet_leaf_90_u_dsync.out_clk ;
 wire \clknet_leaf_91_u_dsync.out_clk ;
 wire \clknet_leaf_92_u_dsync.out_clk ;
 wire \clknet_leaf_93_u_dsync.out_clk ;
 wire \clknet_leaf_94_u_dsync.out_clk ;
 wire \clknet_leaf_95_u_dsync.out_clk ;
 wire \clknet_leaf_96_u_dsync.out_clk ;
 wire \clknet_leaf_97_u_dsync.out_clk ;
 wire \clknet_leaf_98_u_dsync.out_clk ;
 wire \clknet_leaf_99_u_dsync.out_clk ;
 wire \clknet_leaf_9_u_dsync.out_clk ;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net127;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net128;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net129;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net130;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net131;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net132;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net133;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net134;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net135;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net136;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net137;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net138;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net139;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net14;
 wire net140;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net141;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net142;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net143;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net144;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net145;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net146;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net147;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net148;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net149;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net15;
 wire net150;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net151;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net152;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net153;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net154;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net155;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net156;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net157;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net158;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net159;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net16;
 wire net160;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net161;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net162;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net163;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net164;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net165;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net166;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net167;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net168;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net169;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net17;
 wire net170;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net171;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net172;
 wire net1720;
 wire net173;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net174;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net175;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net176;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net177;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1779;
 wire net178;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net179;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net18;
 wire net180;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net181;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net182;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net183;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net184;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net185;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net186;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net187;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net188;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net189;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net19;
 wire net190;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net191;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net192;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net193;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net194;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net195;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net196;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net197;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net198;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net199;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2;
 wire net20;
 wire net200;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net201;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net202;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net203;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net204;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net205;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net206;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net207;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net208;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net209;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire \u_dcg_peri.cfg_mode[0] ;
 wire \u_dcg_peri.cfg_mode[1] ;
 wire \u_dcg_peri.cfg_mode_ss[0] ;
 wire \u_dcg_peri.cfg_mode_ss[1] ;
 wire \u_dcg_peri.clk_enb ;
 wire \u_dcg_peri.reset_n ;
 wire \u_dcg_peri.u_dsync.in_data_2s[0] ;
 wire \u_dcg_peri.u_dsync.in_data_2s[1] ;
 wire \u_dcg_peri.u_dsync.in_data_s[0] ;
 wire \u_dcg_peri.u_dsync.in_data_s[1] ;
 wire \u_dcg_riscv.cfg_mode[0] ;
 wire \u_dcg_riscv.cfg_mode[1] ;
 wire \u_dcg_riscv.cfg_mode_ss[0] ;
 wire \u_dcg_riscv.cfg_mode_ss[1] ;
 wire \u_dcg_riscv.clk_enb ;
 wire \u_dcg_riscv.u_dsync.in_data_2s[0] ;
 wire \u_dcg_riscv.u_dsync.in_data_2s[1] ;
 wire \u_dcg_riscv.u_dsync.in_data_s[0] ;
 wire \u_dcg_riscv.u_dsync.in_data_s[1] ;
 wire \u_dcg_s0.cfg_mode[0] ;
 wire \u_dcg_s0.cfg_mode[1] ;
 wire \u_dcg_s0.cfg_mode_ss[0] ;
 wire \u_dcg_s0.cfg_mode_ss[1] ;
 wire \u_dcg_s0.clk_enb ;
 wire \u_dcg_s0.dst_idle_r ;
 wire \u_dcg_s0.hcnt[0] ;
 wire \u_dcg_s0.hcnt[1] ;
 wire \u_dcg_s0.hcnt[2] ;
 wire \u_dcg_s0.hcnt[3] ;
 wire \u_dcg_s0.idle_his ;
 wire \u_dcg_s0.u_dsync.in_data_2s[0] ;
 wire \u_dcg_s0.u_dsync.in_data_2s[1] ;
 wire \u_dcg_s0.u_dsync.in_data_s[0] ;
 wire \u_dcg_s0.u_dsync.in_data_s[1] ;
 wire \u_dcg_s1.cfg_mode[0] ;
 wire \u_dcg_s1.cfg_mode[1] ;
 wire \u_dcg_s1.cfg_mode_ss[0] ;
 wire \u_dcg_s1.cfg_mode_ss[1] ;
 wire \u_dcg_s1.clk_enb ;
 wire \u_dcg_s1.u_dsync.in_data_2s[0] ;
 wire \u_dcg_s1.u_dsync.in_data_2s[1] ;
 wire \u_dcg_s1.u_dsync.in_data_s[0] ;
 wire \u_dcg_s1.u_dsync.in_data_s[1] ;
 wire \u_dcg_s2.cfg_mode[0] ;
 wire \u_dcg_s2.cfg_mode[1] ;
 wire \u_dcg_s2.cfg_mode_ss[0] ;
 wire \u_dcg_s2.cfg_mode_ss[1] ;
 wire \u_dcg_s2.clk_enb ;
 wire \u_dcg_s2.u_dsync.in_data_2s[0] ;
 wire \u_dcg_s2.u_dsync.in_data_2s[1] ;
 wire \u_dcg_s2.u_dsync.in_data_s[0] ;
 wire \u_dcg_s2.u_dsync.in_data_s[1] ;
 wire \u_dsync.in_data_2s[0] ;
 wire \u_dsync.in_data_2s[1] ;
 wire \u_dsync.in_data_2s[2] ;
 wire \u_dsync.in_data_2s[3] ;
 wire \u_dsync.in_data_2s[4] ;
 wire \u_dsync.in_data_2s[5] ;
 wire \u_dsync.in_data_2s[6] ;
 wire \u_dsync.in_data_2s[7] ;
 wire \u_dsync.in_data_s[0] ;
 wire \u_dsync.in_data_s[1] ;
 wire \u_dsync.in_data_s[2] ;
 wire \u_dsync.in_data_s[3] ;
 wire \u_dsync.in_data_s[4] ;
 wire \u_dsync.in_data_s[5] ;
 wire \u_dsync.in_data_s[6] ;
 wire \u_dsync.in_data_s[7] ;
 wire \u_dsync.out_clk ;
 wire \u_dsync.out_data[0] ;
 wire \u_dsync.out_data[1] ;
 wire \u_dsync.out_data[2] ;
 wire \u_dsync.out_data[3] ;
 wire \u_dsync.out_data[4] ;
 wire \u_dsync.out_data[5] ;
 wire \u_dsync.out_data[6] ;
 wire \u_dsync.out_data[7] ;
 wire \u_reg.cfg_dcg_ctrl[10] ;
 wire \u_reg.cfg_dcg_ctrl[11] ;
 wire \u_reg.cfg_dcg_ctrl[12] ;
 wire \u_reg.cfg_dcg_ctrl[13] ;
 wire \u_reg.cfg_dcg_ctrl[14] ;
 wire \u_reg.cfg_dcg_ctrl[15] ;
 wire \u_reg.cfg_dcg_ctrl[16] ;
 wire \u_reg.cfg_dcg_ctrl[17] ;
 wire \u_reg.cfg_dcg_ctrl[18] ;
 wire \u_reg.cfg_dcg_ctrl[19] ;
 wire \u_reg.cfg_dcg_ctrl[20] ;
 wire \u_reg.cfg_dcg_ctrl[21] ;
 wire \u_reg.cfg_dcg_ctrl[22] ;
 wire \u_reg.cfg_dcg_ctrl[23] ;
 wire \u_reg.cfg_dcg_ctrl[24] ;
 wire \u_reg.cfg_dcg_ctrl[25] ;
 wire \u_reg.cfg_dcg_ctrl[26] ;
 wire \u_reg.cfg_dcg_ctrl[27] ;
 wire \u_reg.cfg_dcg_ctrl[28] ;
 wire \u_reg.cfg_dcg_ctrl[29] ;
 wire \u_reg.cfg_dcg_ctrl[30] ;
 wire \u_reg.cfg_dcg_ctrl[31] ;
 wire \u_reg.reg_2[0] ;
 wire \u_reg.reg_2[10] ;
 wire \u_reg.reg_2[11] ;
 wire \u_reg.reg_2[12] ;
 wire \u_reg.reg_2[13] ;
 wire \u_reg.reg_2[14] ;
 wire \u_reg.reg_2[15] ;
 wire \u_reg.reg_2[16] ;
 wire \u_reg.reg_2[17] ;
 wire \u_reg.reg_2[18] ;
 wire \u_reg.reg_2[19] ;
 wire \u_reg.reg_2[1] ;
 wire \u_reg.reg_2[20] ;
 wire \u_reg.reg_2[21] ;
 wire \u_reg.reg_2[22] ;
 wire \u_reg.reg_2[23] ;
 wire \u_reg.reg_2[24] ;
 wire \u_reg.reg_2[25] ;
 wire \u_reg.reg_2[26] ;
 wire \u_reg.reg_2[27] ;
 wire \u_reg.reg_2[28] ;
 wire \u_reg.reg_2[29] ;
 wire \u_reg.reg_2[2] ;
 wire \u_reg.reg_2[30] ;
 wire \u_reg.reg_2[31] ;
 wire \u_reg.reg_2[3] ;
 wire \u_reg.reg_2[4] ;
 wire \u_reg.reg_2[5] ;
 wire \u_reg.reg_2[6] ;
 wire \u_reg.reg_2[7] ;
 wire \u_reg.reg_2[8] ;
 wire \u_reg.reg_2[9] ;
 wire \u_reg.reg_3[0] ;
 wire \u_reg.reg_3[10] ;
 wire \u_reg.reg_3[11] ;
 wire \u_reg.reg_3[12] ;
 wire \u_reg.reg_3[13] ;
 wire \u_reg.reg_3[14] ;
 wire \u_reg.reg_3[15] ;
 wire \u_reg.reg_3[16] ;
 wire \u_reg.reg_3[17] ;
 wire \u_reg.reg_3[18] ;
 wire \u_reg.reg_3[19] ;
 wire \u_reg.reg_3[1] ;
 wire \u_reg.reg_3[20] ;
 wire \u_reg.reg_3[21] ;
 wire \u_reg.reg_3[22] ;
 wire \u_reg.reg_3[23] ;
 wire \u_reg.reg_3[24] ;
 wire \u_reg.reg_3[25] ;
 wire \u_reg.reg_3[26] ;
 wire \u_reg.reg_3[27] ;
 wire \u_reg.reg_3[28] ;
 wire \u_reg.reg_3[29] ;
 wire \u_reg.reg_3[2] ;
 wire \u_reg.reg_3[30] ;
 wire \u_reg.reg_3[31] ;
 wire \u_reg.reg_3[3] ;
 wire \u_reg.reg_3[4] ;
 wire \u_reg.reg_3[5] ;
 wire \u_reg.reg_3[6] ;
 wire \u_reg.reg_3[7] ;
 wire \u_reg.reg_3[8] ;
 wire \u_reg.reg_3[9] ;
 wire \u_reg.reg_4[0] ;
 wire \u_reg.reg_4[10] ;
 wire \u_reg.reg_4[11] ;
 wire \u_reg.reg_4[12] ;
 wire \u_reg.reg_4[13] ;
 wire \u_reg.reg_4[14] ;
 wire \u_reg.reg_4[15] ;
 wire \u_reg.reg_4[16] ;
 wire \u_reg.reg_4[17] ;
 wire \u_reg.reg_4[18] ;
 wire \u_reg.reg_4[19] ;
 wire \u_reg.reg_4[1] ;
 wire \u_reg.reg_4[20] ;
 wire \u_reg.reg_4[21] ;
 wire \u_reg.reg_4[22] ;
 wire \u_reg.reg_4[23] ;
 wire \u_reg.reg_4[24] ;
 wire \u_reg.reg_4[25] ;
 wire \u_reg.reg_4[26] ;
 wire \u_reg.reg_4[27] ;
 wire \u_reg.reg_4[28] ;
 wire \u_reg.reg_4[29] ;
 wire \u_reg.reg_4[2] ;
 wire \u_reg.reg_4[30] ;
 wire \u_reg.reg_4[31] ;
 wire \u_reg.reg_4[3] ;
 wire \u_reg.reg_4[4] ;
 wire \u_reg.reg_4[5] ;
 wire \u_reg.reg_4[6] ;
 wire \u_reg.reg_4[7] ;
 wire \u_reg.reg_4[8] ;
 wire \u_reg.reg_4[9] ;
 wire \u_reg.reg_5[0] ;
 wire \u_reg.reg_5[10] ;
 wire \u_reg.reg_5[11] ;
 wire \u_reg.reg_5[12] ;
 wire \u_reg.reg_5[13] ;
 wire \u_reg.reg_5[14] ;
 wire \u_reg.reg_5[15] ;
 wire \u_reg.reg_5[16] ;
 wire \u_reg.reg_5[17] ;
 wire \u_reg.reg_5[18] ;
 wire \u_reg.reg_5[19] ;
 wire \u_reg.reg_5[1] ;
 wire \u_reg.reg_5[20] ;
 wire \u_reg.reg_5[21] ;
 wire \u_reg.reg_5[22] ;
 wire \u_reg.reg_5[23] ;
 wire \u_reg.reg_5[24] ;
 wire \u_reg.reg_5[25] ;
 wire \u_reg.reg_5[26] ;
 wire \u_reg.reg_5[27] ;
 wire \u_reg.reg_5[28] ;
 wire \u_reg.reg_5[29] ;
 wire \u_reg.reg_5[2] ;
 wire \u_reg.reg_5[30] ;
 wire \u_reg.reg_5[31] ;
 wire \u_reg.reg_5[3] ;
 wire \u_reg.reg_5[4] ;
 wire \u_reg.reg_5[5] ;
 wire \u_reg.reg_5[6] ;
 wire \u_reg.reg_5[7] ;
 wire \u_reg.reg_5[8] ;
 wire \u_reg.reg_5[9] ;
 wire \u_reg.reg_6[0] ;
 wire \u_reg.reg_6[10] ;
 wire \u_reg.reg_6[11] ;
 wire \u_reg.reg_6[12] ;
 wire \u_reg.reg_6[13] ;
 wire \u_reg.reg_6[14] ;
 wire \u_reg.reg_6[15] ;
 wire \u_reg.reg_6[16] ;
 wire \u_reg.reg_6[17] ;
 wire \u_reg.reg_6[18] ;
 wire \u_reg.reg_6[19] ;
 wire \u_reg.reg_6[1] ;
 wire \u_reg.reg_6[20] ;
 wire \u_reg.reg_6[21] ;
 wire \u_reg.reg_6[22] ;
 wire \u_reg.reg_6[23] ;
 wire \u_reg.reg_6[24] ;
 wire \u_reg.reg_6[25] ;
 wire \u_reg.reg_6[26] ;
 wire \u_reg.reg_6[27] ;
 wire \u_reg.reg_6[28] ;
 wire \u_reg.reg_6[29] ;
 wire \u_reg.reg_6[2] ;
 wire \u_reg.reg_6[30] ;
 wire \u_reg.reg_6[31] ;
 wire \u_reg.reg_6[3] ;
 wire \u_reg.reg_6[4] ;
 wire \u_reg.reg_6[5] ;
 wire \u_reg.reg_6[6] ;
 wire \u_reg.reg_6[7] ;
 wire \u_reg.reg_6[8] ;
 wire \u_reg.reg_6[9] ;
 wire \u_reg.reg_7[0] ;
 wire \u_reg.reg_7[10] ;
 wire \u_reg.reg_7[11] ;
 wire \u_reg.reg_7[12] ;
 wire \u_reg.reg_7[13] ;
 wire \u_reg.reg_7[14] ;
 wire \u_reg.reg_7[15] ;
 wire \u_reg.reg_7[16] ;
 wire \u_reg.reg_7[17] ;
 wire \u_reg.reg_7[18] ;
 wire \u_reg.reg_7[19] ;
 wire \u_reg.reg_7[1] ;
 wire \u_reg.reg_7[20] ;
 wire \u_reg.reg_7[21] ;
 wire \u_reg.reg_7[22] ;
 wire \u_reg.reg_7[23] ;
 wire \u_reg.reg_7[24] ;
 wire \u_reg.reg_7[25] ;
 wire \u_reg.reg_7[26] ;
 wire \u_reg.reg_7[27] ;
 wire \u_reg.reg_7[28] ;
 wire \u_reg.reg_7[29] ;
 wire \u_reg.reg_7[2] ;
 wire \u_reg.reg_7[30] ;
 wire \u_reg.reg_7[31] ;
 wire \u_reg.reg_7[3] ;
 wire \u_reg.reg_7[4] ;
 wire \u_reg.reg_7[5] ;
 wire \u_reg.reg_7[6] ;
 wire \u_reg.reg_7[7] ;
 wire \u_reg.reg_7[8] ;
 wire \u_reg.reg_7[9] ;
 wire \u_reg.reg_ack ;
 wire \u_reg.reg_rdata[0] ;
 wire \u_reg.reg_rdata[10] ;
 wire \u_reg.reg_rdata[11] ;
 wire \u_reg.reg_rdata[12] ;
 wire \u_reg.reg_rdata[13] ;
 wire \u_reg.reg_rdata[14] ;
 wire \u_reg.reg_rdata[15] ;
 wire \u_reg.reg_rdata[16] ;
 wire \u_reg.reg_rdata[17] ;
 wire \u_reg.reg_rdata[18] ;
 wire \u_reg.reg_rdata[19] ;
 wire \u_reg.reg_rdata[1] ;
 wire \u_reg.reg_rdata[20] ;
 wire \u_reg.reg_rdata[21] ;
 wire \u_reg.reg_rdata[22] ;
 wire \u_reg.reg_rdata[23] ;
 wire \u_reg.reg_rdata[24] ;
 wire \u_reg.reg_rdata[25] ;
 wire \u_reg.reg_rdata[26] ;
 wire \u_reg.reg_rdata[27] ;
 wire \u_reg.reg_rdata[28] ;
 wire \u_reg.reg_rdata[29] ;
 wire \u_reg.reg_rdata[2] ;
 wire \u_reg.reg_rdata[30] ;
 wire \u_reg.reg_rdata[31] ;
 wire \u_reg.reg_rdata[3] ;
 wire \u_reg.reg_rdata[4] ;
 wire \u_reg.reg_rdata[5] ;
 wire \u_reg.reg_rdata[6] ;
 wire \u_reg.reg_rdata[7] ;
 wire \u_reg.reg_rdata[8] ;
 wire \u_reg.reg_rdata[9] ;
 wire \u_rst_sync.in_data_2s ;
 wire \u_rst_sync.in_data_s ;
 wire \u_s0.gnt[0] ;
 wire \u_s0.gnt[1] ;
 wire \u_s0.u_sync_wbb.m_bl_cnt[0] ;
 wire \u_s0.u_sync_wbb.m_bl_cnt[1] ;
 wire \u_s0.u_sync_wbb.m_bl_cnt[2] ;
 wire \u_s0.u_sync_wbb.m_bl_cnt[3] ;
 wire \u_s0.u_sync_wbb.m_bl_cnt[4] ;
 wire \u_s0.u_sync_wbb.m_bl_cnt[5] ;
 wire \u_s0.u_sync_wbb.m_bl_cnt[6] ;
 wire \u_s0.u_sync_wbb.m_bl_cnt[7] ;
 wire \u_s0.u_sync_wbb.m_bl_cnt[8] ;
 wire \u_s0.u_sync_wbb.m_bl_cnt[9] ;
 wire \u_s0.u_sync_wbb.m_cmd_wr_en ;
 wire \u_s0.u_sync_wbb.m_resp_rd_en ;
 wire \u_s0.u_sync_wbb.m_state[0] ;
 wire \u_s0.u_sync_wbb.m_state[1] ;
 wire \u_s0.u_sync_wbb.m_state[2] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[0] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[14] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[15] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[16] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[17] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[18] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[19] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[1] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[20] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[21] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[22] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[23] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[24] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[25] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[26] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[27] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[28] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[29] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[2] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[30] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[31] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[32] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[33] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[34] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[35] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[36] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[37] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[38] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[39] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[3] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[40] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[41] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[42] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[43] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[44] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[45] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[46] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[47] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[48] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[49] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[4] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[50] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[53] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[54] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[55] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[56] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[57] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[58] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[59] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[5] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[60] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[61] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[62] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[63] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[64] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[65] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[66] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[67] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[68] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[69] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[6] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[70] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[71] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[72] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[73] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[74] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[75] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[76] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[77] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[78] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[79] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[7] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[80] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[81] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[82] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[8] ;
 wire \u_s0.u_sync_wbb.s_cmd_rd_data_l[9] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][0] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][14] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][15] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][16] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][17] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][18] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][19] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][1] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][20] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][21] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][22] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][23] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][24] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][25] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][26] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][27] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][28] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][29] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][2] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][30] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][31] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][32] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][33] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][34] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][35] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][36] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][37] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][38] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][39] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][3] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][40] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][41] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][42] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][43] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][44] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][45] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][46] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][47] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][48] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][49] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][4] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][50] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][53] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][54] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][55] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][56] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][57] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][58] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][59] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][5] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][60] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][61] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][62] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][63] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][64] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][65] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][66] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][67] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][68] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][69] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][6] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][70] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][71] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][72] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][73] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][74] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][75] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][76] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][77] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][78] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][79] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][7] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][80] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][81] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][82] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][8] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[0][9] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][0] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][14] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][15] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][16] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][17] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][18] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][19] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][1] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][20] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][21] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][22] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][23] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][24] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][25] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][26] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][27] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][28] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][29] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][2] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][30] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][31] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][32] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][33] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][34] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][35] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][36] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][37] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][38] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][39] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][3] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][40] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][41] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][42] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][43] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][44] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][45] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][46] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][47] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][48] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][49] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][4] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][50] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][53] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][54] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][55] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][56] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][57] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][58] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][59] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][5] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][60] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][61] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][62] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][63] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][64] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][65] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][66] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][67] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][68] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][69] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][6] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][70] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][71] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][72] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][73] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][74] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][75] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][76] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][77] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][78] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][79] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][7] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][80] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][81] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][82] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][8] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[1][9] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][0] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][14] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][15] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][16] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][17] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][18] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][19] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][1] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][20] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][21] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][22] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][23] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][24] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][25] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][26] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][27] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][28] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][29] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][2] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][30] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][31] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][32] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][33] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][34] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][35] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][36] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][37] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][38] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][39] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][3] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][40] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][41] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][42] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][43] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][44] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][45] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][46] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][47] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][48] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][49] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][4] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][50] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][53] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][54] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][55] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][56] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][57] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][58] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][59] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][5] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][60] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][61] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][62] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][63] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][64] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][65] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][66] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][67] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][68] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][69] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][6] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][70] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][71] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][72] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][73] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][74] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][75] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][76] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][77] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][78] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][79] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][7] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][80] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][81] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][82] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][8] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[2][9] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][0] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][14] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][15] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][16] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][17] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][18] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][19] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][1] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][20] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][21] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][22] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][23] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][24] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][25] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][26] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][27] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][28] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][29] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][2] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][30] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][31] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][32] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][33] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][34] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][35] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][36] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][37] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][38] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][39] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][3] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][40] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][41] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][42] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][43] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][44] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][45] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][46] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][47] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][48] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][49] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][4] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][50] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][53] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][54] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][55] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][56] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][57] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][58] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][59] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][5] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][60] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][61] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][62] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][63] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][64] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][65] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][66] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][67] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][68] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][69] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][6] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][70] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][71] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][72] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][73] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][74] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][75] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][76] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][77] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][78] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][79] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][7] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][80] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][81] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][82] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][8] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.mem[3][9] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.rd_ptr[0] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.rd_ptr[1] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.rd_ptr[2] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.wr_ptr[0] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.wr_ptr[1] ;
 wire \u_s0.u_sync_wbb.u_cmd_if.wr_ptr[2] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][0] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][10] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][11] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][12] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][13] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][14] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][15] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][16] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][17] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][18] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][19] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][1] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][20] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][21] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][22] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][23] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][24] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][25] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][26] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][27] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][28] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][29] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][2] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][30] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][31] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][3] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][4] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][5] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][6] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][7] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][8] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[0][9] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][0] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][10] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][11] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][12] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][13] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][14] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][15] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][16] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][17] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][18] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][19] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][1] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][20] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][21] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][22] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][23] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][24] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][25] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][26] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][27] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][28] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][29] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][2] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][30] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][31] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][3] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][4] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][5] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][6] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][7] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][8] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[1][9] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][0] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][10] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][11] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][12] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][13] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][14] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][15] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][16] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][17] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][18] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][19] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][1] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][20] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][21] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][22] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][23] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][24] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][25] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][26] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][27] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][28] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][29] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][2] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][30] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][31] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][3] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][4] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][5] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][6] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][7] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][8] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[2][9] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][0] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][10] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][11] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][12] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][13] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][14] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][15] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][16] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][17] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][18] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][19] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][1] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][20] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][21] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][22] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][23] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][24] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][25] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][26] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][27] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][28] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][29] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][2] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][30] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][31] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][3] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][4] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][5] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][6] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][7] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][8] ;
 wire \u_s0.u_sync_wbb.u_resp_if.mem[3][9] ;
 wire \u_s0.u_sync_wbb.u_resp_if.rd_ptr[0] ;
 wire \u_s0.u_sync_wbb.u_resp_if.rd_ptr[1] ;
 wire \u_s0.u_sync_wbb.u_resp_if.rd_ptr[2] ;
 wire \u_s0.u_sync_wbb.u_resp_if.wr_ptr[0] ;
 wire \u_s0.u_sync_wbb.u_resp_if.wr_ptr[1] ;
 wire \u_s0.u_sync_wbb.u_resp_if.wr_ptr[2] ;
 wire \u_s0.u_sync_wbb.wbm_ack_o ;
 wire \u_s0.u_sync_wbb.wbm_lack_o ;
 wire \u_s0.u_sync_wbb.wbs_ack_f ;
 wire \u_s0.u_sync_wbb.wbs_burst ;
 wire \u_s0.u_sync_wbb.wbs_stb_l ;
 wire \u_s1.gnt[0] ;
 wire \u_s1.gnt[1] ;
 wire \u_s1.u_sync_wbb.m_bl_cnt[0] ;
 wire \u_s1.u_sync_wbb.m_bl_cnt[1] ;
 wire \u_s1.u_sync_wbb.m_bl_cnt[2] ;
 wire \u_s1.u_sync_wbb.m_bl_cnt[3] ;
 wire \u_s1.u_sync_wbb.m_bl_cnt[4] ;
 wire \u_s1.u_sync_wbb.m_bl_cnt[5] ;
 wire \u_s1.u_sync_wbb.m_bl_cnt[6] ;
 wire \u_s1.u_sync_wbb.m_bl_cnt[7] ;
 wire \u_s1.u_sync_wbb.m_bl_cnt[8] ;
 wire \u_s1.u_sync_wbb.m_bl_cnt[9] ;
 wire \u_s1.u_sync_wbb.m_cmd_wr_en ;
 wire \u_s1.u_sync_wbb.m_resp_rd_en ;
 wire \u_s1.u_sync_wbb.m_state[0] ;
 wire \u_s1.u_sync_wbb.m_state[1] ;
 wire \u_s1.u_sync_wbb.m_state[2] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[14] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[15] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[16] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[17] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[18] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[19] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[1] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[20] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[21] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[22] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[23] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[24] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[25] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[26] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[27] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[28] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[29] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[2] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[30] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[31] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[32] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[33] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[34] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[35] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[36] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[37] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[38] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[39] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[3] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[40] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[41] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[42] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[43] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[44] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[45] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[46] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[47] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[48] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[49] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[4] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[50] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[53] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[54] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[55] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[56] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[57] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[58] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[59] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[5] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[6] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[7] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[8] ;
 wire \u_s1.u_sync_wbb.s_cmd_rd_data_l[9] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][14] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][15] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][16] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][17] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][18] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][19] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][1] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][20] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][21] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][22] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][23] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][24] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][25] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][26] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][27] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][28] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][29] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][2] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][30] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][31] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][32] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][33] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][34] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][35] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][36] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][37] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][38] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][39] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][3] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][40] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][41] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][42] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][43] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][44] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][45] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][46] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][47] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][48] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][49] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][4] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][50] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][53] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][54] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][55] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][56] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][57] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][58] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][59] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][5] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][6] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][7] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][8] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[0][9] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][14] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][15] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][16] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][17] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][18] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][19] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][1] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][20] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][21] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][22] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][23] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][24] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][25] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][26] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][27] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][28] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][29] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][2] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][30] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][31] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][32] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][33] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][34] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][35] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][36] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][37] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][38] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][39] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][3] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][40] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][41] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][42] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][43] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][44] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][45] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][46] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][47] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][48] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][49] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][4] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][50] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][53] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][54] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][55] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][56] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][57] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][58] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][59] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][5] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][6] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][7] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][8] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[1][9] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][14] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][15] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][16] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][17] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][18] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][19] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][1] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][20] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][21] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][22] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][23] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][24] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][25] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][26] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][27] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][28] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][29] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][2] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][30] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][31] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][32] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][33] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][34] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][35] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][36] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][37] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][38] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][39] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][3] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][40] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][41] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][42] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][43] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][44] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][45] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][46] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][47] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][48] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][49] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][4] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][50] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][53] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][54] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][55] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][56] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][57] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][58] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][59] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][5] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][6] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][7] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][8] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[2][9] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][14] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][15] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][16] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][17] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][18] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][19] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][1] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][20] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][21] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][22] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][23] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][24] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][25] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][26] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][27] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][28] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][29] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][2] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][30] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][31] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][32] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][33] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][34] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][35] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][36] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][37] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][38] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][39] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][3] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][40] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][41] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][42] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][43] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][44] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][45] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][46] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][47] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][48] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][49] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][4] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][50] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][53] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][54] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][55] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][56] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][57] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][58] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][59] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][5] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][6] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][7] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][8] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.mem[3][9] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.rd_ptr[0] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.rd_ptr[1] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.rd_ptr[2] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.wr_ptr[0] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.wr_ptr[1] ;
 wire \u_s1.u_sync_wbb.u_cmd_if.wr_ptr[2] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][0] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][10] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][11] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][12] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][13] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][14] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][15] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][16] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][17] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][18] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][19] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][1] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][20] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][21] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][22] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][23] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][24] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][25] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][26] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][27] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][28] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][29] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][2] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][30] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][31] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][3] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][4] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][5] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][6] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][7] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][8] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[0][9] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][0] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][10] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][11] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][12] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][13] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][14] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][15] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][16] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][17] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][18] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][19] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][1] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][20] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][21] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][22] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][23] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][24] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][25] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][26] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][27] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][28] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][29] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][2] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][30] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][31] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][3] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][4] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][5] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][6] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][7] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][8] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[1][9] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][0] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][10] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][11] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][12] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][13] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][14] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][15] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][16] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][17] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][18] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][19] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][1] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][20] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][21] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][22] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][23] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][24] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][25] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][26] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][27] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][28] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][29] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][2] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][30] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][31] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][3] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][4] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][5] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][6] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][7] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][8] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[2][9] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][0] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][10] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][11] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][12] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][13] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][14] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][15] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][16] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][17] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][18] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][19] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][1] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][20] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][21] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][22] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][23] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][24] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][25] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][26] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][27] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][28] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][29] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][2] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][30] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][31] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][3] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][4] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][5] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][6] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][7] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][8] ;
 wire \u_s1.u_sync_wbb.u_resp_if.mem[3][9] ;
 wire \u_s1.u_sync_wbb.u_resp_if.rd_ptr[0] ;
 wire \u_s1.u_sync_wbb.u_resp_if.rd_ptr[1] ;
 wire \u_s1.u_sync_wbb.u_resp_if.rd_ptr[2] ;
 wire \u_s1.u_sync_wbb.u_resp_if.wr_ptr[0] ;
 wire \u_s1.u_sync_wbb.u_resp_if.wr_ptr[1] ;
 wire \u_s1.u_sync_wbb.u_resp_if.wr_ptr[2] ;
 wire \u_s1.u_sync_wbb.wbm_ack_o ;
 wire \u_s1.u_sync_wbb.wbm_lack_o ;
 wire \u_s1.u_sync_wbb.wbs_ack_f ;
 wire \u_s1.u_sync_wbb.wbs_burst ;
 wire \u_s1.u_sync_wbb.wbs_stb_l ;
 wire \u_s2.gnt[0] ;
 wire \u_s2.gnt[1] ;
 wire \u_s2.u_sync_wbb.m_bl_cnt[0] ;
 wire \u_s2.u_sync_wbb.m_bl_cnt[1] ;
 wire \u_s2.u_sync_wbb.m_bl_cnt[2] ;
 wire \u_s2.u_sync_wbb.m_bl_cnt[3] ;
 wire \u_s2.u_sync_wbb.m_bl_cnt[4] ;
 wire \u_s2.u_sync_wbb.m_bl_cnt[5] ;
 wire \u_s2.u_sync_wbb.m_bl_cnt[6] ;
 wire \u_s2.u_sync_wbb.m_bl_cnt[7] ;
 wire \u_s2.u_sync_wbb.m_bl_cnt[8] ;
 wire \u_s2.u_sync_wbb.m_bl_cnt[9] ;
 wire \u_s2.u_sync_wbb.m_cmd_wr_en ;
 wire \u_s2.u_sync_wbb.m_resp_rd_en ;
 wire \u_s2.u_sync_wbb.m_state[0] ;
 wire \u_s2.u_sync_wbb.m_state[1] ;
 wire \u_s2.u_sync_wbb.m_state[2] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[14] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[15] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[16] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[17] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[18] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[19] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[1] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[20] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[21] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[22] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[23] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[24] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[25] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[26] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[27] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[28] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[29] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[2] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[30] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[31] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[32] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[33] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[34] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[35] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[36] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[37] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[38] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[39] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[3] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[40] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[41] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[42] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[43] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[44] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[45] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[46] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[47] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[48] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[49] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[4] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[50] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[53] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[54] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[55] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[56] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[57] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[58] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[59] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[5] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[60] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[61] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[6] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[7] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[8] ;
 wire \u_s2.u_sync_wbb.s_cmd_rd_data_l[9] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][14] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][15] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][16] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][17] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][18] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][19] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][1] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][20] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][21] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][22] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][23] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][24] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][25] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][26] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][27] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][28] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][29] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][2] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][30] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][31] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][32] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][33] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][34] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][35] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][36] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][37] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][38] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][39] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][3] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][40] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][41] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][42] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][43] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][44] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][45] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][46] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][47] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][48] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][49] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][4] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][50] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][53] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][54] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][55] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][56] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][57] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][58] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][59] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][5] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][60] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][61] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][6] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][7] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][8] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[0][9] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][14] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][15] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][16] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][17] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][18] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][19] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][1] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][20] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][21] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][22] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][23] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][24] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][25] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][26] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][27] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][28] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][29] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][2] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][30] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][31] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][32] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][33] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][34] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][35] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][36] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][37] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][38] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][39] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][3] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][40] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][41] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][42] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][43] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][44] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][45] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][46] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][47] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][48] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][49] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][4] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][50] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][53] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][54] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][55] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][56] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][57] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][58] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][59] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][5] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][60] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][61] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][6] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][7] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][8] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[1][9] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][14] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][15] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][16] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][17] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][18] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][19] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][1] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][20] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][21] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][22] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][23] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][24] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][25] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][26] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][27] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][28] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][29] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][2] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][30] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][31] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][32] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][33] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][34] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][35] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][36] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][37] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][38] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][39] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][3] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][40] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][41] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][42] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][43] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][44] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][45] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][46] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][47] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][48] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][49] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][4] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][50] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][53] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][54] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][55] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][56] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][57] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][58] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][59] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][5] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][60] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][61] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][6] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][7] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][8] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[2][9] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][14] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][15] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][16] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][17] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][18] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][19] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][1] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][20] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][21] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][22] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][23] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][24] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][25] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][26] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][27] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][28] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][29] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][2] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][30] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][31] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][32] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][33] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][34] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][35] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][36] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][37] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][38] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][39] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][3] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][40] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][41] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][42] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][43] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][44] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][45] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][46] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][47] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][48] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][49] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][4] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][50] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][53] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][54] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][55] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][56] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][57] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][58] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][59] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][5] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][60] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][61] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][6] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][7] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][8] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.mem[3][9] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.rd_ptr[0] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.rd_ptr[1] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.rd_ptr[2] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.wr_ptr[0] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.wr_ptr[1] ;
 wire \u_s2.u_sync_wbb.u_cmd_if.wr_ptr[2] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][0] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][10] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][11] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][12] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][13] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][14] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][15] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][16] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][17] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][18] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][19] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][1] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][20] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][21] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][22] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][23] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][24] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][25] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][26] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][27] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][28] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][29] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][2] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][30] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][31] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][3] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][4] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][5] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][6] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][7] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][8] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[0][9] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][0] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][10] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][11] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][12] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][13] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][14] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][15] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][16] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][17] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][18] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][19] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][1] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][20] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][21] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][22] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][23] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][24] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][25] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][26] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][27] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][28] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][29] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][2] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][30] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][31] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][3] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][4] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][5] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][6] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][7] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][8] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[1][9] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][0] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][10] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][11] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][12] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][13] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][14] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][15] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][16] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][17] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][18] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][19] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][1] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][20] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][21] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][22] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][23] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][24] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][25] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][26] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][27] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][28] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][29] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][2] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][30] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][31] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][3] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][4] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][5] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][6] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][7] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][8] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[2][9] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][0] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][10] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][11] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][12] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][13] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][14] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][15] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][16] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][17] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][18] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][19] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][1] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][20] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][21] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][22] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][23] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][24] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][25] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][26] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][27] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][28] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][29] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][2] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][30] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][31] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][3] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][4] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][5] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][6] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][7] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][8] ;
 wire \u_s2.u_sync_wbb.u_resp_if.mem[3][9] ;
 wire \u_s2.u_sync_wbb.u_resp_if.rd_ptr[0] ;
 wire \u_s2.u_sync_wbb.u_resp_if.rd_ptr[1] ;
 wire \u_s2.u_sync_wbb.u_resp_if.rd_ptr[2] ;
 wire \u_s2.u_sync_wbb.u_resp_if.wr_ptr[0] ;
 wire \u_s2.u_sync_wbb.u_resp_if.wr_ptr[1] ;
 wire \u_s2.u_sync_wbb.u_resp_if.wr_ptr[2] ;
 wire \u_s2.u_sync_wbb.wbm_ack_o ;
 wire \u_s2.u_sync_wbb.wbm_lack_o ;
 wire \u_s2.u_sync_wbb.wbs_ack_f ;
 wire \u_s2.u_sync_wbb.wbs_burst ;
 wire \u_s2.u_sync_wbb.wbs_stb_l ;
 wire \u_skew_wi.clk_d1 ;
 wire \u_skew_wi.clk_d10 ;
 wire \u_skew_wi.clk_d11 ;
 wire \u_skew_wi.clk_d12 ;
 wire \u_skew_wi.clk_d13 ;
 wire \u_skew_wi.clk_d14 ;
 wire \u_skew_wi.clk_d15 ;
 wire \u_skew_wi.clk_d2 ;
 wire \u_skew_wi.clk_d3 ;
 wire \u_skew_wi.clk_d4 ;
 wire \u_skew_wi.clk_d5 ;
 wire \u_skew_wi.clk_d6 ;
 wire \u_skew_wi.clk_d7 ;
 wire \u_skew_wi.clk_d8 ;
 wire \u_skew_wi.clk_d9 ;
 wire \u_skew_wi.clk_inbuf ;
 wire \u_skew_wi.clkbuf_1.X1 ;
 wire \u_skew_wi.clkbuf_1.X2 ;
 wire \u_skew_wi.clkbuf_1.X3 ;
 wire \u_skew_wi.clkbuf_10.X1 ;
 wire \u_skew_wi.clkbuf_10.X2 ;
 wire \u_skew_wi.clkbuf_10.X3 ;
 wire \u_skew_wi.clkbuf_11.X1 ;
 wire \u_skew_wi.clkbuf_11.X2 ;
 wire \u_skew_wi.clkbuf_11.X3 ;
 wire \u_skew_wi.clkbuf_12.X1 ;
 wire \u_skew_wi.clkbuf_12.X2 ;
 wire \u_skew_wi.clkbuf_12.X3 ;
 wire \u_skew_wi.clkbuf_13.X1 ;
 wire \u_skew_wi.clkbuf_13.X2 ;
 wire \u_skew_wi.clkbuf_13.X3 ;
 wire \u_skew_wi.clkbuf_14.X1 ;
 wire \u_skew_wi.clkbuf_14.X2 ;
 wire \u_skew_wi.clkbuf_14.X3 ;
 wire \u_skew_wi.clkbuf_15.X1 ;
 wire \u_skew_wi.clkbuf_15.X2 ;
 wire \u_skew_wi.clkbuf_15.X3 ;
 wire \u_skew_wi.clkbuf_2.X1 ;
 wire \u_skew_wi.clkbuf_2.X2 ;
 wire \u_skew_wi.clkbuf_2.X3 ;
 wire \u_skew_wi.clkbuf_3.X1 ;
 wire \u_skew_wi.clkbuf_3.X2 ;
 wire \u_skew_wi.clkbuf_3.X3 ;
 wire \u_skew_wi.clkbuf_4.X1 ;
 wire \u_skew_wi.clkbuf_4.X2 ;
 wire \u_skew_wi.clkbuf_4.X3 ;
 wire \u_skew_wi.clkbuf_5.X1 ;
 wire \u_skew_wi.clkbuf_5.X2 ;
 wire \u_skew_wi.clkbuf_5.X3 ;
 wire \u_skew_wi.clkbuf_6.X1 ;
 wire \u_skew_wi.clkbuf_6.X2 ;
 wire \u_skew_wi.clkbuf_6.X3 ;
 wire \u_skew_wi.clkbuf_7.X1 ;
 wire \u_skew_wi.clkbuf_7.X2 ;
 wire \u_skew_wi.clkbuf_7.X3 ;
 wire \u_skew_wi.clkbuf_8.X1 ;
 wire \u_skew_wi.clkbuf_8.X2 ;
 wire \u_skew_wi.clkbuf_8.X3 ;
 wire \u_skew_wi.clkbuf_9.X1 ;
 wire \u_skew_wi.clkbuf_9.X2 ;
 wire \u_skew_wi.clkbuf_9.X3 ;
 wire \u_skew_wi.d00 ;
 wire \u_skew_wi.d01 ;
 wire \u_skew_wi.d02 ;
 wire \u_skew_wi.d03 ;
 wire \u_skew_wi.d04 ;
 wire \u_skew_wi.d05 ;
 wire \u_skew_wi.d06 ;
 wire \u_skew_wi.d07 ;
 wire \u_skew_wi.d10 ;
 wire \u_skew_wi.d11 ;
 wire \u_skew_wi.d12 ;
 wire \u_skew_wi.d13 ;
 wire \u_skew_wi.d20 ;
 wire \u_skew_wi.d21 ;
 wire \u_skew_wi.d30 ;
 wire \u_skew_wi.in0 ;
 wire \u_skew_wi.in1 ;
 wire \u_skew_wi.in10 ;
 wire \u_skew_wi.in11 ;
 wire \u_skew_wi.in12 ;
 wire \u_skew_wi.in13 ;
 wire \u_skew_wi.in14 ;
 wire \u_skew_wi.in15 ;
 wire \u_skew_wi.in2 ;
 wire \u_skew_wi.in3 ;
 wire \u_skew_wi.in4 ;
 wire \u_skew_wi.in5 ;
 wire \u_skew_wi.in6 ;
 wire \u_skew_wi.in7 ;
 wire \u_skew_wi.in8 ;
 wire \u_skew_wi.in9 ;
 wire \u_wbi_arb.gnt[0] ;
 wire \u_wbi_arb.gnt[1] ;

 sky130_fd_sc_hd__diode_2 ANTENNA__3614__A (.DIODE(m2_wbd_bl_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__A (.DIODE(net1404));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__A (.DIODE(net1405));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__A (.DIODE(net1409));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__A (.DIODE(net1408));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__A (.DIODE(m2_wbd_bry_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3622__A (.DIODE(\u_s2.u_sync_wbb.m_bl_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3625__A (.DIODE(net1396));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__A (.DIODE(m0_wbd_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__A (.DIODE(m0_wbd_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__A (.DIODE(m0_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__A (.DIODE(m3_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__A (.DIODE(m2_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__A (.DIODE(m1_wbd_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__A (.DIODE(m1_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A (.DIODE(\u_s1.u_sync_wbb.m_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__A (.DIODE(\u_s1.u_sync_wbb.wbm_lack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__A (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__A (.DIODE(s0_wbd_lack_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__A (.DIODE(net1276));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__A (.DIODE(net1274));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__A (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__A_N (.DIODE(net1328));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__B (.DIODE(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__A (.DIODE(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__B (.DIODE(net1328));
 sky130_fd_sc_hd__diode_2 ANTENNA__3657__A_N (.DIODE(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3657__B (.DIODE(net1338));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__A (.DIODE(net1338));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__B (.DIODE(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__B (.DIODE(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__A2 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__A (.DIODE(_1719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__A (.DIODE(\u_s0.u_sync_wbb.m_cmd_wr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__B (.DIODE(net1254));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__A (.DIODE(net1264));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__A_N (.DIODE(net1371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__B (.DIODE(net1375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__C (.DIODE(net1563));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__A (.DIODE(net1371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__B (.DIODE(net1375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__C (.DIODE(m3_wbd_bry_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A (.DIODE(net1371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__B (.DIODE(net1375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__A_N (.DIODE(\u_s0.gnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__B (.DIODE(net1371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__A (.DIODE(net1193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__A1 (.DIODE(net1259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__A2 (.DIODE(m2_wbd_bry_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__D1 (.DIODE(net1205));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__B1_N (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__A (.DIODE(m3_wbd_adr_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__B (.DIODE(m3_wbd_adr_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__C (.DIODE(m3_wbd_adr_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__D (.DIODE(m3_wbd_adr_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__A (.DIODE(m3_wbd_adr_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__B (.DIODE(m3_wbd_adr_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__C (.DIODE(m3_wbd_adr_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__D_N (.DIODE(m3_wbd_adr_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__A (.DIODE(m3_wbd_adr_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__B (.DIODE(m3_wbd_adr_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__C (.DIODE(m3_wbd_adr_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__D (.DIODE(m3_wbd_adr_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__A (.DIODE(m3_wbd_adr_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__B (.DIODE(m3_wbd_adr_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__A (.DIODE(m3_wbd_adr_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__B (.DIODE(m3_wbd_adr_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__C_N (.DIODE(m3_wbd_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__A (.DIODE(m3_wbd_adr_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__B (.DIODE(m3_wbd_adr_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__C_N (.DIODE(m3_wbd_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__A (.DIODE(net1208));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__B (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__C (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__A (.DIODE(m0_wbd_adr_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__B (.DIODE(m0_wbd_adr_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__A (.DIODE(m0_wbd_adr_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__B (.DIODE(m0_wbd_adr_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__C (.DIODE(m0_wbd_adr_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__D_N (.DIODE(m0_wbd_adr_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__A (.DIODE(m0_wbd_adr_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__B (.DIODE(m0_wbd_adr_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__C (.DIODE(m0_wbd_adr_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__D (.DIODE(m0_wbd_adr_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__A (.DIODE(m0_wbd_adr_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__B (.DIODE(m0_wbd_adr_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__C (.DIODE(m0_wbd_adr_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__D (.DIODE(m0_wbd_adr_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__B (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__C (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__D (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__B (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__C (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__B (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__C (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__D (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__B (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__A (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__A (.DIODE(m0_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__A1 (.DIODE(m0_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__A2 (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__B2 (.DIODE(m3_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__A (.DIODE(m1_wbd_adr_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__B (.DIODE(m1_wbd_adr_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__C_N (.DIODE(m1_wbd_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3705__A (.DIODE(m1_wbd_adr_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3705__B (.DIODE(m1_wbd_adr_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3705__C (.DIODE(m1_wbd_adr_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3705__D_N (.DIODE(m1_wbd_adr_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__A (.DIODE(m1_wbd_adr_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__B (.DIODE(m1_wbd_adr_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__C (.DIODE(m1_wbd_adr_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__D (.DIODE(m1_wbd_adr_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__A (.DIODE(m1_wbd_adr_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__B (.DIODE(m1_wbd_adr_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__C (.DIODE(m1_wbd_adr_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__D (.DIODE(m1_wbd_adr_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__A (.DIODE(m1_wbd_adr_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__B (.DIODE(m1_wbd_adr_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__C_N (.DIODE(m1_wbd_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__A (.DIODE(m2_wbd_adr_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__B (.DIODE(m2_wbd_adr_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__C (.DIODE(m2_wbd_adr_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__D (.DIODE(m2_wbd_adr_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__A (.DIODE(m2_wbd_adr_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__B (.DIODE(m2_wbd_adr_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__C (.DIODE(m2_wbd_adr_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__D_N (.DIODE(m2_wbd_adr_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__A (.DIODE(m2_wbd_adr_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__B (.DIODE(m2_wbd_adr_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__C (.DIODE(m2_wbd_adr_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__D (.DIODE(m2_wbd_adr_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__A (.DIODE(m2_wbd_adr_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__B (.DIODE(m2_wbd_adr_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__A (.DIODE(m2_wbd_adr_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__B (.DIODE(m2_wbd_adr_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__C_N (.DIODE(m2_wbd_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__A (.DIODE(m2_wbd_adr_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__B (.DIODE(m2_wbd_adr_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__C_N (.DIODE(m2_wbd_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__A (.DIODE(net1193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__A (.DIODE(m2_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__A1 (.DIODE(m1_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__B1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__B2 (.DIODE(m2_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__A1 (.DIODE(_1759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__A2 (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__B1 (.DIODE(\u_s0.u_sync_wbb.wbm_lack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__A1 (.DIODE(_1759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__A2 (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__B1 (.DIODE(\u_s0.u_sync_wbb.wbm_lack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__C1 (.DIODE(_1735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__A1 (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__A2 (.DIODE(m2_wbd_bl_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__B2 (.DIODE(m3_wbd_bl_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__C1 (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__A1 (.DIODE(net1564));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__A2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__A1 (.DIODE(m3_wbd_bl_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__B1 (.DIODE(net1193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__B2 (.DIODE(m2_wbd_bl_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__A1 (.DIODE(m3_wbd_bl_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__B1 (.DIODE(net1193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__B2 (.DIODE(m2_wbd_bl_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__A1 (.DIODE(m1_wbd_bl_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__A2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__B1 (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__A (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__B (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__C_N (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__A1 (.DIODE(m3_wbd_bl_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__B1 (.DIODE(net1193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__B2 (.DIODE(m2_wbd_bl_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__A1 (.DIODE(m1_wbd_bl_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__A2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__A1 (.DIODE(m3_wbd_bl_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__B1 (.DIODE(net1193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__B2 (.DIODE(m2_wbd_bl_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__A1 (.DIODE(m3_wbd_bl_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__B1 (.DIODE(net1193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__B2 (.DIODE(m2_wbd_bl_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__A (.DIODE(_1792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__B (.DIODE(_1794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__A1 (.DIODE(m3_wbd_bl_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__B1 (.DIODE(net1193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__B2 (.DIODE(m2_wbd_bl_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__A1 (.DIODE(m3_wbd_bl_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__B1 (.DIODE(net1193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__B2 (.DIODE(m2_wbd_bl_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__A (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__B (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__A1 (.DIODE(m3_wbd_bl_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__B1 (.DIODE(net1193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__B2 (.DIODE(m2_wbd_bl_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A1 (.DIODE(m3_wbd_bl_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A2 (.DIODE(net1209));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__B1 (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__B2 (.DIODE(m2_wbd_bl_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__B (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__C (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__B (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__D (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3748__A (.DIODE(net1271));
 sky130_fd_sc_hd__diode_2 ANTENNA__3748__B (.DIODE(net1375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3748__C (.DIODE(m1_wbd_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__A1 (.DIODE(net1259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__A2 (.DIODE(m2_wbd_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__B1 (.DIODE(net1208));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__B2 (.DIODE(m3_wbd_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__C1 (.DIODE(net1204));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__A1 (.DIODE(m0_wbd_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__A2 (.DIODE(net1199));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__A (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__A_N (.DIODE(\u_s0.u_sync_wbb.wbm_lack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__C (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__B (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A_N (.DIODE(net1315));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__A_N (.DIODE(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__B (.DIODE(net1320));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__B (.DIODE(net1315));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__B (.DIODE(_1814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__A (.DIODE(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__B (.DIODE(net1321));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__A (.DIODE(\u_s0.u_sync_wbb.wbm_ack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3764__A1 (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3764__A2 (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3764__B1 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__A1 (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__A2 (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__B1 (.DIODE(\u_s0.u_sync_wbb.m_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__C1 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__B (.DIODE(_1735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__B (.DIODE(\u_s0.u_sync_wbb.m_bl_cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__C (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__C (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__B (.DIODE(\u_s0.u_sync_wbb.m_bl_cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3773__C (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__A2 (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__B1 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A (.DIODE(net1404));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__B (.DIODE(net1405));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__A (.DIODE(net1404));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__B (.DIODE(net1405));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__A (.DIODE(net1404));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__B (.DIODE(net1405));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__A_N (.DIODE(\u_s1.gnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__A (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__B (.DIODE(net1405));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__A (.DIODE(m1_wbd_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__B (.DIODE(net1183));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__A1 (.DIODE(net1240));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__A2 (.DIODE(m2_wbd_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__B1 (.DIODE(net1185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__B2 (.DIODE(m3_wbd_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__C1 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__A1 (.DIODE(m0_wbd_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__A2 (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__A_N (.DIODE(net1358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__B (.DIODE(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A (.DIODE(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__B (.DIODE(net1365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__A (.DIODE(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__B (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__A_N (.DIODE(net1365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A1 (.DIODE(net1404));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__A1 (.DIODE(net1252));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__A2 (.DIODE(net1563));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__B1 (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__B2 (.DIODE(m3_wbd_bry_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__A (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__B (.DIODE(_1849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__A_N (.DIODE(net1405));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__B (.DIODE(net1404));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__A (.DIODE(m2_wbd_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__C_N (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A (.DIODE(m3_wbd_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__B (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__A (.DIODE(m3_wbd_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__C (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__D_N (.DIODE(net1185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__C (.DIODE(m0_wbd_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__D (.DIODE(_1830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__A1 (.DIODE(m3_wbd_bl_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__A2 (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__B1 (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__B2 (.DIODE(m2_wbd_bl_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__A (.DIODE(net1404));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__C (.DIODE(m3_wbd_bl_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A1 (.DIODE(m1_wbd_bl_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A2 (.DIODE(net1183));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__B1 (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__B2 (.DIODE(m2_wbd_bl_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__A1 (.DIODE(m3_wbd_bl_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__A2 (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__B1 (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__B2 (.DIODE(m2_wbd_bl_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__A (.DIODE(_1860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__A (.DIODE(net1404));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__B (.DIODE(net1405));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__C (.DIODE(m3_wbd_bl_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__A1 (.DIODE(m1_wbd_bl_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__A2 (.DIODE(net1184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__B1 (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__B2 (.DIODE(m2_wbd_bl_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__A (.DIODE(_1856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__B (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__C (.DIODE(_1860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__D (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__A1 (.DIODE(m3_wbd_bl_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__A2 (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__B1 (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__B2 (.DIODE(m2_wbd_bl_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__A1 (.DIODE(m3_wbd_bl_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__A2 (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__B1 (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__B2 (.DIODE(m2_wbd_bl_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A1 (.DIODE(m3_wbd_bl_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A2 (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__B1 (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__B2 (.DIODE(m2_wbd_bl_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__A1 (.DIODE(m3_wbd_bl_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__A2 (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__B1 (.DIODE(_1851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__B2 (.DIODE(m2_wbd_bl_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__A (.DIODE(_1867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__B (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__C (.DIODE(_1869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__A (.DIODE(_1866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__A (.DIODE(_1866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A1 (.DIODE(m3_wbd_bl_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A2 (.DIODE(_1832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__B1 (.DIODE(_1851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__B2 (.DIODE(m2_wbd_bl_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__A2 (.DIODE(\u_s1.gnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A1 (.DIODE(net1564));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A2 (.DIODE(net1252));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__B1 (.DIODE(_1832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__B2 (.DIODE(m3_wbd_bl_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__B (.DIODE(_1872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__C (.DIODE(_1873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__D_N (.DIODE(_1875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__A (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__B (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__C (.DIODE(_1849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__A (.DIODE(m0_wbd_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__C (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__A (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__C (.DIODE(_1834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__A (.DIODE(m2_wbd_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__D_N (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A1 (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A2 (.DIODE(_1878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__B1 (.DIODE(_1880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__B (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__B (.DIODE(net1345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__B (.DIODE(net1344));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__A2 (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__B1 (.DIODE(\u_s1.u_sync_wbb.wbm_ack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__A2 (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__A1 (.DIODE(\u_s1.u_sync_wbb.wbm_ack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__B (.DIODE(\u_s1.u_sync_wbb.u_resp_if.rd_ptr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__A1 (.DIODE(_1888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__A2 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__B1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__B (.DIODE(_1892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__B (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__C (.DIODE(_1849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__A (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__D (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__D_N (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__B (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__C (.DIODE(_1896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A (.DIODE(\u_s1.u_sync_wbb.m_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__D_N (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__A (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__C (.DIODE(_1896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__A2 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A1 (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A2 (.DIODE(_1902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__B1 (.DIODE(_1903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__C1 (.DIODE(_1900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__S0 (.DIODE(net1339));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__S1 (.DIODE(net1329));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__A1 (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__S (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__S0 (.DIODE(net1341));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__S1 (.DIODE(net1331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__A1 (.DIODE(_1905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__S (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__S0 (.DIODE(net1341));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__S1 (.DIODE(net1331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__A1 (.DIODE(_1906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__S (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__S0 (.DIODE(net1340));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__S1 (.DIODE(net1330));
 sky130_fd_sc_hd__diode_2 ANTENNA__3857__A1 (.DIODE(_1907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3857__S (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__S0 (.DIODE(net1340));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__S1 (.DIODE(net1330));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__A1 (.DIODE(_1908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__S (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__S0 (.DIODE(net1340));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__S1 (.DIODE(net1330));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__A1 (.DIODE(_1909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__S (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__S0 (.DIODE(net1341));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__S1 (.DIODE(net1331));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__A1 (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__S (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__S0 (.DIODE(net1340));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__S1 (.DIODE(net1330));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__A1 (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__S (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__S0 (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__S1 (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__A1 (.DIODE(_1912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__S (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__B (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__A1 (.DIODE(_1735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__A_N (.DIODE(net1410));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__B (.DIODE(net1408));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__A (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__B (.DIODE(net1407));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__A (.DIODE(net1410));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__B (.DIODE(\u_s2.gnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__A1 (.DIODE(m2_wbd_bl_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__A2 (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__B2 (.DIODE(m3_wbd_bl_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__A (.DIODE(m3_wbd_bl_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__B (.DIODE(net1410));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__C (.DIODE(net1408));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__A_N (.DIODE(net1407));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__B (.DIODE(net1409));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__A1 (.DIODE(m2_wbd_bl_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__A2 (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__B1 (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__B2 (.DIODE(m1_wbd_bl_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__A1 (.DIODE(m2_wbd_bl_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__A2 (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__B2 (.DIODE(m3_wbd_bl_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__A (.DIODE(m3_wbd_bl_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__B (.DIODE(net1410));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__C (.DIODE(net1408));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__A1 (.DIODE(m2_wbd_bl_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__A2 (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__B1 (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__B2 (.DIODE(m1_wbd_bl_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__A (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__B (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__C (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__D (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__A1 (.DIODE(m2_wbd_bl_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__A2 (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__B2 (.DIODE(m3_wbd_bl_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__A1 (.DIODE(m2_wbd_bl_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__A2 (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__B2 (.DIODE(m3_wbd_bl_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__A1 (.DIODE(m2_wbd_bl_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__A2 (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__B2 (.DIODE(m3_wbd_bl_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A1 (.DIODE(m2_wbd_bl_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A2 (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__B2 (.DIODE(m3_wbd_bl_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__A1 (.DIODE(m2_wbd_bl_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__A2 (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__B1 (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__B2 (.DIODE(m3_wbd_bl_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__B (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__C (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__A1 (.DIODE(m2_wbd_bl_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__B2 (.DIODE(m3_wbd_bl_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__A (.DIODE(net1409));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__B (.DIODE(net1407));
 sky130_fd_sc_hd__diode_2 ANTENNA__3892__A (.DIODE(net1409));
 sky130_fd_sc_hd__diode_2 ANTENNA__3892__B (.DIODE(net1407));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__A2 (.DIODE(\u_s2.gnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__B1 (.DIODE(\u_s2.gnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__A1 (.DIODE(net1564));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__A2 (.DIODE(net1225));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__B2 (.DIODE(m3_wbd_bl_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__A1 (.DIODE(net1564));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__A2 (.DIODE(net1225));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__B2 (.DIODE(m3_wbd_bl_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__B (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__B (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__A (.DIODE(net1410));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__B (.DIODE(net1408));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__C (.DIODE(m3_wbd_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__A1 (.DIODE(net1233));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__A2 (.DIODE(m2_wbd_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__B1 (.DIODE(m1_wbd_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__B2 (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__C1 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__A1 (.DIODE(m0_wbd_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__A2 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__A_N (.DIODE(net1389));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__A (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__B (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.rd_ptr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__B (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__B (.DIODE(net1389));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A1 (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__A (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__C1 (.DIODE(\u_s2.u_sync_wbb.m_cmd_wr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__A1 (.DIODE(m3_wbd_bry_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__B1 (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__B2 (.DIODE(net1563));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__A1 (.DIODE(\u_s2.gnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__B1 (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__A1 (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__B1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__A (.DIODE(m1_wbd_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__C_N (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__A (.DIODE(m1_wbd_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__B (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__D_N (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__A (.DIODE(m3_wbd_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__B (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__A (.DIODE(m3_wbd_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__C (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__D_N (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__A (.DIODE(m2_wbd_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__A (.DIODE(m2_wbd_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__B (.DIODE(m0_wbd_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__C (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__A1 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__A2 (.DIODE(_1962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__D1 (.DIODE(_1957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__A (.DIODE(m3_wbd_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3921__A (.DIODE(m2_wbd_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3921__D_N (.DIODE(m2_wbd_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__A (.DIODE(m3_wbd_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__C_N (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__D_N (.DIODE(m3_wbd_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__B (.DIODE(m0_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__A_N (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__C (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__A1 (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__A2 (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__B1 (.DIODE(_1969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__A1 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__A2 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__B1 (.DIODE(net1400));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__C1 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__A1 (.DIODE(net1400));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__A2 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__A3 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__A_N (.DIODE(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__B (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__A (.DIODE(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__B (.DIODE(net1379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__A1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__A2 (.DIODE(net1383));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__B1 (.DIODE(\u_s2.u_sync_wbb.wbm_ack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__B2 (.DIODE(_1974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__A1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__A2 (.DIODE(net1383));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__B1 (.DIODE(_1974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__A1 (.DIODE(\u_s2.u_sync_wbb.wbm_ack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__A3 (.DIODE(_1980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__B1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__B (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__B (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__A (.DIODE(_1982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__B (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A (.DIODE(\u_s2.u_sync_wbb.m_bl_cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__B (.DIODE(\u_s2.u_sync_wbb.m_bl_cnt[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__C (.DIODE(\u_s2.u_sync_wbb.m_bl_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__B (.DIODE(\u_s2.u_sync_wbb.m_bl_cnt[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__C (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__A (.DIODE(_1987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__A (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__B (.DIODE(_1971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__B1 (.DIODE(_1987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__A1 (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__A2 (.DIODE(_1987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__A1 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__A2 (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__B1 (.DIODE(net1400));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__C1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__D1 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A1 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A2 (.DIODE(_1987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__C (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__D (.DIODE(_1971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__A (.DIODE(\u_s1.u_sync_wbb.m_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__A2 (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__C1 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__D1 (.DIODE(\u_s0.u_sync_wbb.wbm_lack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A1 (.DIODE(_1759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A2 (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__B1 (.DIODE(_1997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__B2 (.DIODE(\u_s0.u_sync_wbb.m_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__A1 (.DIODE(_1892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__A2 (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__B1 (.DIODE(\u_s1.u_sync_wbb.m_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__A_N (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__B (.DIODE(_1849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__C (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__D (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__A (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__B (.DIODE(net1492));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__A (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__A2 (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.mem[2][50] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__A3 (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.mem[3][50] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__S0 (.DIODE(net1396));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__S1 (.DIODE(net1389));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__S (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__S0 (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__S1 (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__A1 (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__S (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__S0 (.DIODE(net1339));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__S1 (.DIODE(net1329));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__A1 (.DIODE(_2007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__S (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__A2 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__A2 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__A2 (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__B1 (.DIODE(net1278));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__A (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__B (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__A (.DIODE(m2_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__B (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__A (.DIODE(net1277));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__B (.DIODE(net1274));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__B (.DIODE(net1277));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__A1 (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__A2 (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__A (.DIODE(net1278));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__B (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__A (.DIODE(net1276));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__B (.DIODE(net1274));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__A (.DIODE(m0_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__B (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__B1 (.DIODE(_2019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__A (.DIODE(\u_reg.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__B (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__A (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__A1 (.DIODE(net1366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__B2 (.DIODE(\u_reg.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__A1 (.DIODE(\u_s0.u_sync_wbb.wbm_lack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__A2 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__B2 (.DIODE(net1401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__A1 (.DIODE(net1367));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__B2 (.DIODE(\u_reg.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__A1 (.DIODE(\u_s0.u_sync_wbb.wbm_ack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__B2 (.DIODE(net1402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__S0 (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__S1 (.DIODE(net1314));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__A1 (.DIODE(net1312));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__B1 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__S0 (.DIODE(net1383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__S1 (.DIODE(net1379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__S0 (.DIODE(net1349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__S1 (.DIODE(net1345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__A2 (.DIODE(net1140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__B1 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__B2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__S0 (.DIODE(net1350));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__S1 (.DIODE(net1346));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__A1 (.DIODE(\u_reg.reg_rdata[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__B1 (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__S0 (.DIODE(net1321));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__S1 (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__S0 (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__S1 (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__A2 (.DIODE(_2036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__B1 (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4015__S0 (.DIODE(net1322));
 sky130_fd_sc_hd__diode_2 ANTENNA__4015__S1 (.DIODE(net1315));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__A1 (.DIODE(\u_reg.reg_rdata[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__B1 (.DIODE(net1134));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__S0 (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__S1 (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__S0 (.DIODE(net1350));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__S1 (.DIODE(net1346));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__A2 (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__B1 (.DIODE(net1129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__S0 (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__S1 (.DIODE(net1344));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__A1 (.DIODE(\u_reg.reg_rdata[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__B1 (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__B2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__S0 (.DIODE(net1321));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__S1 (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__A1 (.DIODE(\u_s2.u_sync_wbb.u_resp_if.mem[1][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__S0 (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__S1 (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4025__A2 (.DIODE(_2046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4025__B1 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__S0 (.DIODE(net1320));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__S1 (.DIODE(net1317));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__A1 (.DIODE(net1311));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__B1 (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__S0 (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__S1 (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__S0 (.DIODE(net1349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__S1 (.DIODE(net1345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__A2 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__B1 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__S0 (.DIODE(net1350));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__S1 (.DIODE(net1346));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__A1 (.DIODE(net1310));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__B1 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__B2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__S0 (.DIODE(net1320));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__S1 (.DIODE(net1317));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__S0 (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__S1 (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__A2 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__B1 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__S0 (.DIODE(net1350));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__S1 (.DIODE(net1346));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__A1 (.DIODE(\u_reg.reg_rdata[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__B1 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__B2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__S0 (.DIODE(net1320));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__S1 (.DIODE(net1315));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__S0 (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__S1 (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__A1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__A2 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__B1 (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__S0 (.DIODE(net1322));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__S1 (.DIODE(net1315));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__A1 (.DIODE(net1309));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__B1 (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__A2 (.DIODE(\u_s2.u_sync_wbb.u_resp_if.mem[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__S0 (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__S1 (.DIODE(net1376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__S0 (.DIODE(net1349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__S1 (.DIODE(net1345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__A2 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__B1 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__B2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__4051__S0 (.DIODE(net1349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4051__S1 (.DIODE(net1346));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__A1 (.DIODE(net1308));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__A2 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__B1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__S0 (.DIODE(net1321));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__S1 (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__S0 (.DIODE(net1383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__S1 (.DIODE(net1379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__A2 (.DIODE(_2071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__B1 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__S0 (.DIODE(net1349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__S1 (.DIODE(net1345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__A1 (.DIODE(net1307));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__B1 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__S0 (.DIODE(net1321));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__S1 (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__S0 (.DIODE(net1383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__S1 (.DIODE(net1379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__A1 (.DIODE(_1780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__A2 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__B1 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__S0 (.DIODE(net1347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__S1 (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__A1 (.DIODE(net1306));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__A2 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__B1 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__S0 (.DIODE(net1321));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__S1 (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__S0 (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__S1 (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__A1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__A2 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__B1 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__S0 (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__S1 (.DIODE(net1314));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__A1 (.DIODE(net1305));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__B1 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__S0 (.DIODE(net1381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__S1 (.DIODE(net1377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__S0 (.DIODE(net1347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__S1 (.DIODE(net1344));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__A1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__A2 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__B1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__B2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__4075__S0 (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA__4075__S1 (.DIODE(net1344));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__A1 (.DIODE(net1304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__A2 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__B1 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__B2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__S0 (.DIODE(net1318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__S1 (.DIODE(net1313));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__S0 (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__S1 (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__A1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__A2 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__B1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__S0 (.DIODE(net1351));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__S1 (.DIODE(net1344));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__A1 (.DIODE(net1302));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__B1 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__B2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__S0 (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__S1 (.DIODE(net1314));
 sky130_fd_sc_hd__diode_2 ANTENNA__4084__S0 (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4084__S1 (.DIODE(net1376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__A1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__A2 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__B1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__S0 (.DIODE(net1349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__S1 (.DIODE(net1345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__A1 (.DIODE(net1300));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__A2 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__B1 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__B2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__4089__S0 (.DIODE(net1318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4089__S1 (.DIODE(net1313));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__S0 (.DIODE(net1381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__S1 (.DIODE(net1377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__A1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__A2 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__B1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__S0 (.DIODE(net1320));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__S1 (.DIODE(net1315));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__A1 (.DIODE(net1298));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__A2 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__B1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__B2 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__S0 (.DIODE(net1383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__S1 (.DIODE(net1379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__S0 (.DIODE(net1349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__S1 (.DIODE(net1345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__A1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__A2 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__B1 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__B2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__S0 (.DIODE(net1349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__S1 (.DIODE(net1345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__A1 (.DIODE(net1296));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__B1 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__B2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__4101__S0 (.DIODE(net1318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4101__S1 (.DIODE(net1313));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__S0 (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__S1 (.DIODE(net1376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4103__A2 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA__4103__B1 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__S0 (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__S1 (.DIODE(net1344));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__A1 (.DIODE(net1295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__A2 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__B1 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__B2 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__S0 (.DIODE(net1320));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__S1 (.DIODE(net1315));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__S0 (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__S1 (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__A1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__A2 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__B1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__S0 (.DIODE(net1322));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__S1 (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__A1 (.DIODE(\u_reg.reg_rdata[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__B1 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__B2 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__4113__S0 (.DIODE(net1383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4113__S1 (.DIODE(net1379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__S0 (.DIODE(net1349));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__S1 (.DIODE(net1345));
 sky130_fd_sc_hd__diode_2 ANTENNA__4115__A2 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA__4115__B1 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__S0 (.DIODE(net1347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__S1 (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__A1 (.DIODE(\u_reg.reg_rdata[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__B1 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__S0 (.DIODE(net1318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__S1 (.DIODE(net1313));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__A2 (.DIODE(\u_s2.u_sync_wbb.u_resp_if.mem[2][19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__S0 (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__S1 (.DIODE(net1376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__A2 (.DIODE(_2126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__B1 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__S0 (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__S1 (.DIODE(net1344));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__A1 (.DIODE(net1293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__A2 (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__B1 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__B2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__S0 (.DIODE(net1318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__S1 (.DIODE(net1313));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__S0 (.DIODE(net1383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__S1 (.DIODE(net1379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__A2 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__B1 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__B2 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__4129__S0 (.DIODE(net1320));
 sky130_fd_sc_hd__diode_2 ANTENNA__4129__S1 (.DIODE(net1315));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__A1 (.DIODE(net1291));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__A2 (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__B1 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__S0 (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__S1 (.DIODE(net1376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4132__S0 (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA__4132__S1 (.DIODE(net1344));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__A1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__A2 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__B1 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__B2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__4135__S0 (.DIODE(net1318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4135__S1 (.DIODE(net1313));
 sky130_fd_sc_hd__diode_2 ANTENNA__4136__A1 (.DIODE(net1290));
 sky130_fd_sc_hd__diode_2 ANTENNA__4136__A2 (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4136__B1 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA__4137__S0 (.DIODE(net1381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4137__S1 (.DIODE(net1377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__S0 (.DIODE(net1347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__S1 (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__A1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__A2 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__B1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__B2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__S0 (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__S1 (.DIODE(net1314));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__A1 (.DIODE(\u_reg.reg_rdata[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__A2 (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__B1 (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__B2 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__4143__S0 (.DIODE(net1383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4143__S1 (.DIODE(net1379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4144__S0 (.DIODE(net1347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4144__S1 (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__4145__A1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__4145__A2 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA__4145__B1 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA__4145__B2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__4147__S0 (.DIODE(net1321));
 sky130_fd_sc_hd__diode_2 ANTENNA__4147__S1 (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA__4148__A1 (.DIODE(net1289));
 sky130_fd_sc_hd__diode_2 ANTENNA__4148__B1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA__4149__S0 (.DIODE(net1381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4149__S1 (.DIODE(net1377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__S0 (.DIODE(net1347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__S1 (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__A2 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__B1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__S0 (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__S1 (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__A1 (.DIODE(net1288));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__B1 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA__4155__S0 (.DIODE(net1321));
 sky130_fd_sc_hd__diode_2 ANTENNA__4155__S1 (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__S0 (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__S1 (.DIODE(net1376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4157__A2 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA__4157__B1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__S0 (.DIODE(net1347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__S1 (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__A1 (.DIODE(net1286));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__A2 (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__B1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__B2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__S0 (.DIODE(net1318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__S1 (.DIODE(net1313));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__A1 (.DIODE(\u_s2.u_sync_wbb.u_resp_if.mem[1][26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__S0 (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__S1 (.DIODE(net1376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4163__A1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__4163__A2 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA__4163__B1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA__4163__B2 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__S0 (.DIODE(net1347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__S1 (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__A1 (.DIODE(net1285));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__A2 (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__B1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__B2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__4167__S0 (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA__4167__S1 (.DIODE(net1314));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__A0 (.DIODE(\u_s2.u_sync_wbb.u_resp_if.mem[0][27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__S0 (.DIODE(net1381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__S1 (.DIODE(net1377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__A2 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__B1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__B2 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__4171__S0 (.DIODE(net1318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4171__S1 (.DIODE(net1313));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__A1 (.DIODE(net1284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__B1 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__B2 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__S0 (.DIODE(net1381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__S1 (.DIODE(net1377));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__S0 (.DIODE(net1347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__S1 (.DIODE(net1344));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__A2 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__B1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA__4177__S0 (.DIODE(net1351));
 sky130_fd_sc_hd__diode_2 ANTENNA__4177__S1 (.DIODE(\u_s1.u_sync_wbb.u_resp_if.rd_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__A1 (.DIODE(net1282));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__A2 (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__B1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__B2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__4179__S0 (.DIODE(net1318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4179__S1 (.DIODE(net1313));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__S0 (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__S1 (.DIODE(net1376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4181__A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA__4181__B1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA__4181__B2 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__4183__S0 (.DIODE(net1347));
 sky130_fd_sc_hd__diode_2 ANTENNA__4183__S1 (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__A1 (.DIODE(net1281));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__B1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA__4185__S0 (.DIODE(net1318));
 sky130_fd_sc_hd__diode_2 ANTENNA__4185__S1 (.DIODE(net1313));
 sky130_fd_sc_hd__diode_2 ANTENNA__4186__S0 (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4186__S1 (.DIODE(net1376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__A1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__A2 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__B1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA__4189__S0 (.DIODE(net1321));
 sky130_fd_sc_hd__diode_2 ANTENNA__4189__S1 (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA__4190__A1 (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA__4190__A2 (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4190__B1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__A0 (.DIODE(\u_s2.u_sync_wbb.u_resp_if.mem[0][31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__S0 (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__S1 (.DIODE(net1376));
 sky130_fd_sc_hd__diode_2 ANTENNA__4192__S0 (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA__4192__S1 (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__4193__A1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__4193__A2 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA__4193__B1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA__4193__B2 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__4195__B (.DIODE(_1833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__A1 (.DIODE(\u_reg.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__A2 (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__B1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__B2 (.DIODE(net1366));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__A1 (.DIODE(\u_s0.u_sync_wbb.wbm_lack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__A2 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__B1 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__B2 (.DIODE(net1401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__A1 (.DIODE(\u_reg.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__A2 (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__B1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__B2 (.DIODE(net1367));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__A1 (.DIODE(\u_s0.u_sync_wbb.wbm_ack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__A2 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__B1 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__B2 (.DIODE(net1402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__A1 (.DIODE(net1312));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__B1 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__A2 (.DIODE(net1140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__B1 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__A1 (.DIODE(\u_reg.reg_rdata[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__A2 (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__B1 (.DIODE(_2036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__B2 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__A1 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__A2 (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__B1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__B2 (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4208__A1 (.DIODE(\u_reg.reg_rdata[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4208__A2 (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4208__B1 (.DIODE(net1129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4208__B2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__A1 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__A2 (.DIODE(net1134));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__B1 (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__B2 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__4211__A1 (.DIODE(\u_reg.reg_rdata[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4211__A2 (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4211__B1 (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4211__B2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__A1 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__A2 (.DIODE(_2046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__B1 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__B2 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__A1 (.DIODE(net1311));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__A2 (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__B1 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__B2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__A2 (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__B1 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA__4217__A1 (.DIODE(net1310));
 sky130_fd_sc_hd__diode_2 ANTENNA__4217__B1 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__A2 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__B1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__B2 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__A1 (.DIODE(\u_reg.reg_rdata[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__B1 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__A2 (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__B2 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4223__A1 (.DIODE(net1309));
 sky130_fd_sc_hd__diode_2 ANTENNA__4223__A2 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4223__B1 (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA__4223__B2 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__A2 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__B1 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__A1 (.DIODE(net1308));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__B1 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__A1 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__A2 (.DIODE(_2071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__B1 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__B2 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__4229__A1 (.DIODE(net1307));
 sky130_fd_sc_hd__diode_2 ANTENNA__4229__A2 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4229__B1 (.DIODE(_2076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4230__A1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__4230__A2 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA__4230__B2 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4232__A1 (.DIODE(net1306));
 sky130_fd_sc_hd__diode_2 ANTENNA__4232__B1 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA__4233__A2 (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4233__B1 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA__4235__A1 (.DIODE(net1305));
 sky130_fd_sc_hd__diode_2 ANTENNA__4235__A2 (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4235__B1 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA__4235__B2 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__A1 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__A2 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__B1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__B2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__A1 (.DIODE(net1304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__B1 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__B2 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__4239__A2 (.DIODE(_2091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4239__B1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA__4241__A1 (.DIODE(net1302));
 sky130_fd_sc_hd__diode_2 ANTENNA__4241__A2 (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4241__B1 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA__4241__B2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__A1 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__A2 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__B1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__B2 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__A1 (.DIODE(net1300));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__A2 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__B1 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__B2 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__4245__A2 (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4245__B1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__A1 (.DIODE(net1298));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__B1 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__A2 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__B1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__A1 (.DIODE(net1296));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__A2 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__B1 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__B2 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__A1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__A2 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__B1 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__B2 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__A1 (.DIODE(net1295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__B1 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__A1 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__A2 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__B1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__A1 (.DIODE(\u_reg.reg_rdata[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__B1 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA__4257__A2 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA__4257__B1 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA__4257__B2 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__A1 (.DIODE(\u_reg.reg_rdata[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__A2 (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__B1 (.DIODE(_2126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4260__A1 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__4260__A2 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA__4260__B2 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA__4262__A1 (.DIODE(net1293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4262__B1 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__A1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__A2 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__B1 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__B2 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__A1 (.DIODE(net1291));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__B1 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__B2 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__4266__A1 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__4266__A2 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA__4266__B1 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA__4266__B2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__A1 (.DIODE(net1290));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__A2 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__B1 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__B2 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__A1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__A2 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__B1 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__B2 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__A1 (.DIODE(\u_reg.reg_rdata[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__B1 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__B2 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__A2 (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__B1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA__4274__A1 (.DIODE(net1289));
 sky130_fd_sc_hd__diode_2 ANTENNA__4274__B1 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__A2 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__B1 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA__4277__A1 (.DIODE(net1288));
 sky130_fd_sc_hd__diode_2 ANTENNA__4277__B1 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__A2 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__B2 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__A1 (.DIODE(net1286));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__B1 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__A2 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__B1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__A1 (.DIODE(net1285));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__A2 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__B1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__B2 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__A1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__A2 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__B1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__B2 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__A1 (.DIODE(net1284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__A2 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__B1 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__B2 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__4287__A2 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA__4287__B1 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__A1 (.DIODE(net1282));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__A2 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__B1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__B2 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__A1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__B1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__B2 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__A1 (.DIODE(net1281));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__A2 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__B1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__B2 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__A1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__A2 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__B1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__B2 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__4295__A1 (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA__4295__B1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__A2 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__B1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__A1 (.DIODE(net1366));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__A2 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__B1 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__B2 (.DIODE(\u_reg.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__C (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__A1 (.DIODE(\u_s0.u_sync_wbb.wbm_lack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__A2 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__B1 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__B2 (.DIODE(net1401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__A1 (.DIODE(net1367));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__B1 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__B2 (.DIODE(\u_reg.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__A1 (.DIODE(\u_s0.u_sync_wbb.wbm_ack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__A2 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__B1 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__B2 (.DIODE(net1402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__A1 (.DIODE(net1312));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__B1 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__A2 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__B2 (.DIODE(net1140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__A1 (.DIODE(\u_reg.reg_rdata[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__A2 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__B1 (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__B2 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__A1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__A2 (.DIODE(_2036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__B1 (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__B2 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__A1 (.DIODE(\u_reg.reg_rdata[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__B1 (.DIODE(net1134));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__A2 (.DIODE(net1129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__B2 (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA__4314__A1 (.DIODE(\u_reg.reg_rdata[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4314__A2 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4314__B1 (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4314__B2 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__A1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__A2 (.DIODE(_2046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__B1 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__B2 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__A1 (.DIODE(net1311));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__B1 (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4318__A2 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__4318__B2 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__A1 (.DIODE(net1310));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__A2 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__B1 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__B2 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__A1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__A2 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__B1 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__B2 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__A1 (.DIODE(\u_reg.reg_rdata[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__A2 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__B1 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__A2 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__B1 (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__A1 (.DIODE(net1309));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__B1 (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__A1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__A2 (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__B1 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__A1 (.DIODE(net1308));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__A2 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__B1 (.DIODE(_2071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__B2 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__A1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__A2 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__B1 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__B2 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__A1 (.DIODE(net1307));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__B1 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__A2 (.DIODE(_2076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__B1 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA__4335__A1 (.DIODE(net1306));
 sky130_fd_sc_hd__diode_2 ANTENNA__4335__B1 (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__A2 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__B1 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA__4338__A1 (.DIODE(net1305));
 sky130_fd_sc_hd__diode_2 ANTENNA__4338__B1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__A1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__A2 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__B1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__B2 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__A1 (.DIODE(net1304));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__B1 (.DIODE(_2091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__A2 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__B1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__A1 (.DIODE(net1302));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__A2 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__B1 (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__B2 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__A1 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__A2 (.DIODE(_2096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__B1 (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__B2 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__A1 (.DIODE(net1300));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__A2 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__B1 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__B2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__A1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__A2 (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__B1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__A1 (.DIODE(net1298));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__B1 (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__A2 (.DIODE(_2104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__B1 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__A1 (.DIODE(net1296));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__A2 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__B1 (.DIODE(_2111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__A2 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__B1 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA__4356__A1 (.DIODE(net1295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4356__A2 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4356__B1 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__A1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__A2 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__B1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__B2 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__4359__A1 (.DIODE(\u_reg.reg_rdata[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4359__A2 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4359__B1 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA__4359__B2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__A1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__A2 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__B1 (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__A1 (.DIODE(\u_reg.reg_rdata[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__B1 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA__4363__A2 (.DIODE(_2126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4363__B1 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA__4365__A1 (.DIODE(net1293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4365__B1 (.DIODE(_2131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A2 (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__B1 (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__A1 (.DIODE(net1291));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__A2 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__B1 (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__B2 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__A1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__A2 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__B1 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__B2 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__A1 (.DIODE(net1290));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__A2 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__B1 (.DIODE(_2139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__B2 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__4372__A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__4372__A2 (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA__4372__B2 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__A1 (.DIODE(\u_reg.reg_rdata[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__B1 (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA__4375__A2 (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4375__B1 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA__4377__A1 (.DIODE(net1289));
 sky130_fd_sc_hd__diode_2 ANTENNA__4377__A2 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4377__B1 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA__4378__A1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__4378__A2 (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA__4378__B2 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA__4380__A1 (.DIODE(net1288));
 sky130_fd_sc_hd__diode_2 ANTENNA__4380__B1 (.DIODE(_2156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4380__B2 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__A1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__A2 (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__B1 (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__A1 (.DIODE(net1286));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__B1 (.DIODE(_2161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4384__A2 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA__4384__B1 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__A1 (.DIODE(net1285));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__A2 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__B1 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__B2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__A2 (.DIODE(_2166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__B1 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__A1 (.DIODE(net1284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__B1 (.DIODE(_2169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__A2 (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__B2 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__A1 (.DIODE(net1282));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__A2 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__B1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__B2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__4393__A2 (.DIODE(_2176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4393__B1 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__A1 (.DIODE(net1281));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__A2 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__B1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__B2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__4396__A2 (.DIODE(_2181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4396__B1 (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__A1 (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__A2 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__B1 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__B2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__A2 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__B1 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__A1 (.DIODE(\u_dcg_s0.cfg_mode_ss[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__A3 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__B1 (.DIODE(\u_dcg_s0.cfg_mode_ss[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__A1 (.DIODE(\u_dcg_s0.cfg_mode_ss[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__B1 (.DIODE(\u_dcg_s0.cfg_mode_ss[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__S0 (.DIODE(net1397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__S1 (.DIODE(net1390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4405__A1 (.DIODE(_2329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4405__S (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__S0 (.DIODE(net1398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__S1 (.DIODE(net1391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__A1 (.DIODE(_2330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__S (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__S0 (.DIODE(net1396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__S1 (.DIODE(net1389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__A1 (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__S (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__S0 (.DIODE(net1393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__S1 (.DIODE(net1386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__A1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__S (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__S0 (.DIODE(net1394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__S1 (.DIODE(net1388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__A1 (.DIODE(_2333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__S (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__S0 (.DIODE(net1395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__S1 (.DIODE(net1388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__A1 (.DIODE(_2334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__S (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__S0 (.DIODE(net1397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__S1 (.DIODE(net1390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__A1 (.DIODE(_2335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__S (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__S0 (.DIODE(net1394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__S1 (.DIODE(net1387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__S (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__S0 (.DIODE(net1397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__S1 (.DIODE(net1390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__S (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__S0 (.DIODE(net1395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__S1 (.DIODE(net1388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__A1 (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__S (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA__4424__A0 (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.mem[0][24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4424__S0 (.DIODE(net1395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4424__S1 (.DIODE(net1387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__A1 (.DIODE(_2339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__S (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__S0 (.DIODE(net1397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__S1 (.DIODE(net1390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4427__A1 (.DIODE(_2340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4427__S (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__S0 (.DIODE(net1393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__S1 (.DIODE(net1386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__A1 (.DIODE(_2341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__S (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__S0 (.DIODE(net1394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__S1 (.DIODE(net1387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__A1 (.DIODE(_2342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__S (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__A3 (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.mem[3][28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__S0 (.DIODE(net1397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__S1 (.DIODE(net1390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__A1 (.DIODE(_2343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__S (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__S0 (.DIODE(net1393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__S1 (.DIODE(net1386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__A1 (.DIODE(_2344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__S (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__S0 (.DIODE(net1394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__S1 (.DIODE(net1387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__A1 (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__S (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__S0 (.DIODE(net1392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__S1 (.DIODE(net1385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__A1 (.DIODE(_2346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__S (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__S0 (.DIODE(net1396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__S1 (.DIODE(net1389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__A1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__S (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__S0 (.DIODE(net1396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__S1 (.DIODE(net1389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4443__A1 (.DIODE(_2348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4443__S (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__S0 (.DIODE(net1396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__S1 (.DIODE(net1389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__A1 (.DIODE(_2349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__S (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__S0 (.DIODE(net1396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__S1 (.DIODE(net1389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__A1 (.DIODE(_2350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__S (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__S0 (.DIODE(net1397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__S1 (.DIODE(net1390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__A1 (.DIODE(_2351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__S (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__S0 (.DIODE(net1397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__S1 (.DIODE(net1390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__A1 (.DIODE(_2352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__S (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__S0 (.DIODE(net1392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__S1 (.DIODE(net1385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__A1 (.DIODE(_2353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__S (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__S0 (.DIODE(net1392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__S1 (.DIODE(net1385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__A1 (.DIODE(_2354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__S (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__S0 (.DIODE(net1393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__S1 (.DIODE(net1386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__A1 (.DIODE(_2355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__S (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__S0 (.DIODE(net1392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__S1 (.DIODE(net1385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__A1 (.DIODE(_2356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__S (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__S0 (.DIODE(net1393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__S1 (.DIODE(net1386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__A1 (.DIODE(_2357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__S (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__S0 (.DIODE(net1395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__S1 (.DIODE(net1388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__A1 (.DIODE(_2358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__S (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__S0 (.DIODE(net1398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__S1 (.DIODE(net1390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__A1 (.DIODE(_2359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__S (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__S0 (.DIODE(net1399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__S1 (.DIODE(net1391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__A1 (.DIODE(_2360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__S (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__S0 (.DIODE(net1392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__S1 (.DIODE(net1385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__A1 (.DIODE(_2361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__S (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__S0 (.DIODE(net1392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__S1 (.DIODE(net1385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__A1 (.DIODE(_2362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__S (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__S0 (.DIODE(net1394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__S1 (.DIODE(net1387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__A1 (.DIODE(_2363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__S (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__S0 (.DIODE(net1392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__S1 (.DIODE(net1386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__A1 (.DIODE(_2364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__S (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__A0 (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.mem[0][53] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__S0 (.DIODE(net1394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__S1 (.DIODE(net1387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__A1 (.DIODE(_2365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__S (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__S0 (.DIODE(net1394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__S1 (.DIODE(net1387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__A1 (.DIODE(_2366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__S (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__A2 (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.mem[2][55] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__S0 (.DIODE(net1394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__S1 (.DIODE(net1387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__A1 (.DIODE(_2367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__S (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__S0 (.DIODE(net1393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__S1 (.DIODE(net1386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__A1 (.DIODE(_2368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__S (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__S0 (.DIODE(net1395));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__S1 (.DIODE(net1388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__A1 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__S (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__S0 (.DIODE(net1392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__S1 (.DIODE(net1385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__A1 (.DIODE(_2370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__S (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__S0 (.DIODE(net1394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__S1 (.DIODE(net1387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4489__A1 (.DIODE(_2371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4489__S (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__A1 (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.mem[1][60] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__S0 (.DIODE(net1393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__S1 (.DIODE(net1385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__A1 (.DIODE(_2372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__S (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__S0 (.DIODE(net1392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__S1 (.DIODE(net1385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__A1 (.DIODE(_2373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__S (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__S0 (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__S1 (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__A1 (.DIODE(_2374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__S (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__S0 (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__S1 (.DIODE(net1353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__A1 (.DIODE(_2375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__S (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__S0 (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__S1 (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__S (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__S0 (.DIODE(net1363));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__S1 (.DIODE(net1356));
 sky130_fd_sc_hd__diode_2 ANTENNA__4501__S (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__S0 (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__S1 (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__A1 (.DIODE(_2378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__S (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__S0 (.DIODE(net1363));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__S1 (.DIODE(net1356));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__A1 (.DIODE(_2379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__S (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__S0 (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__S1 (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__S0 (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__S1 (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__S (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__S0 (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__S1 (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__A1 (.DIODE(_2382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__S0 (.DIODE(net1363));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__S1 (.DIODE(net1356));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__A1 (.DIODE(_2383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__S (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__S0 (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__S1 (.DIODE(net1353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__S (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__S0 (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__S1 (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__S (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__S0 (.DIODE(net1363));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__S1 (.DIODE(net1356));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__A1 (.DIODE(_2386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__S0 (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__S1 (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__A1 (.DIODE(_2387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__S0 (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__S1 (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__S (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__S0 (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__S1 (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__A1 (.DIODE(_2389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__S (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__S0 (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__S1 (.DIODE(net1358));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__S (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__S0 (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__S1 (.DIODE(net1353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__S (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__S0 (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__S1 (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__A1 (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__S (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__S0 (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__S1 (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__S (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__S0 (.DIODE(net1363));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__S1 (.DIODE(net1356));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__A1 (.DIODE(_2394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__S (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__S0 (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__S1 (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__A1 (.DIODE(_2395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__S0 (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__S1 (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__S (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__S0 (.DIODE(net1363));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__S1 (.DIODE(net1356));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__A1 (.DIODE(_2397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__S (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__S0 (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__S1 (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__S (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__S0 (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__S1 (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__A1 (.DIODE(_2399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__S (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__S0 (.DIODE(net1361));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__S1 (.DIODE(net1354));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__S (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__S0 (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__S1 (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__S0 (.DIODE(net1363));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__S1 (.DIODE(net1356));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__A1 (.DIODE(_2402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__S (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__S0 (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__S1 (.DIODE(net1353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__A1 (.DIODE(_2403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__S (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__S0 (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__S1 (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__S (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__S0 (.DIODE(net1365));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__S1 (.DIODE(net1358));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__S (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__S0 (.DIODE(net1365));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__S1 (.DIODE(net1358));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__A1 (.DIODE(_2406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__S (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__S0 (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__S1 (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__S (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__S0 (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__S1 (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__A1 (.DIODE(_2408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__S (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__S0 (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__S1 (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__S (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__S0 (.DIODE(net1361));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__S1 (.DIODE(net1354));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__S (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__S0 (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__S1 (.DIODE(net1353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__S (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__S0 (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__S1 (.DIODE(net1353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__S (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__S0 (.DIODE(net1361));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__S1 (.DIODE(net1354));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__S (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__S0 (.DIODE(net1361));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__S1 (.DIODE(net1354));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__A1 (.DIODE(_2414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__S (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__S0 (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__S1 (.DIODE(net1353));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__S (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__S0 (.DIODE(net1361));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__S1 (.DIODE(net1354));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__S (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__A_N (.DIODE(_1719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__B (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__A0 (.DIODE(s0_wbd_lack_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__A1 (.DIODE(s0_wbd_ack_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__A (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__B (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__A (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__B (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__C_N (.DIODE(net2049));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__A (.DIODE(_2423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__A (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__D (.DIODE(_2423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__A1 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__S0 (.DIODE(net1338));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__S1 (.DIODE(net1328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__A1 (.DIODE(_2426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__S (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__S0 (.DIODE(net1342));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__S1 (.DIODE(net1332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__A1 (.DIODE(_2427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__S (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__S0 (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__S1 (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__A1 (.DIODE(_2428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__S0 (.DIODE(net1335));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__S1 (.DIODE(net1325));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__A1 (.DIODE(_2429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__S (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__S0 (.DIODE(net1335));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__S1 (.DIODE(net1325));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__S0 (.DIODE(net1340));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__S1 (.DIODE(net1330));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__S (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__S0 (.DIODE(net1340));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__S1 (.DIODE(net1330));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__S (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__S0 (.DIODE(net1341));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__S1 (.DIODE(net1331));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__S (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__S0 (.DIODE(net1340));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__S1 (.DIODE(net1330));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__S (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__S0 (.DIODE(net1338));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__S1 (.DIODE(net1328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__S (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__S0 (.DIODE(net1339));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__S1 (.DIODE(net1329));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__A1 (.DIODE(_2436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__S (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__S0 (.DIODE(net1339));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__S1 (.DIODE(net1329));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__S (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__S0 (.DIODE(net1337));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__S1 (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__A1 (.DIODE(_2438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__S (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__S0 (.DIODE(net1339));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__S1 (.DIODE(net1329));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__A1 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__S (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__S0 (.DIODE(net1341));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__S1 (.DIODE(net1331));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__S (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__S0 (.DIODE(net1340));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__S1 (.DIODE(net1330));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__A1 (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__S (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__S0 (.DIODE(net1341));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__S1 (.DIODE(net1331));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__S (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__S0 (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__S1 (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__S (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__S0 (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__S1 (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__S (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__S0 (.DIODE(net1341));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__S1 (.DIODE(net1331));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__S (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__S0 (.DIODE(net1338));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__S1 (.DIODE(net1328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__A1 (.DIODE(_2446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__S (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__S0 (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__S1 (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__A1 (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__S (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__S0 (.DIODE(net1340));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__S1 (.DIODE(net1330));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__A1 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__S (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__S0 (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__S1 (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__S (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__S0 (.DIODE(net1338));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__S1 (.DIODE(net1328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__S (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__S0 (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__S1 (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__S (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__S0 (.DIODE(net1339));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__S1 (.DIODE(net1329));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__S (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__S0 (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__S1 (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__S (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__S0 (.DIODE(net1339));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__S1 (.DIODE(net1329));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__A1 (.DIODE(_2454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__S (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__S0 (.DIODE(net1337));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__S1 (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__A1 (.DIODE(_2455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__S (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__S0 (.DIODE(net1338));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__S1 (.DIODE(net1328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__A1 (.DIODE(_2456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__S (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__S0 (.DIODE(net1337));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__S1 (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__S (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__S0 (.DIODE(net1337));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__S1 (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__A1 (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__S (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__S0 (.DIODE(net1335));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__S1 (.DIODE(net1325));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__S0 (.DIODE(net1337));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__S1 (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__A1 (.DIODE(_2460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__S (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__S0 (.DIODE(net1338));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__S1 (.DIODE(net1328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__A1 (.DIODE(_2461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__S (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__S0 (.DIODE(net1335));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__S1 (.DIODE(net1325));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__A1 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__S (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__S0 (.DIODE(net1338));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__S1 (.DIODE(net1328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__A1 (.DIODE(_2463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__S (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__S0 (.DIODE(net1342));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__S1 (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__A1 (.DIODE(_2464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__S (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__S0 (.DIODE(net1338));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__S1 (.DIODE(net1328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__A1 (.DIODE(_2465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__S (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__S0 (.DIODE(net1337));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__S1 (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__A1 (.DIODE(_2466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__S (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__S0 (.DIODE(net1335));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__S1 (.DIODE(net1325));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__S (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__S0 (.DIODE(net1333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__S1 (.DIODE(net1325));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__S0 (.DIODE(net1337));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__S1 (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__A1 (.DIODE(_2469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__S (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__S0 (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__S1 (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__A1 (.DIODE(_2470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__S (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__S0 (.DIODE(net1337));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__S1 (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__A1 (.DIODE(_2471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__S (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__S0 (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__S1 (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__A1 (.DIODE(_2472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__S (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__S0 (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__S1 (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__A1 (.DIODE(_2473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__S (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__S0 (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__S1 (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__A1 (.DIODE(_2474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__S (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__S0 (.DIODE(net1333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__S1 (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__A1 (.DIODE(_2475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__S0 (.DIODE(net1333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__S1 (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__A1 (.DIODE(_2476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__S0 (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__S1 (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__A1 (.DIODE(_2477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__S0 (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__S1 (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__A1 (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__S0 (.DIODE(net1333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__S1 (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__S0 (.DIODE(net1333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__S1 (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__S0 (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__S1 (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__A1 (.DIODE(_2481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__S (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__S0 (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__S1 (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__A1 (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__S (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__S0 (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__S1 (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__A1 (.DIODE(_2483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__S (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__S0 (.DIODE(net1333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__S1 (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__A1 (.DIODE(_2484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__S0 (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__S1 (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__A1 (.DIODE(_2485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__S (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__S0 (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__S1 (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__A1 (.DIODE(_2486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__S0 (.DIODE(net1333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__S1 (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__A1 (.DIODE(_2487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__S0 (.DIODE(net1333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__S1 (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__A1 (.DIODE(_2488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__S (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__S0 (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__S1 (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__A1 (.DIODE(_2489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__S0 (.DIODE(net1333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__S1 (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__A1 (.DIODE(_2490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__S0 (.DIODE(net1333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__S1 (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__A1 (.DIODE(_2491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__S0 (.DIODE(net1335));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__S1 (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__A1 (.DIODE(_2492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__S (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__A (.DIODE(\u_s0.u_sync_wbb.wbm_lack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__B (.DIODE(net1208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__A (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__B (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__A (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__B (.DIODE(_1958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__A (.DIODE(net1366));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__B (.DIODE(net1185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__A1 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__A2 (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__B1 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__B2 (.DIODE(\u_reg.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__A1 (.DIODE(net1366));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__A2 (.DIODE(net1185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__A3 (.DIODE(_1853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__A1 (.DIODE(net1401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__A2 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__A (.DIODE(net1401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__B (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__A (.DIODE(net1185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__B (.DIODE(_1853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__A1 (.DIODE(\u_reg.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__B1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__B2 (.DIODE(net1367));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__A1 (.DIODE(\u_s0.u_sync_wbb.wbm_ack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__B2 (.DIODE(net1402));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__A1 (.DIODE(net1312));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__A2 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__B1 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__B2 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__A1 (.DIODE(net1141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__B2 (.DIODE(net1139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__A (.DIODE(_2504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__A1 (.DIODE(\u_reg.reg_rdata[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__A2 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__B1 (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__B2 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__A1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__A2 (.DIODE(_2036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__B1 (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__B2 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__A1 (.DIODE(\u_reg.reg_rdata[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__A2 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__B1 (.DIODE(net1134));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__B2 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__A1 (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__A2 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__B2 (.DIODE(net1130));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__A1 (.DIODE(\u_reg.reg_rdata[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__A2 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__B1 (.DIODE(_2046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__B2 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__A1 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__B1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__B2 (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__A1 (.DIODE(net1311));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__A2 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__B1 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__A2 (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__B1 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__A1 (.DIODE(\u_reg.reg_rdata[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__A2 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__B1 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__B2 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__A2 (.DIODE(_2056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__B1 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__B2 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__A1 (.DIODE(\u_reg.reg_rdata[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__B1 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__A1 (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__B1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__B2 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__A2 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__B1 (.DIODE(_2064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__B2 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__A1 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__A2 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__B1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__B2 (.DIODE(_2067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__A1 (.DIODE(\u_reg.reg_rdata[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__A2 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__B1 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__A2 (.DIODE(_2071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__B1 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__A2 (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__B1 (.DIODE(_2074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__B2 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__A2 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__B1 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__B2 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__A1 (.DIODE(\u_reg.reg_rdata[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__A2 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__B1 (.DIODE(_2079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__B2 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__A2 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__B1 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__A1 (.DIODE(net1305));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__A2 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__B1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__B2 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__A1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__A2 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__B1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__A1 (.DIODE(\u_reg.reg_rdata[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__A2 (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__B1 (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__B2 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__A1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__A2 (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__B1 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__B2 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__A1 (.DIODE(net1303));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__A2 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__B1 (.DIODE(_2094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__A2 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__B1 (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__A1 (.DIODE(net1301));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__A2 (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__B1 (.DIODE(_2099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__B2 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__A1 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__A2 (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__B1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__B2 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__A1 (.DIODE(net1299));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__A2 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__B1 (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__B2 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__A1 (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__A2 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__B2 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__A1 (.DIODE(net1297));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__A2 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__B1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__B2 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__A2 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__B1 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__A1 (.DIODE(net1295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__A2 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__B1 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__A2 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__B1 (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__A1 (.DIODE(\u_reg.reg_rdata[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__A2 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__B1 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__B2 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__A1 (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__B1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__B2 (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__A1 (.DIODE(\u_reg.reg_rdata[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__A2 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__B1 (.DIODE(_2126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__B2 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__A1 (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__A2 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__B1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__B2 (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__A1 (.DIODE(net1294));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__A2 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__B1 (.DIODE(_2129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__B2 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__A2 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__B1 (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__A1 (.DIODE(net1292));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__B1 (.DIODE(_2137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__B2 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__A2 (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__B1 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__B1 (.DIODE(_2142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__B2 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__A2 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__B1 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__B2 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__A1 (.DIODE(\u_reg.reg_rdata[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__A2 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__B1 (.DIODE(_2144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__B2 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__A1 (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__A2 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__B2 (.DIODE(_2147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4808__A (.DIODE(_2550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4808__B (.DIODE(_2551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__A1 (.DIODE(net1289));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__A2 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__B1 (.DIODE(_2152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__A2 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__B1 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__B2 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__A1 (.DIODE(\u_reg.reg_rdata[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__A2 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__B1 (.DIODE(_2154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__B2 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__A2 (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__B1 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__B2 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__A1 (.DIODE(net1287));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__A2 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__B1 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__A1 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__B1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__B2 (.DIODE(_2159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__A1 (.DIODE(\u_reg.reg_rdata[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__A2 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__B1 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__A1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__B1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__B2 (.DIODE(_2164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__A1 (.DIODE(\u_reg.reg_rdata[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__A2 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__B1 (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__A2 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__B1 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__A1 (.DIODE(net1283));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__B1 (.DIODE(_2174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__B2 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__A1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__A2 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__B1 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__A1 (.DIODE(\u_reg.reg_rdata[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__A2 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__B1 (.DIODE(_2179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__B2 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__A1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__A2 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__B1 (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__A1 (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__A2 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__B1 (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__A1 (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__B1 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__B2 (.DIODE(_2187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__A2 (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.mem[2][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__S0 (.DIODE(net1397));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__S1 (.DIODE(net1390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__S (.DIODE(net1502));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__S0 (.DIODE(net1396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__S1 (.DIODE(net1391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__S (.DIODE(net1501));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__S0 (.DIODE(net1398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__S1 (.DIODE(net1391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__S (.DIODE(net1501));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__S0 (.DIODE(net1398));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__S1 (.DIODE(net1391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__A1 (.DIODE(_2571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__S (.DIODE(net1501));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__S0 (.DIODE(net1392));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__S1 (.DIODE(net1385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__A1 (.DIODE(net1816));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__S (.DIODE(net1501));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__S0 (.DIODE(net1396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__S1 (.DIODE(net1389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__A1 (.DIODE(_2573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__S (.DIODE(net1501));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__A1 (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.mem[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__S0 (.DIODE(net1393));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__S1 (.DIODE(net1386));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__A1 (.DIODE(net1804));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__S (.DIODE(net1502));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__S0 (.DIODE(net1394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__S1 (.DIODE(net1387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__A1 (.DIODE(_2575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__S (.DIODE(net1501));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__S0 (.DIODE(net1396));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__S1 (.DIODE(net1389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__A0 (.DIODE(\u_s2.u_sync_wbb.s_cmd_rd_data_l[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__A1 (.DIODE(_2576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__S (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__A1 (.DIODE(_2329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__S (.DIODE(net1496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__A1 (.DIODE(_2330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__S (.DIODE(net1502));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__A1 (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__S (.DIODE(net1500));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__A1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__S (.DIODE(net1495));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__A1 (.DIODE(_2333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__S (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__A1 (.DIODE(_2334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__S (.DIODE(net1502));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__A1 (.DIODE(_2335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__S (.DIODE(net1500));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__S (.DIODE(net1496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__S (.DIODE(net1502));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__A1 (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__S (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__A1 (.DIODE(_2339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__S (.DIODE(net1497));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__A1 (.DIODE(_2340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__S (.DIODE(net1500));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__A1 (.DIODE(_2341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__S (.DIODE(net1496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__A1 (.DIODE(_2342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__S (.DIODE(net1497));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__A1 (.DIODE(_2343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__S (.DIODE(net1501));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__A1 (.DIODE(_2344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__S (.DIODE(net1496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__A1 (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__S (.DIODE(net1496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__A1 (.DIODE(_2346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__S (.DIODE(net1495));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__A1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__S (.DIODE(net1497));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__A1 (.DIODE(_2348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__S (.DIODE(net1500));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__A1 (.DIODE(_2349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__S (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__A1 (.DIODE(_2350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__S (.DIODE(net1500));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__A1 (.DIODE(_2351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__S (.DIODE(net1500));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__A1 (.DIODE(_2352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__S (.DIODE(net1496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__A1 (.DIODE(_2353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__S (.DIODE(net1500));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__A1 (.DIODE(_2354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__S (.DIODE(net1495));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__A1 (.DIODE(_2355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__S (.DIODE(net1498));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__A1 (.DIODE(_2356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__S (.DIODE(net1496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__A1 (.DIODE(_2357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__S (.DIODE(net1495));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__A1 (.DIODE(_2358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__S (.DIODE(net1495));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__A1 (.DIODE(_2359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__S (.DIODE(net1500));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__A1 (.DIODE(_2360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__S (.DIODE(net1497));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__A1 (.DIODE(_2361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__S (.DIODE(net1495));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__A1 (.DIODE(_2362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__S (.DIODE(net1497));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__A1 (.DIODE(_2363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__S (.DIODE(net1496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__A1 (.DIODE(_2364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__S (.DIODE(net1496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__S (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__A1 (.DIODE(_2365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__S (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__A1 (.DIODE(_2366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__S (.DIODE(net1496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__A1 (.DIODE(_2367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__S (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__A1 (.DIODE(_2368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__S (.DIODE(net1495));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__A1 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__S (.DIODE(net1495));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__A1 (.DIODE(_2370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__S (.DIODE(net1495));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__A1 (.DIODE(_2371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__S (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__S (.DIODE(net1498));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__S (.DIODE(net1495));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__A1 (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__B2 (.DIODE(net1409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__A (.DIODE(net1407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__B (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__A (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__C (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__A1 (.DIODE(net1407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__A2 (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__B1 (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__A1 (.DIODE(_1962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__A1 (.DIODE(net1409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__B1 (.DIODE(net1224));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__A1 (.DIODE(m3_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__A2 (.DIODE(_1958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A1 (.DIODE(_1967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A2 (.DIODE(_1970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__B1 (.DIODE(net1401));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__A0 (.DIODE(net1409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__A1_N (.DIODE(net1224));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__B1 (.DIODE(_1962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__B2 (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__B (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__A0 (.DIODE(net1407));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__A (.DIODE(\u_s0.u_sync_wbb.m_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__A (.DIODE(\u_s0.u_sync_wbb.m_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__A (.DIODE(\u_s0.u_sync_wbb.m_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__B (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__A1 (.DIODE(\u_s0.u_sync_wbb.m_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__B2 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__A2 (.DIODE(_1735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__B1 (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__A (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__A1 (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__B1 (.DIODE(_2589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__A2 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__C1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__A2 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__A1 (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__B1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__A (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__B (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4922__C1 (.DIODE(_2589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__B (.DIODE(\u_s0.u_sync_wbb.m_bl_cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__B (.DIODE(\u_s0.u_sync_wbb.m_bl_cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4925__A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA__4925__B1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__B1 (.DIODE(\u_s0.u_sync_wbb.m_bl_cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__B2 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__B1 (.DIODE(_1792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__A (.DIODE(_1792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__A (.DIODE(_2589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__B (.DIODE(\u_s0.u_sync_wbb.m_bl_cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__B1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__B2 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__A1 (.DIODE(_1792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__B1 (.DIODE(_1794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__B1 (.DIODE(_2589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__A (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__S (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__A2 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__B1 (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__A (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4943__A (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__4943__B (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__C1 (.DIODE(_2589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__S (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__A (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__B (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__C (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4949__A1 (.DIODE(_1998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4949__A2 (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4949__B1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__A (.DIODE(_2589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__B1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__B2 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__A1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__A2 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__A3 (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__B1 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__A (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__B (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__C (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__D (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4957__A (.DIODE(_2589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A1 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A2 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A3 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A4 (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__B1 (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__C (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__D (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__C (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__D (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__B1 (.DIODE(_2589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__A1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__B2 (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__C1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__A1 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__A2 (.DIODE(_1998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__A3 (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__B1 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__A (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__B (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__C (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__D (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__A (.DIODE(_2589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__A1 (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__A (.DIODE(net1223));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__B (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__A_N (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__B (.DIODE(m1_wbd_adr_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__C (.DIODE(net1276));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__A (.DIODE(net1276));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__B (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__C (.DIODE(m3_wbd_adr_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__A_N (.DIODE(net1276));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__B (.DIODE(m2_wbd_adr_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__A (.DIODE(net1276));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__B (.DIODE(\u_wbi_arb.gnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__C (.DIODE(net1597));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__A1 (.DIODE(_2019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__A (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__B (.DIODE(net1274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__C (.DIODE(m2_wbd_adr_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__A1 (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__A2 (.DIODE(m1_wbd_adr_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__B2 (.DIODE(m3_wbd_adr_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__C1 (.DIODE(_2019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__A1 (.DIODE(net1596));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__A2 (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__A_N (.DIODE(net1274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__B (.DIODE(m1_wbd_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__C (.DIODE(net1277));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__A (.DIODE(net1277));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__B (.DIODE(net1274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__C (.DIODE(m3_wbd_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__A_N (.DIODE(net1277));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__B (.DIODE(m2_wbd_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__A (.DIODE(net1276));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__B (.DIODE(net1274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__C (.DIODE(net1598));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__A1 (.DIODE(net1152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__A1 (.DIODE(net1152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__A (.DIODE(_2653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__B (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__C (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__A0 (.DIODE(m0_wbd_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__A1 (.DIODE(m1_wbd_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__A2 (.DIODE(m2_wbd_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__A3 (.DIODE(m3_wbd_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__S0 (.DIODE(net1276));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__S1 (.DIODE(net1274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__A_N (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__B (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__A (.DIODE(m1_wbd_sel_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__B (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__A1 (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__A2 (.DIODE(m2_wbd_sel_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__B2 (.DIODE(m3_wbd_sel_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__C1 (.DIODE(_2019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__A1 (.DIODE(m0_wbd_sel_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__A2 (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__A_N (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__B (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__C (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__D (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__A (.DIODE(net1586));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__B (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__A2 (.DIODE(net1555));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__B1 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__A2 (.DIODE(net1529));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__S (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A (.DIODE(net1585));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__B (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__A2 (.DIODE(net1554));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__B1 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A2 (.DIODE(net1528));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__A1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__S (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__A (.DIODE(net1584));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__B (.DIODE(net1152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__A1 (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__A2 (.DIODE(m2_wbd_dat_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__B1 (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__A1 (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__A2 (.DIODE(net1553));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__B1 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__A1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__S (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__A (.DIODE(net1583));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__B (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__A1 (.DIODE(net1221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__A2 (.DIODE(net1527));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__A1 (.DIODE(net1221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__A2 (.DIODE(net1552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__A1 (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__S (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__A (.DIODE(net1581));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__B (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__A2 (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__B1 (.DIODE(net1221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__A2 (.DIODE(net1526));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__A1 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__S (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__A1 (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__A2 (.DIODE(net1549));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__B1 (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__A1 (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__A2 (.DIODE(net1525));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__B1 (.DIODE(net1580));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__B2 (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__A1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__S (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__A1 (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__A2 (.DIODE(net1548));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__B1 (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__A1 (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__A2 (.DIODE(net2051));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__B1 (.DIODE(net1579));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__B2 (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__A1 (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__S (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__A1 (.DIODE(net1212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__A2 (.DIODE(net1547));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__B1 (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A1 (.DIODE(net1212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A2 (.DIODE(net1524));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__B1 (.DIODE(net1578));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__B2 (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A1 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__S (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__A (.DIODE(_2661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__B (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__C_N (.DIODE(_2653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__A (.DIODE(net1276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__B (.DIODE(net1274));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__C (.DIODE(m3_wbd_sel_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__A1 (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__A2 (.DIODE(m2_wbd_sel_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__B1 (.DIODE(m1_wbd_sel_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__B2 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__C1 (.DIODE(_2019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A1 (.DIODE(net1565));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A2 (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__A_N (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__B (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__C (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__A1 (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__A2 (.DIODE(net1562));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__B1 (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__A1 (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__A2 (.DIODE(net2050));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__B1 (.DIODE(net1593));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__B2 (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__A1 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__S (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__A (.DIODE(net1582));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__B (.DIODE(net1152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__A1 (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__A2 (.DIODE(net1551));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__B1 (.DIODE(net1223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__A1 (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__A2 (.DIODE(m2_wbd_dat_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__A1 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__S (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__A (.DIODE(net1574));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__B (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__A1 (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__A2 (.DIODE(net1543));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__B1 (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__A1 (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__A2 (.DIODE(m2_wbd_dat_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A1 (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__S (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__A1 (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__A2 (.DIODE(m1_wbd_dat_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__B1 (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__A1 (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__A2 (.DIODE(net2088));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__B1 (.DIODE(m0_wbd_dat_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__B2 (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__A1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__S (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__A2 (.DIODE(net1540));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__B1 (.DIODE(net1221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__A2 (.DIODE(net1518));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__B1 (.DIODE(net1571));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__B2 (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__A1 (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__S (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__A2 (.DIODE(net1539));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__B1 (.DIODE(net1221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__A2 (.DIODE(net1517));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__B1 (.DIODE(net1570));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__B2 (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A1 (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__S (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__A (.DIODE(net1569));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__B (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__A1 (.DIODE(net1217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__A2 (.DIODE(net1538));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__B1 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A1 (.DIODE(net1217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A2 (.DIODE(net1516));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__A1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__S (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A2 (.DIODE(net1537));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__B1 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__A2 (.DIODE(net1515));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__B1 (.DIODE(net1568));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__B2 (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__A1 (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__S (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__A (.DIODE(net1276));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__B (.DIODE(net1274));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__C (.DIODE(m3_wbd_sel_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__A1 (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__A2 (.DIODE(m2_wbd_sel_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__B1 (.DIODE(m1_wbd_sel_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__B2 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__C1 (.DIODE(_2019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__A1 (.DIODE(m0_wbd_sel_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__A2 (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__A_N (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__B (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__C (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__A (.DIODE(net1567));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__B (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A1 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A2 (.DIODE(net1514));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__A1 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__A2 (.DIODE(net1536));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__A1 (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__S (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5071__A2 (.DIODE(net1535));
 sky130_fd_sc_hd__diode_2 ANTENNA__5071__B1 (.DIODE(net1223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__A2 (.DIODE(net1513));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__B1 (.DIODE(net1566));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__B2 (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__A1 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__S (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__A2 (.DIODE(net1561));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__B1 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__A2 (.DIODE(net1534));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__B1 (.DIODE(net1592));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__B2 (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__A1 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__S (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__A2 (.DIODE(net1560));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__B1 (.DIODE(net1221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__A2 (.DIODE(net1533));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__B1 (.DIODE(net1591));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__B2 (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__A1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__S (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__A2 (.DIODE(net1559));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__B1 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A2 (.DIODE(net1532));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__B1 (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__B2 (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__A1 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__S (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A1 (.DIODE(net1212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A2 (.DIODE(net1558));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__B1 (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__A1 (.DIODE(net1212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__A2 (.DIODE(m2_wbd_dat_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__B1 (.DIODE(net1589));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__B2 (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__A1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__S (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A1 (.DIODE(net1212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A2 (.DIODE(net1557));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__B1 (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__A1 (.DIODE(net1212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__A2 (.DIODE(net1531));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__B1 (.DIODE(net1588));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__B2 (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__A1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__S (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A1 (.DIODE(net1212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A2 (.DIODE(net1556));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__B1 (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__A1 (.DIODE(net1212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__A2 (.DIODE(net1530));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__B1 (.DIODE(net1587));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__B2 (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__A1 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__S (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__A_N (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__B (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__C (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__S (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__S (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__A1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__S (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A1 (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__S (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__A0 (.DIODE(\u_reg.reg_6[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__A1 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__S (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__A1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__S (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A1 (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__S (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A1 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__S (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__A (.DIODE(_2653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__B (.DIODE(_2661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A_N (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__B (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__C (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__A1 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__S (.DIODE(_2739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__A1 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__S (.DIODE(_2739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__A1 (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__S (.DIODE(_2739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__A1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__S (.DIODE(_2739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__A1 (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__S (.DIODE(_2739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A1 (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__S (.DIODE(_2739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__A1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__S (.DIODE(_2739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A1 (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__S (.DIODE(_2739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__A_N (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__C (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__A1 (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__S (.DIODE(_2740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__A1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__S (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A1 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__S (.DIODE(_2740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__A1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__S (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__A1 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__S (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__A1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__S (.DIODE(_2740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__A1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__S (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__A1 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__S (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__A_N (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__B (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__C (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__S (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A0 (.DIODE(\u_reg.reg_7[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__S (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__A1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__S (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__A1 (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__S (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A1 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__S (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__A1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__S (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__A1 (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__S (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__A1 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__S (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__A_N (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__B (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__C (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__D (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__A0 (.DIODE(\u_reg.reg_5[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__A1 (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__A1 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__S (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__A1 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__S (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__A0 (.DIODE(\u_reg.reg_5[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__A1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__S (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__A1 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__S (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__A1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__S (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__A1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__S (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__A1 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__S (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__A_N (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__B (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__C (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__D (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__A1 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__S (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__A1 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__S (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__A1 (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__A0 (.DIODE(\u_reg.reg_5[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__A1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A1 (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__S (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__A1 (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__S (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__A1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__S (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A1 (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__S (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__A (.DIODE(_2653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__B (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__C (.DIODE(_2661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__A_N (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__B (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__C (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__A0 (.DIODE(\u_reg.reg_4[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__S (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__A1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__S (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__A1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__S (.DIODE(_2745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__A1 (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__S (.DIODE(_2745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__A1 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__S (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__A1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__S (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__A1 (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__S (.DIODE(_2745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__A1 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__S (.DIODE(_2745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__A_N (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__C (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__A1 (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__S (.DIODE(_2746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__S (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__A1 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__S (.DIODE(_2746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__A1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__S (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__A1 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__S (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__A1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__S (.DIODE(_2746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__A1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__S (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__A1 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__S (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__A_N (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__B (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__C (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__A1 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__S (.DIODE(_2747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__A1 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__S (.DIODE(_2747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__A1 (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__S (.DIODE(_2747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__A1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__S (.DIODE(_2747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__A1 (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__S (.DIODE(_2747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__A1 (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__S (.DIODE(_2747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__A1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__S (.DIODE(_2747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__A1 (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__S (.DIODE(_2747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__A (.DIODE(_2653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__B (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__C (.DIODE(_2661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__A (.DIODE(net1223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__B (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__C (.DIODE(m2_wbd_sel_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__A1 (.DIODE(m3_wbd_sel_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__B1 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__B2 (.DIODE(m1_wbd_sel_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__A0 (.DIODE(m0_wbd_sel_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__S (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__A_N (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__B (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__C (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__A (.DIODE(m0_wbd_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__B (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__A1 (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__A2 (.DIODE(m1_wbd_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__B1 (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__A1 (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__A2 (.DIODE(m2_wbd_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__A1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__S (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__A1 (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__A2 (.DIODE(m1_wbd_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__B1 (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__A1 (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__A2 (.DIODE(m2_wbd_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__B1 (.DIODE(m0_wbd_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__B2 (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__A0 (.DIODE(\u_reg.reg_3[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__A1 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__S (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__A2 (.DIODE(net1546));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__B1 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__A2 (.DIODE(net1523));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__B1 (.DIODE(net1577));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__B2 (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__A1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__S (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__A2 (.DIODE(net1545));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__B1 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__A2 (.DIODE(net1522));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__B1 (.DIODE(net1576));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__B2 (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__A1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__S (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__A (.DIODE(m0_wbd_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__B (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A1 (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A2 (.DIODE(m1_wbd_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__B1 (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__A1 (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__S (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__A (.DIODE(net1575));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__B (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A1 (.DIODE(net1221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A2 (.DIODE(net1521));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__A1 (.DIODE(net1221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__A2 (.DIODE(net1544));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__A1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__S (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__A1 (.DIODE(net1212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__A2 (.DIODE(net1542));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__B1 (.DIODE(net1221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__A1 (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__A2 (.DIODE(net1520));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__B1 (.DIODE(net1573));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__B2 (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__S (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A (.DIODE(net1572));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__B (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__A2 (.DIODE(net1541));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__B1 (.DIODE(net1221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A2 (.DIODE(net1519));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__S (.DIODE(_2752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__A_N (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__C (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A1 (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__S (.DIODE(_2773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__A1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__S (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A1 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__S (.DIODE(_2773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__A1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__S (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__A1 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__S (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__A1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__S (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__A1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__S (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A1 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__S (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__A_N (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__B (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__C (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__A1 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__S (.DIODE(_2774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__A1 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__S (.DIODE(_2774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__A1 (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__S (.DIODE(_2774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__S (.DIODE(_2774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__A1 (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__S (.DIODE(_2774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__A1 (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__S (.DIODE(_2774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__S (.DIODE(_2774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__A1 (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__S (.DIODE(_2774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__A (.DIODE(_2653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__B (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__C (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__A_N (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__C (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__A1 (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__S (.DIODE(_2776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__A1 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__S (.DIODE(_2776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__A1 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__S (.DIODE(_2776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__A0 (.DIODE(\u_reg.reg_2[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__A1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__S (.DIODE(_2776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A1 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__S (.DIODE(_2776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__A1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__S (.DIODE(_2776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__A1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__S (.DIODE(_2776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__A1 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__S (.DIODE(_2776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__A_N (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__B (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__C (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__S (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__S (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__A1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__S (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__A1 (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__S (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__A1 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__S (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__S (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A1 (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__S (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A1 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__S (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__A_N (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__B (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__C (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__A1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__S (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A1 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__S (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__A1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__S (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__A1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__S (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__A1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__S (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__A1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__S (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__A1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A_N (.DIODE(_2653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__B (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__A (.DIODE(_2661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__B (.DIODE(_2779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A_N (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__C (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__A0 (.DIODE(\u_dcg_riscv.cfg_mode[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__A1 (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__S (.DIODE(_2781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A1 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__S (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__A1 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__S (.DIODE(_2781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__S (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__A1 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__S (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A1 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__S (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__A1 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__S (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__A1 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__S (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__A_N (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__B (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__C (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__S (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__A1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__S (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__A1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__S (.DIODE(_2782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__A1 (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__S (.DIODE(_2782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__A1 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__S (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__A1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__S (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__A1 (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__S (.DIODE(_2782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__S (.DIODE(_2782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__A_N (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__B (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__C (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__S (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A0 (.DIODE(\u_reg.cfg_dcg_ctrl[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A1 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__S (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__S (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__A1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__S (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__S (.DIODE(_2783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__S (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__S (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__A1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__S (.DIODE(_2783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A (.DIODE(_1711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__B (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__C_N (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__B (.DIODE(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A0 (.DIODE(net1802));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__S (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A0 (.DIODE(net1805));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__S (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A0 (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__S (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__A0 (.DIODE(net1795));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__S (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A0 (.DIODE(net1779));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__S (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__A0 (.DIODE(net1796));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__S (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__S (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A0 (.DIODE(net1493));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__S (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__A0 (.DIODE(net1831));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__S (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__S (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__A0 (.DIODE(net1781));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__S (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__A0 (.DIODE(net1813));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__S (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__A0 (.DIODE(net1791));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__S (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__A0 (.DIODE(net1814));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__S (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__A0 (.DIODE(net1811));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__S (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A0 (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__S (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A0 (.DIODE(net1808));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__S (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__A0 (.DIODE(net1806));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__S (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__S (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__A0 (.DIODE(net1809));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__S (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__S (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A0 (.DIODE(net1812));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__S (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A0 (.DIODE(net1807));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__S (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__S (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A0 (.DIODE(net1927));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__S (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A0 (.DIODE(net1941));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__S (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__A0 (.DIODE(net1937));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__S (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__A0 (.DIODE(net1810));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__A1 (.DIODE(\u_s2.u_sync_wbb.u_resp_if.mem[0][27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__S (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A0 (.DIODE(net1930));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__S (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A0 (.DIODE(net1494));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__S (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A0 (.DIODE(net1939));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__S (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A0 (.DIODE(net1943));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A1 (.DIODE(\u_s2.u_sync_wbb.u_resp_if.mem[0][31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__S (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__A (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__B (.DIODE(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__A0 (.DIODE(net1802));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__S (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__A0 (.DIODE(net1805));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__S (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__A0 (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__S (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A0 (.DIODE(net1795));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A1 (.DIODE(\u_s2.u_sync_wbb.u_resp_if.mem[1][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__S (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A0 (.DIODE(net1779));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__S (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A0 (.DIODE(net1796));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__S (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__S (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__A0 (.DIODE(net1493));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__S (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__A0 (.DIODE(net1831));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__S (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__S (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A0 (.DIODE(net1781));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__S (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A0 (.DIODE(net1813));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__S (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__A0 (.DIODE(net1791));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__S (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__A0 (.DIODE(net1814));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__S (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__A0 (.DIODE(net1811));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__S (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__A0 (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__S (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__A0 (.DIODE(net1808));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__S (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A0 (.DIODE(net1806));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__S (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__S (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__A0 (.DIODE(net1809));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__S (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__S (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__A0 (.DIODE(net1812));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__S (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A0 (.DIODE(net1807));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__S (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__S (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A0 (.DIODE(net1927));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__S (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__A0 (.DIODE(net1941));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__S (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__A0 (.DIODE(net1937));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__A1 (.DIODE(\u_s2.u_sync_wbb.u_resp_if.mem[1][26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__S (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__A0 (.DIODE(net1810));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__S (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__A0 (.DIODE(net1930));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__S (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__A0 (.DIODE(net1494));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__S (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__A0 (.DIODE(net1939));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__S (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__A0 (.DIODE(net1943));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__S (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__C_N (.DIODE(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A0 (.DIODE(net1802));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__S (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__A0 (.DIODE(net1805));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__S (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__A0 (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__S (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A0 (.DIODE(net1795));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__S (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A0 (.DIODE(net1779));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__S (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__A0 (.DIODE(net1796));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__S (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__S (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A0 (.DIODE(net1493));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A1 (.DIODE(\u_s2.u_sync_wbb.u_resp_if.mem[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__S (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__A0 (.DIODE(net1831));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__S (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__S (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__A0 (.DIODE(net1781));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__S (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A0 (.DIODE(net1813));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__S (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A0 (.DIODE(net1791));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__S (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A0 (.DIODE(net1814));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__S (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A0 (.DIODE(net1811));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__S (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__A0 (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__S (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A0 (.DIODE(net1808));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__S (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__A0 (.DIODE(net1806));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__S (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__S (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__A0 (.DIODE(net1809));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__A1 (.DIODE(\u_s2.u_sync_wbb.u_resp_if.mem[2][19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__S (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__S (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__A0 (.DIODE(net1812));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__S (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A0 (.DIODE(net1807));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__S (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__S (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__A0 (.DIODE(net1927));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__S (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__A0 (.DIODE(net1941));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__S (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__A0 (.DIODE(net1937));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__S (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A0 (.DIODE(net1810));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__S (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A0 (.DIODE(net1930));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__S (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__A0 (.DIODE(net1494));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__S (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__A0 (.DIODE(net1939));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__S (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__A0 (.DIODE(net1943));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__S (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__A (.DIODE(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__A1 (.DIODE(net1802));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__S (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__A1 (.DIODE(net1805));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__S (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__A1 (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__S (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__A1 (.DIODE(net1795));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__S (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A1 (.DIODE(net1779));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__S (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A1 (.DIODE(net1796));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__S (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__S (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__A1 (.DIODE(net1493));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__S (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__A1 (.DIODE(net1831));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__S (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__S (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A1 (.DIODE(net1781));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__S (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__A1 (.DIODE(net1813));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__S (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A1 (.DIODE(net1791));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__S (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__A1 (.DIODE(net1814));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__S (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__A1 (.DIODE(net1811));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__S (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__A1 (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__S (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__A1 (.DIODE(net1808));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__S (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A1 (.DIODE(net1806));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__S (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__S (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__A1 (.DIODE(net1809));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__S (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__S (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A1 (.DIODE(net1812));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__S (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__A1 (.DIODE(net1807));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__S (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__S (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__A1 (.DIODE(net1927));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__S (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__A1 (.DIODE(net1941));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__S (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__A1 (.DIODE(net1937));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__S (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A1 (.DIODE(net1810));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__S (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A1 (.DIODE(net1930));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__S (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__A1 (.DIODE(net1494));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__S (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__A1 (.DIODE(net1939));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__S (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__A1 (.DIODE(net1943));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__S (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__S0 (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__S1 (.DIODE(net1353));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__A1 (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__S (.DIODE(net1510));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__S0 (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__S1 (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__A1 (.DIODE(_2791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__S (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__S0 (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__S1 (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__S (.DIODE(net1509));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__S0 (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__S1 (.DIODE(net1353));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__A1 (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__S (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__S0 (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__S1 (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__S (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__S0 (.DIODE(net1363));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__S1 (.DIODE(net1356));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__S (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__S0 (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__S1 (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__A1 (.DIODE(_2796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__S (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__S0 (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__S1 (.DIODE(net1353));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__S (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__S0 (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__S1 (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__A1 (.DIODE(_2798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__S (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__A1 (.DIODE(_2374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__S (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__A1 (.DIODE(_2375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__S (.DIODE(net1504));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__S (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__S (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__A1 (.DIODE(_2378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__S (.DIODE(net1504));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__A1 (.DIODE(_2379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__S (.DIODE(net1506));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__S (.DIODE(net1509));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__S (.DIODE(net1509));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__A1 (.DIODE(_2382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__S (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__A1 (.DIODE(_2383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__S (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__S (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__S (.DIODE(net1509));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__A1 (.DIODE(_2386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__S (.DIODE(net1509));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__A1 (.DIODE(_2387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__S (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__S (.DIODE(net1509));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__A1 (.DIODE(_2389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__S (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__S (.DIODE(net1509));
 sky130_fd_sc_hd__diode_2 ANTENNA__5453__S (.DIODE(net1506));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__A1 (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__S (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__S (.DIODE(net1503));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__A1 (.DIODE(_2394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__S (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__A1 (.DIODE(_2395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__S (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__S (.DIODE(net1503));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__A1 (.DIODE(_2397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__S (.DIODE(net1503));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__S (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__A1 (.DIODE(_2399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__S (.DIODE(net1503));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__S (.DIODE(net1503));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__S (.DIODE(net1509));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__A1 (.DIODE(_2402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__S (.DIODE(net1503));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__A1 (.DIODE(_2403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__S (.DIODE(net1506));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__S (.DIODE(net1503));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__S (.DIODE(net1509));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__A1 (.DIODE(_2406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__S (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__S (.DIODE(net1503));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__A1 (.DIODE(_2408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__S (.DIODE(net1506));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__S (.DIODE(net1503));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__A1 (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__S (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__S (.DIODE(net1504));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__S (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__S (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__S (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__A1 (.DIODE(_2414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__S (.DIODE(net1503));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__S (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__S (.DIODE(net1504));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__A (.DIODE(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__S (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__S (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__A1 (.DIODE(_1860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__S (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__A1 (.DIODE(_1856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__S (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__A1 (.DIODE(_1869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__S (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__A1 (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__S (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__A1 (.DIODE(_1867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__S (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__A1 (.DIODE(_1866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__S (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__A1 (.DIODE(_1873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__S (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__A1 (.DIODE(net1240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__A2 (.DIODE(m2_wbd_sel_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__B1 (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__B2 (.DIODE(m3_wbd_sel_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__C1 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__A (.DIODE(m1_wbd_sel_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__B (.DIODE(net1184));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A1 (.DIODE(net1565));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A2 (.DIODE(_1831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__A1 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__S (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__A (.DIODE(net1404));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__B (.DIODE(net1405));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__C (.DIODE(m3_wbd_sel_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__A1 (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__A2 (.DIODE(m2_wbd_sel_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__B1 (.DIODE(m1_wbd_sel_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__B2 (.DIODE(net1183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__C1 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__A1 (.DIODE(m0_wbd_sel_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__A2 (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__A1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__S (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__A (.DIODE(m1_wbd_sel_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__B (.DIODE(_1833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__A1 (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__A2 (.DIODE(m2_wbd_sel_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__B1 (.DIODE(net1185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__B2 (.DIODE(m3_wbd_sel_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__C1 (.DIODE(_1830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__A1 (.DIODE(m0_wbd_sel_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__A2 (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__A1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__S (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A (.DIODE(m1_wbd_sel_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__B (.DIODE(net1183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__A1 (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__A2 (.DIODE(m2_wbd_sel_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__B1 (.DIODE(net1185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__B2 (.DIODE(m3_wbd_sel_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__C1 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__A1 (.DIODE(m0_wbd_sel_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__A2 (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__A1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__S (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__A1 (.DIODE(net1246));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__A2 (.DIODE(net1562));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__B1 (.DIODE(net1240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__A1 (.DIODE(net1246));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__A2 (.DIODE(m2_wbd_dat_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__B1 (.DIODE(net1593));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__B2 (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__A1 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__S (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__A1 (.DIODE(net1246));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__A2 (.DIODE(net1551));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__B1 (.DIODE(net1240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__A1 (.DIODE(net1246));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__A2 (.DIODE(m2_wbd_dat_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__B1 (.DIODE(net1582));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__B2 (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__A1 (.DIODE(_2816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__S (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__A2 (.DIODE(net1543));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__B1 (.DIODE(net1244));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__A2 (.DIODE(m2_wbd_dat_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__B1 (.DIODE(net1574));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__B2 (.DIODE(net1191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__A1 (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__S (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__A1 (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__A2 (.DIODE(m1_wbd_dat_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__B1 (.DIODE(net1240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__A1 (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__A2 (.DIODE(net2088));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__B1 (.DIODE(m0_wbd_dat_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__B2 (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__A1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__S (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A (.DIODE(net1571));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__B (.DIODE(net1191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__A1 (.DIODE(net1244));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__A2 (.DIODE(net1518));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__A1 (.DIODE(net1244));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__A2 (.DIODE(net1540));
 sky130_fd_sc_hd__diode_2 ANTENNA__5522__A1 (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5522__S (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__A1 (.DIODE(net1251));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__A2 (.DIODE(net1539));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__B1 (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__A1 (.DIODE(net1251));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__A2 (.DIODE(net1517));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__B1 (.DIODE(net1570));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__B2 (.DIODE(net1190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__A1 (.DIODE(_2825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__S (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA__5526__A2 (.DIODE(net1538));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__A2 (.DIODE(net1516));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__B1 (.DIODE(net1569));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__B2 (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__S (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__A (.DIODE(net1568));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__B (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__A2 (.DIODE(net1515));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__A2 (.DIODE(net1537));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__A1 (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__S (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__A2 (.DIODE(net1536));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__A2 (.DIODE(net1514));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__B1 (.DIODE(net1567));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__B2 (.DIODE(net1190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__A1 (.DIODE(_2832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__S (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__A (.DIODE(net1566));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__B (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__A2 (.DIODE(net1513));
 sky130_fd_sc_hd__diode_2 ANTENNA__5538__A2 (.DIODE(net1535));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__A1 (.DIODE(_2835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__S (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__A (.DIODE(net1592));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__B (.DIODE(net1190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__A1 (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__A2 (.DIODE(net1534));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__B1 (.DIODE(net1251));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__A1 (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__A2 (.DIODE(net1561));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__A1 (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__S (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__A (.DIODE(net1591));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__B (.DIODE(net1190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__A1 (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__A2 (.DIODE(net1533));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__B1 (.DIODE(net1251));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__A1 (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__A2 (.DIODE(net1560));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__A1 (.DIODE(_2841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__S (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__A (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__B (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__A2 (.DIODE(net1532));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__B1 (.DIODE(net1250));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__A2 (.DIODE(net1559));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__A1 (.DIODE(_2844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__S (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A2 (.DIODE(net1558));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__B1 (.DIODE(net1244));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__A2 (.DIODE(net2066));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__B1 (.DIODE(net1589));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__B2 (.DIODE(net1191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__A1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__S (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__A (.DIODE(net1588));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__B (.DIODE(net1190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__A1 (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__A2 (.DIODE(net1531));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__B1 (.DIODE(net1251));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A1 (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A2 (.DIODE(net1557));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__A1 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__S (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__A2 (.DIODE(net1556));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__B1 (.DIODE(net1244));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__A2 (.DIODE(net1530));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__B1 (.DIODE(net1587));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__B2 (.DIODE(net1191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__A1 (.DIODE(_2851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__S (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__A (.DIODE(net1586));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__B (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__A2 (.DIODE(net1529));
 sky130_fd_sc_hd__diode_2 ANTENNA__5564__A2 (.DIODE(net1555));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__A1 (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__S (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__A1 (.DIODE(net1250));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__A2 (.DIODE(net1554));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__A1 (.DIODE(net1250));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__A2 (.DIODE(net1528));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__B1 (.DIODE(net1585));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__B2 (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5568__A1 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5568__S (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__A1 (.DIODE(net1246));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__A2 (.DIODE(net1553));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__B1 (.DIODE(net1240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__A1 (.DIODE(net1246));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__A2 (.DIODE(net2056));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__B1 (.DIODE(net1584));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__B2 (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__A1 (.DIODE(_2858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__S (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__A (.DIODE(net1583));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__B (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__A2 (.DIODE(net1527));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__B1 (.DIODE(net1250));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__A2 (.DIODE(net1552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__A1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__S (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A1 (.DIODE(net1251));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A2 (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__B1 (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__A2 (.DIODE(net1526));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__B1 (.DIODE(net1581));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__B2 (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__A1 (.DIODE(_2863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__S (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__A2 (.DIODE(net1549));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__B1 (.DIODE(net1244));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__A2 (.DIODE(net1525));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__B1 (.DIODE(net1580));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__B2 (.DIODE(net1191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__S (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__A1 (.DIODE(net1246));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__A2 (.DIODE(net1548));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__B1 (.DIODE(net1244));
 sky130_fd_sc_hd__diode_2 ANTENNA__5583__A1 (.DIODE(net1246));
 sky130_fd_sc_hd__diode_2 ANTENNA__5583__A2 (.DIODE(net2051));
 sky130_fd_sc_hd__diode_2 ANTENNA__5583__B1 (.DIODE(net1579));
 sky130_fd_sc_hd__diode_2 ANTENNA__5583__B2 (.DIODE(net1191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__A1 (.DIODE(_2867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__S (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__A2 (.DIODE(net1547));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__B1 (.DIODE(net1244));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__A2 (.DIODE(net1524));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__B1 (.DIODE(net1578));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__B2 (.DIODE(net1191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__A1 (.DIODE(_2869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__S (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A1 (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A2 (.DIODE(m1_wbd_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__B1 (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__A1 (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__A2 (.DIODE(m2_wbd_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__B1 (.DIODE(m0_wbd_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__B2 (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A1 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__S (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A1 (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A2 (.DIODE(m1_wbd_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__B1 (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A1 (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__B1 (.DIODE(m0_wbd_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__B2 (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A1 (.DIODE(net2080));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__S (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__A2 (.DIODE(net1546));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A2 (.DIODE(net1523));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__B1 (.DIODE(net1577));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__B2 (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A1 (.DIODE(_2875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__S (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__A1 (.DIODE(net1250));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__A2 (.DIODE(net1545));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A1 (.DIODE(net1250));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A2 (.DIODE(net1522));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__B1 (.DIODE(net1576));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__B2 (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__A1 (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__S (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A1 (.DIODE(net1246));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A2 (.DIODE(m1_wbd_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__B1 (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__A1 (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__A2 (.DIODE(m2_wbd_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__B1 (.DIODE(m0_wbd_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__B2 (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__A1 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__S (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__A2 (.DIODE(net1544));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__B1 (.DIODE(net1244));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__A2 (.DIODE(net1521));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__B1 (.DIODE(net1575));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__B2 (.DIODE(net1191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__A1 (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__S (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__A2 (.DIODE(net1542));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__B1 (.DIODE(net1244));
 sky130_fd_sc_hd__diode_2 ANTENNA__5607__A2 (.DIODE(net1520));
 sky130_fd_sc_hd__diode_2 ANTENNA__5607__B1 (.DIODE(net1573));
 sky130_fd_sc_hd__diode_2 ANTENNA__5607__B2 (.DIODE(net1191));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__S (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA__5609__A1 (.DIODE(net1251));
 sky130_fd_sc_hd__diode_2 ANTENNA__5609__A2 (.DIODE(net1541));
 sky130_fd_sc_hd__diode_2 ANTENNA__5609__B1 (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__A1 (.DIODE(net1251));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__A2 (.DIODE(net1519));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__B1 (.DIODE(net1572));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__B2 (.DIODE(net1190));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__A1 (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__S (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__A1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__S (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__A (.DIODE(net1404));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__C (.DIODE(m3_wbd_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__A1 (.DIODE(net1240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__A2 (.DIODE(m2_wbd_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__B1 (.DIODE(m1_wbd_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__B2 (.DIODE(net1183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__C1 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__A1 (.DIODE(net1598));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__A2 (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__A1 (.DIODE(_2888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__S (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__A (.DIODE(\u_s1.gnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__C (.DIODE(m3_wbd_adr_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__A1 (.DIODE(net1240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__A2 (.DIODE(m2_wbd_adr_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__B1 (.DIODE(m1_wbd_adr_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__B2 (.DIODE(net1184));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__C1 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__A1 (.DIODE(net1597));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__A2 (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__A1 (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__S (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A (.DIODE(m1_wbd_adr_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__B (.DIODE(net1183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__A1 (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__A2 (.DIODE(m2_wbd_adr_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__B1 (.DIODE(net1185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__B2 (.DIODE(m3_wbd_adr_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__C1 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__A1 (.DIODE(net1596));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__A2 (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__A1 (.DIODE(_2894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__S (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__A (.DIODE(m1_wbd_adr_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__B (.DIODE(net1184));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__A1 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__A2 (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__B1 (.DIODE(_1832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__B2 (.DIODE(m3_wbd_adr_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__C1 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A1 (.DIODE(net1595));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A2 (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__A1 (.DIODE(_2897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__S (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__A (.DIODE(m1_wbd_adr_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__B (.DIODE(net1183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__A1 (.DIODE(net1240));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__A2 (.DIODE(m2_wbd_adr_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__B1 (.DIODE(net1185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__B2 (.DIODE(m3_wbd_adr_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__C1 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__A1 (.DIODE(net2035));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__A2 (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A1 (.DIODE(_2900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__S (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__A (.DIODE(m1_wbd_adr_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__B (.DIODE(net1184));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__A1 (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__A2 (.DIODE(m2_wbd_adr_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__B1 (.DIODE(net1185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__B2 (.DIODE(m3_wbd_adr_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__C1 (.DIODE(_1830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__A1 (.DIODE(net1594));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__A2 (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__A1 (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__S (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__A (.DIODE(m1_wbd_adr_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__B (.DIODE(net1183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A1 (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A2 (.DIODE(m2_wbd_adr_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__B1 (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__B2 (.DIODE(m3_wbd_adr_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__C1 (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__A1 (.DIODE(net2021));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__A2 (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__A1 (.DIODE(_2906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__S (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__A1 (.DIODE(m2_wbd_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__B1 (.DIODE(net1405));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__A1 (.DIODE(m3_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__A2 (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__A3 (.DIODE(_1853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__A (.DIODE(_1878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__A (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__B (.DIODE(net1183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__C_N (.DIODE(_1879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__A (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__B (.DIODE(_1878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__A1 (.DIODE(m1_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__A2 (.DIODE(_1834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__A3 (.DIODE(_1879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__A1 (.DIODE(m2_wbd_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__B1 (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__A (.DIODE(net1183));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__A1 (.DIODE(m3_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__A2 (.DIODE(_1853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__B (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__A0 (.DIODE(net1405));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__S (.DIODE(_2916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A1 (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A2 (.DIODE(_1878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__A1 (.DIODE(m3_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__A2 (.DIODE(_1853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__A0 (.DIODE(\u_s1.gnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__A1 (.DIODE(_2919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__S (.DIODE(_2916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__B (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__A2 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__A1 (.DIODE(\u_s2.u_sync_wbb.wbm_ack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__B (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__A2 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__B2 (.DIODE(net1400));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__A1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__A2 (.DIODE(_1971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__A3 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__A2 (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__A1 (.DIODE(_1971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__A2 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__B1 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__A0 (.DIODE(\u_s2.u_sync_wbb.m_cmd_wr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__A0 (.DIODE(\u_s2.u_sync_wbb.m_resp_rd_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__A1 (.DIODE(_1982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__S (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__A (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__A (.DIODE(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__A (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__B (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__5677__A (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5677__B (.DIODE(\u_s2.u_sync_wbb.m_cmd_wr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__A (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__C (.DIODE(\u_s2.u_sync_wbb.m_cmd_wr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__A1 (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__A2 (.DIODE(\u_s2.u_sync_wbb.m_cmd_wr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__A (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA__5681__A (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5681__B (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__B (.DIODE(_2571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__C (.DIODE(net1816));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__D (.DIODE(_2573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__D_N (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__A (.DIODE(net1804));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__B (.DIODE(_2575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__C (.DIODE(_2576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__A (.DIODE(\u_s2.u_sync_wbb.s_cmd_rd_data_l[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__C (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__B1 (.DIODE(_1711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__A (.DIODE(net1397));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__B (.DIODE(net1501));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__A1 (.DIODE(net1397));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__A2 (.DIODE(net1501));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__B1 (.DIODE(net1391));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__A (.DIODE(net1390));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__B (.DIODE(net1398));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__C (.DIODE(net1501));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__A (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.rd_ptr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__A (.DIODE(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__S (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__S (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__A1 (.DIODE(_1860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__S (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__A1 (.DIODE(_1856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__S (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A1 (.DIODE(_1869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__S (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__A1 (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__S (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__A1 (.DIODE(_1867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__S (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__A1 (.DIODE(_1866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__S (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__A1 (.DIODE(_1873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__S (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__A1 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__S (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__A1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__S (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__A1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__S (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__A1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__S (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__A1 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__S (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__A1 (.DIODE(_2816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__S (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__A1 (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__S (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__5711__A1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA__5711__S (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__A1 (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__S (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__A1 (.DIODE(_2825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__S (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__S (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__A1 (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__S (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__A1 (.DIODE(_2832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__S (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A1 (.DIODE(_2835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__S (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__A1 (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__S (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__A1 (.DIODE(_2841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__S (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__A1 (.DIODE(_2844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__S (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__A1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__S (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__A1 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__S (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__A1 (.DIODE(_2851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__S (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__A1 (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__S (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__A1 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__S (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__A1 (.DIODE(_2858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__S (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__A1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__S (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__A1 (.DIODE(_2863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__S (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__S (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__A1 (.DIODE(_2867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__S (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__A1 (.DIODE(_2869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__S (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__A1 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__S (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__A1 (.DIODE(net2080));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__S (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__A1 (.DIODE(_2875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__S (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__A1 (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__S (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__A1 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__S (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA__5737__A1 (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5737__S (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__S (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__A1 (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__S (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__A1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__S (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__A1 (.DIODE(_2888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__S (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__A1 (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__S (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__A1 (.DIODE(_2894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__S (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__A1 (.DIODE(_2897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__S (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__5745__A1 (.DIODE(_2900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5745__S (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A1 (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__S (.DIODE(_2944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__A1 (.DIODE(_2906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__S (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__A (.DIODE(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__B (.DIODE(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__C_N (.DIODE(\u_s0.u_sync_wbb.m_cmd_wr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__A0 (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__S (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__A0 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__S (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__A0 (.DIODE(_1792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__S (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__A0 (.DIODE(_1794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__S (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__A0 (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__S (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__A0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__S (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__A0 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__S (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A0 (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__S (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__A0 (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__S (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__A0 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__S (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__A (.DIODE(net1371));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__B (.DIODE(net1375));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__C (.DIODE(m3_wbd_sel_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__A1 (.DIODE(net1259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__A2 (.DIODE(net2082));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__B1 (.DIODE(net2085));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__B2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__C1 (.DIODE(net1205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__A1 (.DIODE(net1565));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__A2 (.DIODE(net1199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__A0 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__S (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__A1 (.DIODE(net1259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__A2 (.DIODE(m2_wbd_sel_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__B1 (.DIODE(net1208));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__B2 (.DIODE(m3_wbd_sel_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__C1 (.DIODE(net1204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__A1 (.DIODE(m1_wbd_sel_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__A2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__B1 (.DIODE(_2949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__A1 (.DIODE(net2030));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__A2 (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__S (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__A1 (.DIODE(net1259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__A2 (.DIODE(m2_wbd_sel_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__B1 (.DIODE(net1206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__B2 (.DIODE(m3_wbd_sel_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__C1 (.DIODE(net1205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__A1 (.DIODE(m1_wbd_sel_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__A2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__B1 (.DIODE(_2952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__A0 (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__S (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__A1 (.DIODE(net1259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__A2 (.DIODE(m2_wbd_sel_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__B1 (.DIODE(net1206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__B2 (.DIODE(m3_wbd_sel_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__C1 (.DIODE(net1205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__A1 (.DIODE(m1_wbd_sel_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__A2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__B1 (.DIODE(_2955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__A2 (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__A0 (.DIODE(_2957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__S (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__A (.DIODE(net1593));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__B (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__A1 (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__A2 (.DIODE(m2_wbd_dat_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A1 (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A2 (.DIODE(net1562));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__S (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A1 (.DIODE(net1273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A2 (.DIODE(net1551));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__B1 (.DIODE(net1263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A1 (.DIODE(net1273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A2 (.DIODE(m2_wbd_dat_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__B1 (.DIODE(net1582));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__B2 (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A0 (.DIODE(_2962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__S (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__A2 (.DIODE(net1543));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__B1 (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__A1 (.DIODE(net1273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__A2 (.DIODE(m2_wbd_dat_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__B1 (.DIODE(net1574));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__B2 (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A0 (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__S (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__A1 (.DIODE(net1270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__A2 (.DIODE(m1_wbd_dat_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__B1 (.DIODE(net1261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__A1 (.DIODE(net1270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__A2 (.DIODE(net2088));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__B1 (.DIODE(m0_wbd_dat_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__B2 (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__A0 (.DIODE(_2966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__S (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__A (.DIODE(m0_wbd_dat_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__B (.DIODE(net1199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__A1 (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__A2 (.DIODE(m2_wbd_dat_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__B1 (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A1 (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A2 (.DIODE(net2006));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__S (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__A1 (.DIODE(net1273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__A2 (.DIODE(net1539));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__B1 (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__A1 (.DIODE(net1273));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__A2 (.DIODE(net1517));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__B1 (.DIODE(net1570));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__B2 (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__S (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A1 (.DIODE(net1270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A2 (.DIODE(net1538));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__B1 (.DIODE(net1261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__A1 (.DIODE(net1270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__A2 (.DIODE(net1516));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__B1 (.DIODE(net1569));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__B2 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__S (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__A (.DIODE(m0_wbd_dat_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__B (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__A2 (.DIODE(m2_wbd_dat_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__A2 (.DIODE(net2084));
 sky130_fd_sc_hd__diode_2 ANTENNA__5801__A0 (.DIODE(_2976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5801__S (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__A (.DIODE(m0_wbd_dat_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__B (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__A1 (.DIODE(net1261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__A2 (.DIODE(m2_wbd_dat_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__B1 (.DIODE(net1270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__A1 (.DIODE(net1261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__A2 (.DIODE(net2077));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__S (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__A2 (.DIODE(net1535));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__B1 (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__A2 (.DIODE(net1513));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__B1 (.DIODE(net1566));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__B2 (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__S (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__A2 (.DIODE(net1561));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__B1 (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__A2 (.DIODE(net1534));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__B1 (.DIODE(net1592));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__B2 (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__S (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__A2 (.DIODE(net1560));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__B1 (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__A2 (.DIODE(net1533));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__B1 (.DIODE(net1591));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__B2 (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5814__S (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__A (.DIODE(m0_wbd_dat_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__B (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__A2 (.DIODE(m2_wbd_dat_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__B1 (.DIODE(net1267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__A2 (.DIODE(net2055));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__A0 (.DIODE(_2988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__S (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__A (.DIODE(net1589));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__B (.DIODE(net1198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__A2 (.DIODE(m2_wbd_dat_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__A2 (.DIODE(net1558));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__A0 (.DIODE(_2991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__S (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__A2 (.DIODE(net1557));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__B1 (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__A2 (.DIODE(net1531));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__B1 (.DIODE(net1588));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__B2 (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__S (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__A2 (.DIODE(net1556));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__B1 (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__A2 (.DIODE(net2036));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__B1 (.DIODE(net1587));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__B2 (.DIODE(net1199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__S (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__A (.DIODE(m0_wbd_dat_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__B (.DIODE(net1199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__A2 (.DIODE(m2_wbd_dat_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A2 (.DIODE(net2039));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__A0 (.DIODE(_2998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__S (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A (.DIODE(net1585));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__B (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__A1 (.DIODE(net1261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__A2 (.DIODE(net1528));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__B1 (.DIODE(net1270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__A1 (.DIODE(net1261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__A2 (.DIODE(net1554));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A0 (.DIODE(_3001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__S (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__A (.DIODE(net1584));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__B (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__A2 (.DIODE(m2_wbd_dat_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__A2 (.DIODE(net1553));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__C1 (.DIODE(_3003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__A0 (.DIODE(_3004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__S (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA__5841__A (.DIODE(net1583));
 sky130_fd_sc_hd__diode_2 ANTENNA__5841__B (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__A1 (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__A2 (.DIODE(m2_wbd_dat_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__B1 (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__A1 (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__A2 (.DIODE(net2008));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__S (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__A (.DIODE(m0_wbd_dat_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__B (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5846__A2 (.DIODE(m2_wbd_dat_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__A2 (.DIODE(net2064));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__A0 (.DIODE(_3010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__S (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__A1 (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__A2 (.DIODE(net1549));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__B1 (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__A1 (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__A2 (.DIODE(net1525));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__B1 (.DIODE(net1580));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__B2 (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__A0 (.DIODE(_3012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__S (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__A2 (.DIODE(net1548));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__A2 (.DIODE(net2051));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__B1 (.DIODE(net1579));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__B2 (.DIODE(net1198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__A0 (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__S (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__A1 (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__A2 (.DIODE(net1547));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__B1 (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A1 (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A2 (.DIODE(net1524));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__B1 (.DIODE(net1578));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__B2 (.DIODE(net1199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__A0 (.DIODE(_3016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__S (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__A (.DIODE(m0_wbd_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__B (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__A2 (.DIODE(m2_wbd_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__A2 (.DIODE(net2016));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__S (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__A (.DIODE(m0_wbd_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__B (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__A1 (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__A2 (.DIODE(m2_wbd_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__B1 (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__A1 (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__A2 (.DIODE(net2037));
 sky130_fd_sc_hd__diode_2 ANTENNA__5865__S (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__A2 (.DIODE(m1_wbd_dat_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__A2 (.DIODE(net2067));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__B1 (.DIODE(net2018));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__B2 (.DIODE(net1198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A0 (.DIODE(_3024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__S (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A1 (.DIODE(net1267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A2 (.DIODE(net2043));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__A1 (.DIODE(net1267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__A2 (.DIODE(net2041));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__B1 (.DIODE(net2010));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__B2 (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5871__S (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__A (.DIODE(m0_wbd_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__B (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5873__A2 (.DIODE(m2_wbd_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5873__B1 (.DIODE(net1267));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__A2 (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__A0 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__S (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__A2 (.DIODE(m1_wbd_dat_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5877__B1 (.DIODE(net1575));
 sky130_fd_sc_hd__diode_2 ANTENNA__5877__B2 (.DIODE(net1199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__A0 (.DIODE(_3031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__S (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA__5879__A1 (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5879__A2 (.DIODE(net1542));
 sky130_fd_sc_hd__diode_2 ANTENNA__5879__B1 (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A1 (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A2 (.DIODE(net1520));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__B1 (.DIODE(net1573));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__B2 (.DIODE(net1199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5881__S (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__A1 (.DIODE(net1268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__A2 (.DIODE(m1_wbd_dat_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__B1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5883__A1 (.DIODE(net1268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5883__A2 (.DIODE(m2_wbd_dat_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5883__B2 (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__S (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__A0 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__S (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__A (.DIODE(net1371));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__B (.DIODE(net1375));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__C (.DIODE(m3_wbd_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__A1 (.DIODE(net1258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__A2 (.DIODE(m2_wbd_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__B1 (.DIODE(m1_wbd_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__B2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__C1 (.DIODE(net1204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__A1 (.DIODE(net1598));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__A2 (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__B1 (.DIODE(_3036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5889__S (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__A (.DIODE(net1271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__B (.DIODE(net1375));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__C (.DIODE(m1_wbd_adr_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__A1 (.DIODE(net1263));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__A2 (.DIODE(m2_wbd_adr_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__B1 (.DIODE(net1208));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__B2 (.DIODE(m3_wbd_adr_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__C1 (.DIODE(net1205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__A1 (.DIODE(net1597));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__A2 (.DIODE(net1199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5893__A0 (.DIODE(_3041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5893__S (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__A (.DIODE(net1271));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__B (.DIODE(net1375));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__C (.DIODE(m1_wbd_adr_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__A1 (.DIODE(net1259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__A2 (.DIODE(m2_wbd_adr_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__B1 (.DIODE(net1208));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__B2 (.DIODE(m3_wbd_adr_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__C1 (.DIODE(net1204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5896__A1 (.DIODE(net1596));
 sky130_fd_sc_hd__diode_2 ANTENNA__5896__A2 (.DIODE(net1199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__A0 (.DIODE(_3044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__S (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__A (.DIODE(net1270));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__B (.DIODE(net1375));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__C (.DIODE(m1_wbd_adr_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__A1 (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__A2 (.DIODE(m2_wbd_adr_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__B2 (.DIODE(m3_wbd_adr_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__C1 (.DIODE(net1205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__A1 (.DIODE(net1595));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__A2 (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__A0 (.DIODE(_3047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__S (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__A1 (.DIODE(net1259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__A2 (.DIODE(m2_wbd_adr_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__B1 (.DIODE(net1208));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__B2 (.DIODE(m3_wbd_adr_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__C1 (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__A1 (.DIODE(net1983));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__A2 (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__B1 (.DIODE(_3048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__A1 (.DIODE(net1832));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__A2 (.DIODE(net1198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__A0 (.DIODE(_3050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__S (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__A1 (.DIODE(net1261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__A2 (.DIODE(m2_wbd_adr_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__B1 (.DIODE(net1208));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__B2 (.DIODE(m3_wbd_adr_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__C1 (.DIODE(net1205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__A1 (.DIODE(m1_wbd_adr_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__A2 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__B1 (.DIODE(_3051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5908__A1 (.DIODE(net1594));
 sky130_fd_sc_hd__diode_2 ANTENNA__5908__A2 (.DIODE(net1194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__A0 (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__S (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__A (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__B (.DIODE(net1375));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__C (.DIODE(m1_wbd_adr_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__A1 (.DIODE(net1261));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__A2 (.DIODE(m2_wbd_adr_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__B1 (.DIODE(net1208));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__B2 (.DIODE(m3_wbd_adr_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__C1 (.DIODE(net1205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__A1 (.DIODE(net2021));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__A2 (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5913__S (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__A (.DIODE(net1268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__B (.DIODE(net1374));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__C (.DIODE(m1_wbd_adr_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__A1 (.DIODE(net1258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__A2 (.DIODE(m2_wbd_adr_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__B1 (.DIODE(net1206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__B2 (.DIODE(m3_wbd_adr_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__C1 (.DIODE(net1204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A1 (.DIODE(net2031));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A2 (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__S (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__A (.DIODE(net1370));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__B (.DIODE(net1374));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__C (.DIODE(m3_wbd_adr_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__A1 (.DIODE(net1258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__A2 (.DIODE(m2_wbd_adr_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__B1 (.DIODE(m1_wbd_adr_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__B2 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__C1 (.DIODE(net1204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__A1 (.DIODE(m0_wbd_adr_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__A2 (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__S (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__A1 (.DIODE(net1264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__A2 (.DIODE(m2_wbd_adr_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__B1 (.DIODE(net1254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__A1 (.DIODE(net1264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__A2 (.DIODE(m1_wbd_adr_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__B1 (.DIODE(net1206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__B2 (.DIODE(m3_wbd_adr_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5924__A1 (.DIODE(m0_wbd_adr_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5924__A2 (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA__5925__S (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__A1 (.DIODE(net1264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__A2 (.DIODE(m2_wbd_adr_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__B1 (.DIODE(net1254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__A1 (.DIODE(net1264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__A2 (.DIODE(m1_wbd_adr_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__B1 (.DIODE(net1206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__B2 (.DIODE(m3_wbd_adr_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__A1 (.DIODE(m0_wbd_adr_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__A2 (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__A0 (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__S (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__A1 (.DIODE(net1264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__A2 (.DIODE(m2_wbd_adr_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__B1 (.DIODE(net1258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__A1 (.DIODE(net1268));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__A2 (.DIODE(m1_wbd_adr_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__B1 (.DIODE(net1206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__B2 (.DIODE(m3_wbd_adr_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__A1 (.DIODE(net1908));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__A2 (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__S (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__A1 (.DIODE(net1264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__A2 (.DIODE(net1997));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A1 (.DIODE(net1264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A2 (.DIODE(m1_wbd_adr_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__B1 (.DIODE(net1206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__B2 (.DIODE(m3_wbd_adr_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__A2 (.DIODE(net1194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__B1 (.DIODE(_3072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__B2 (.DIODE(_3073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__S (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__A1 (.DIODE(net1264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__A2 (.DIODE(m2_wbd_adr_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__B1 (.DIODE(net1254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__A1 (.DIODE(net1264));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__A2 (.DIODE(m1_wbd_adr_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__B1 (.DIODE(net1206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__B2 (.DIODE(m3_wbd_adr_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__B2 (.DIODE(_3076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__S (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__A1 (.DIODE(net1258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__A2 (.DIODE(m2_wbd_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__B1 (.DIODE(net1209));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__B2 (.DIODE(m3_wbd_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__C1 (.DIODE(net1204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5943__A1 (.DIODE(m1_wbd_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5943__A2 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__5943__B1 (.DIODE(_3078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__A2 (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__B1 (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__A0 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__S (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__A1 (.DIODE(net1259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__A2 (.DIODE(m2_wbd_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__B1 (.DIODE(net1209));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__B2 (.DIODE(m3_wbd_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__C1 (.DIODE(net1204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__A1 (.DIODE(m1_wbd_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__A2 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__B1 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__A2 (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5949__A0 (.DIODE(_3083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5949__S (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__C (.DIODE(m3_wbd_adr_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5951__A2 (.DIODE(m2_wbd_adr_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__A2 (.DIODE(net1194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__B1 (.DIODE(_3084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__S (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__A1 (.DIODE(net1259));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__A2 (.DIODE(m2_wbd_adr_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__B1 (.DIODE(net1206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__B2 (.DIODE(m3_wbd_adr_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__C1 (.DIODE(net1205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__B1 (.DIODE(_3087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__A2 (.DIODE(net1194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__B1 (.DIODE(_3088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__S (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__C (.DIODE(m3_wbd_adr_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__A2 (.DIODE(m2_wbd_adr_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__B1 (.DIODE(m1_wbd_adr_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__A2 (.DIODE(net1194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__B1 (.DIODE(_3090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__A0 (.DIODE(_3092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__S (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__C (.DIODE(m3_wbd_adr_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5963__A2 (.DIODE(m2_wbd_adr_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5963__B2 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__5964__B1 (.DIODE(_3093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5965__A0 (.DIODE(_3095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5965__S (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA__5966__C (.DIODE(m3_wbd_adr_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A1 (.DIODE(net1254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A2 (.DIODE(m2_wbd_adr_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__B1 (.DIODE(m1_wbd_adr_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__B2 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__C1 (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__A2 (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__B2 (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__A0 (.DIODE(_3098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__S (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__C (.DIODE(m3_wbd_adr_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__A2 (.DIODE(m2_wbd_adr_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__A2 (.DIODE(net1194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__B1 (.DIODE(_3099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__S (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__C (.DIODE(m3_wbd_adr_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__A2 (.DIODE(m2_wbd_adr_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__B1 (.DIODE(m1_wbd_adr_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__B2 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__B1 (.DIODE(_3102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__B2 (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__S (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__C (.DIODE(m3_wbd_adr_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__A1 (.DIODE(net1254));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__A2 (.DIODE(m2_wbd_adr_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__B1 (.DIODE(m1_wbd_adr_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__B2 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__5980__A2 (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA__5980__B1 (.DIODE(_3105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5980__B2 (.DIODE(_3106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__S (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA__5982__A (.DIODE(net1370));
 sky130_fd_sc_hd__diode_2 ANTENNA__5982__C (.DIODE(m3_wbd_adr_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5983__A2 (.DIODE(m2_wbd_adr_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5983__B2 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__B1 (.DIODE(_3108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__B2 (.DIODE(_3109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5985__S (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__C (.DIODE(m3_wbd_adr_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__A2 (.DIODE(m2_wbd_adr_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__B1 (.DIODE(m1_wbd_adr_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5988__A2 (.DIODE(net1194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5988__B1 (.DIODE(_3111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5988__B2 (.DIODE(_3112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__S (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__A1 (.DIODE(net1258));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__A2 (.DIODE(m2_wbd_adr_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__B1 (.DIODE(net1209));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__B2 (.DIODE(m3_wbd_adr_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__C1 (.DIODE(net1204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__A1 (.DIODE(m1_wbd_adr_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__B1 (.DIODE(_3114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5992__A2 (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5992__B1 (.DIODE(_3115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__S (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA__5994__A (.DIODE(net1370));
 sky130_fd_sc_hd__diode_2 ANTENNA__5994__B (.DIODE(net1374));
 sky130_fd_sc_hd__diode_2 ANTENNA__5994__C (.DIODE(m3_wbd_adr_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__A2 (.DIODE(m2_wbd_adr_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__B1 (.DIODE(m1_wbd_adr_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__A2 (.DIODE(net1194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__B1 (.DIODE(_3117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__B2 (.DIODE(_3118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__S (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA__5998__A (.DIODE(net1370));
 sky130_fd_sc_hd__diode_2 ANTENNA__5998__B (.DIODE(net1374));
 sky130_fd_sc_hd__diode_2 ANTENNA__5998__C (.DIODE(m3_wbd_adr_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__A2 (.DIODE(m2_wbd_adr_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6000__A2 (.DIODE(net1194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6000__B1 (.DIODE(_3120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6001__S (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA__6002__A1 (.DIODE(net1258));
 sky130_fd_sc_hd__diode_2 ANTENNA__6002__A2 (.DIODE(m2_wbd_adr_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6002__B1 (.DIODE(net1206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6002__B2 (.DIODE(m3_wbd_adr_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6002__C1 (.DIODE(net1204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__A1 (.DIODE(m1_wbd_adr_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__B1 (.DIODE(_3123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6004__A2 (.DIODE(net1194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6005__S (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA__6006__A (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__6006__B (.DIODE(\u_s2.u_sync_wbb.m_resp_rd_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__A1 (.DIODE(net1384));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__A2 (.DIODE(\u_s2.u_sync_wbb.m_resp_rd_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__B1 (.DIODE(\u_s2.u_sync_wbb.u_resp_if.rd_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__A (.DIODE(net1379));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__B (.DIODE(net1384));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__C (.DIODE(\u_s2.u_sync_wbb.m_resp_rd_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6011__A (.DIODE(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6011__C (.DIODE(_2423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__S (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__A0 (.DIODE(net1902));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__S (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__A0 (.DIODE(net2060));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__S (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__A0 (.DIODE(net1903));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__S (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__A0 (.DIODE(net2063));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__S (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__6017__A0 (.DIODE(net2065));
 sky130_fd_sc_hd__diode_2 ANTENNA__6017__S (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__A0 (.DIODE(net1880));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__S (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__A0 (.DIODE(net1886));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__S (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__A0 (.DIODE(net1904));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__S (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__6021__A0 (.DIODE(net1892));
 sky130_fd_sc_hd__diode_2 ANTENNA__6021__S (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__A0 (.DIODE(net1898));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__S (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__6023__S (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__S (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__S (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__6026__S (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__6027__A0 (.DIODE(net1881));
 sky130_fd_sc_hd__diode_2 ANTENNA__6027__S (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__A0 (.DIODE(net1851));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__S (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__6029__A0 (.DIODE(net1879));
 sky130_fd_sc_hd__diode_2 ANTENNA__6029__S (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__A0 (.DIODE(net1889));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__S (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__A0 (.DIODE(net1993));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__S (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__S (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__A0 (.DIODE(net1912));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__S (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__S (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__6035__S (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__A0 (.DIODE(net1893));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__S (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__6037__S (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__S (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__S (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__S (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__A0 (.DIODE(net1845));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__S (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__S (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__A0 (.DIODE(net1899));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__S (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__B (.DIODE(_2423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__C_N (.DIODE(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__S (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__A0 (.DIODE(net1902));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__A0 (.DIODE(net1882));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__S (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__6048__A0 (.DIODE(net1903));
 sky130_fd_sc_hd__diode_2 ANTENNA__6048__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__A0 (.DIODE(net2063));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__S (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__A0 (.DIODE(net2065));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__S (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__A0 (.DIODE(net1880));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__S (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__A0 (.DIODE(net1886));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__S (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__A0 (.DIODE(net1904));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__A0 (.DIODE(net1892));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__S (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__A0 (.DIODE(net1898));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__S (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__S (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__6058__A0 (.DIODE(net2003));
 sky130_fd_sc_hd__diode_2 ANTENNA__6058__S (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__S (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__6060__A0 (.DIODE(net1881));
 sky130_fd_sc_hd__diode_2 ANTENNA__6060__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__A0 (.DIODE(net1851));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__S (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__6062__A0 (.DIODE(net1879));
 sky130_fd_sc_hd__diode_2 ANTENNA__6062__S (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__A0 (.DIODE(net1889));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__S (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__A0 (.DIODE(net1993));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__S (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__6066__A0 (.DIODE(net1912));
 sky130_fd_sc_hd__diode_2 ANTENNA__6066__S (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__S (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__S (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__A0 (.DIODE(net1893));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__A0 (.DIODE(net1907));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__A0 (.DIODE(net1891));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__S (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__S (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__A0 (.DIODE(net1845));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__S (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__6075__S (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__6076__A0 (.DIODE(net1899));
 sky130_fd_sc_hd__diode_2 ANTENNA__6076__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__A (.DIODE(_2423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__B (.DIODE(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__S (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__A0 (.DIODE(net1902));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__S (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__A0 (.DIODE(net1882));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__S (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__A0 (.DIODE(net1903));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__S (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__A0 (.DIODE(net1890));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__S (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__A0 (.DIODE(net2065));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__S (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__A0 (.DIODE(net1880));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__S (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__A0 (.DIODE(net1886));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__S (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__A0 (.DIODE(net1904));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__S (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__A0 (.DIODE(net1892));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__S (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__A0 (.DIODE(net1898));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__S (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__S (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__S (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__A0 (.DIODE(net2003));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__S (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__S (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__A0 (.DIODE(net1881));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__S (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A0 (.DIODE(net1851));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__S (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__6095__A0 (.DIODE(net1879));
 sky130_fd_sc_hd__diode_2 ANTENNA__6095__S (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__A0 (.DIODE(net1889));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__S (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__A0 (.DIODE(net1993));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__S (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__S (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__A0 (.DIODE(net1912));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__S (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__S (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__S (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__6102__A0 (.DIODE(net1893));
 sky130_fd_sc_hd__diode_2 ANTENNA__6102__S (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__6103__A0 (.DIODE(net1907));
 sky130_fd_sc_hd__diode_2 ANTENNA__6103__S (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__A0 (.DIODE(net1891));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__S (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__S (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__S (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__A0 (.DIODE(net1845));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__S (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__S (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__A0 (.DIODE(net1899));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__S (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__A (.DIODE(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__S (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__A1 (.DIODE(net1902));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__S (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__A1 (.DIODE(net1882));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__S (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__A1 (.DIODE(net1903));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__S (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__A1 (.DIODE(net2063));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__S (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__A1 (.DIODE(net2065));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__S (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__6117__A1 (.DIODE(net1880));
 sky130_fd_sc_hd__diode_2 ANTENNA__6117__S (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__A1 (.DIODE(net1886));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__S (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__A1 (.DIODE(net1904));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__S (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__A1 (.DIODE(net1892));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__S (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__A1 (.DIODE(net1999));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__S (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__6122__S (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__S (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__6124__A1 (.DIODE(net2003));
 sky130_fd_sc_hd__diode_2 ANTENNA__6124__S (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__6125__S (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__A1 (.DIODE(net1881));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__S (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__A1 (.DIODE(net1851));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__S (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__A1 (.DIODE(net1879));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__S (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__A1 (.DIODE(net1889));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__S (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__A1 (.DIODE(net1993));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__S (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__S (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__A1 (.DIODE(net1912));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__S (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__6133__S (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__6134__S (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__6135__A1 (.DIODE(net1893));
 sky130_fd_sc_hd__diode_2 ANTENNA__6135__S (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__A1 (.DIODE(net1907));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__S (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__A1 (.DIODE(net1891));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__S (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__S (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__S (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__A1 (.DIODE(net1845));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__S (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__6141__S (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__A1 (.DIODE(net1899));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__S (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__S (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA__6144__A1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__6144__S (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__S (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__A1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__S (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__A1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__S (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__A1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__S (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__S (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__A1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__S (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__A1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__S (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__A (.DIODE(m1_wbd_sel_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__A1 (.DIODE(net1238));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__A2 (.DIODE(net2082));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__B1 (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__B2 (.DIODE(m3_wbd_sel_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__C1 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6154__A1 (.DIODE(net1565));
 sky130_fd_sc_hd__diode_2 ANTENNA__6154__A2 (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__A1 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__S (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA__6156__A (.DIODE(net1410));
 sky130_fd_sc_hd__diode_2 ANTENNA__6156__B (.DIODE(net1408));
 sky130_fd_sc_hd__diode_2 ANTENNA__6156__C (.DIODE(m3_wbd_sel_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6157__A1 (.DIODE(net1233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6157__A2 (.DIODE(m2_wbd_sel_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6157__B1 (.DIODE(m1_wbd_sel_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6157__B2 (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6157__C1 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__A1 (.DIODE(net1915));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__A2 (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__A1 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__S (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__A (.DIODE(net1410));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__B (.DIODE(net1408));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__C (.DIODE(m3_wbd_sel_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6161__A1 (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6161__A2 (.DIODE(m2_wbd_sel_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6161__B1 (.DIODE(m1_wbd_sel_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6161__B2 (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6161__C1 (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__A1 (.DIODE(net1974));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__A2 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__A1 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__S (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__A (.DIODE(net1410));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__B (.DIODE(net1407));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__C (.DIODE(m3_wbd_sel_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__A1 (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__B1 (.DIODE(net2059));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__B2 (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__C1 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__A1 (.DIODE(net1970));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__A2 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__A1 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__S (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__A1 (.DIODE(net1225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__A2 (.DIODE(net1562));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__B1 (.DIODE(net1233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__A1 (.DIODE(net1225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__A2 (.DIODE(net2050));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__B1 (.DIODE(net1593));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__B2 (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6170__A1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__6170__S (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__A1 (.DIODE(net1225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__A2 (.DIODE(net1551));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__B1 (.DIODE(net1233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__A1 (.DIODE(net1225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__A2 (.DIODE(net2078));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__B1 (.DIODE(net1582));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__B2 (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6173__A1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__6173__S (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__A (.DIODE(net1574));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__B (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__A2 (.DIODE(net1543));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__B1 (.DIODE(net1237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__A2 (.DIODE(net1855));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__A1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__S (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__A (.DIODE(m0_wbd_dat_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__B (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6179__A1 (.DIODE(net1224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6179__A2 (.DIODE(m1_wbd_dat_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6179__B1 (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__A1 (.DIODE(net1224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__A2 (.DIODE(net2088));
 sky130_fd_sc_hd__diode_2 ANTENNA__6181__A1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__6181__S (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA__6182__A1 (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6182__A2 (.DIODE(net1540));
 sky130_fd_sc_hd__diode_2 ANTENNA__6182__B1 (.DIODE(net1237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__A1 (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__A2 (.DIODE(net1518));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__B1 (.DIODE(net1571));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__B2 (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__A1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__S (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA__6185__A2 (.DIODE(net1539));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__A2 (.DIODE(net1517));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__B1 (.DIODE(net1570));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__B2 (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__A1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__S (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__A (.DIODE(net1569));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__B (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6189__A1 (.DIODE(net1235));
 sky130_fd_sc_hd__diode_2 ANTENNA__6189__A2 (.DIODE(net1516));
 sky130_fd_sc_hd__diode_2 ANTENNA__6189__B1 (.DIODE(net1230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__A1 (.DIODE(net1235));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__A2 (.DIODE(net1538));
 sky130_fd_sc_hd__diode_2 ANTENNA__6191__A1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__6191__S (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA__6192__A1 (.DIODE(net1230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6192__A2 (.DIODE(net1537));
 sky130_fd_sc_hd__diode_2 ANTENNA__6192__B1 (.DIODE(net1235));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__A1 (.DIODE(net1230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__A2 (.DIODE(net1515));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__B1 (.DIODE(net1568));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__B2 (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__A1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__S (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__A2 (.DIODE(net1536));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__A2 (.DIODE(net1514));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__B1 (.DIODE(net1567));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__B2 (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__A1 (.DIODE(_3164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__S (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__A (.DIODE(net1566));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__B (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__A2 (.DIODE(net1535));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__A2 (.DIODE(net1513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__A1 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__S (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA__6202__A (.DIODE(net1592));
 sky130_fd_sc_hd__diode_2 ANTENNA__6202__B (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__A2 (.DIODE(net1534));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__A2 (.DIODE(net1561));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__A0 (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.mem[3][28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__A1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__S (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__A2 (.DIODE(net1560));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__A2 (.DIODE(net1533));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__B1 (.DIODE(net1591));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__B2 (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__A1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__S (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__A1 (.DIODE(net1230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__A2 (.DIODE(net1559));
 sky130_fd_sc_hd__diode_2 ANTENNA__6210__A1 (.DIODE(net1230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6210__A2 (.DIODE(net1532));
 sky130_fd_sc_hd__diode_2 ANTENNA__6210__B1 (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__6210__B2 (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6211__A1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__6211__S (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__A1 (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__A2 (.DIODE(net1558));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__B1 (.DIODE(net1237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A1 (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A2 (.DIODE(net2066));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__B1 (.DIODE(net1589));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__B2 (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__A1 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__S (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__A (.DIODE(net1588));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__B (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6216__A2 (.DIODE(net1557));
 sky130_fd_sc_hd__diode_2 ANTENNA__6217__A2 (.DIODE(net1531));
 sky130_fd_sc_hd__diode_2 ANTENNA__6218__A1 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA__6218__S (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__A (.DIODE(net1587));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__B (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6220__A2 (.DIODE(net1556));
 sky130_fd_sc_hd__diode_2 ANTENNA__6220__B1 (.DIODE(net1237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__A2 (.DIODE(net1530));
 sky130_fd_sc_hd__diode_2 ANTENNA__6222__A1 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA__6222__S (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__A (.DIODE(net1586));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__B (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__A2 (.DIODE(net1529));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__A2 (.DIODE(net1555));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__A1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__S (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA__6227__A (.DIODE(net1585));
 sky130_fd_sc_hd__diode_2 ANTENNA__6227__B (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6228__A2 (.DIODE(net1528));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__A2 (.DIODE(net1554));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__A1 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__S (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__A (.DIODE(net1584));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__B (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__A1 (.DIODE(net1225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__A2 (.DIODE(net1553));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__B1 (.DIODE(net1233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__A1 (.DIODE(net1225));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__A2 (.DIODE(net1928));
 sky130_fd_sc_hd__diode_2 ANTENNA__6234__A1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__6234__S (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__A2 (.DIODE(net1552));
 sky130_fd_sc_hd__diode_2 ANTENNA__6236__A2 (.DIODE(net1527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6236__B1 (.DIODE(net1583));
 sky130_fd_sc_hd__diode_2 ANTENNA__6236__B2 (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6237__A1 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__6237__S (.DIODE(_2934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6238__A1 (.DIODE(net1230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6238__A2 (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__6238__B1 (.DIODE(net1235));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__A1 (.DIODE(net1230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__A2 (.DIODE(net1526));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__B1 (.DIODE(net1581));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__B2 (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__A1 (.DIODE(_3195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__S (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__A1 (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__A2 (.DIODE(net1549));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__B1 (.DIODE(net1237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__A1 (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__A2 (.DIODE(net1525));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__B1 (.DIODE(net1580));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__B2 (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__A1 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__S (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA__6244__A (.DIODE(net1579));
 sky130_fd_sc_hd__diode_2 ANTENNA__6244__B (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__A1 (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__A2 (.DIODE(net1548));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__B1 (.DIODE(net1237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__A1 (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__A2 (.DIODE(net2051));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__A1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__S (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__A1 (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__A2 (.DIODE(net1547));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__B1 (.DIODE(net1237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6249__A1 (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA__6249__A2 (.DIODE(net1524));
 sky130_fd_sc_hd__diode_2 ANTENNA__6249__B1 (.DIODE(net1578));
 sky130_fd_sc_hd__diode_2 ANTENNA__6249__B2 (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6250__A1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__6250__S (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__A1 (.DIODE(net1224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__A2 (.DIODE(m1_wbd_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__B1 (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__A1 (.DIODE(net1224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__B1 (.DIODE(m0_wbd_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__B2 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6253__A1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__6253__S (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__A1 (.DIODE(net1224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__A2 (.DIODE(m1_wbd_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__B1 (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__A1 (.DIODE(net1224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__B1 (.DIODE(m0_wbd_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__B2 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6256__A1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__6256__S (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA__6257__A (.DIODE(net1577));
 sky130_fd_sc_hd__diode_2 ANTENNA__6257__B (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6258__A2 (.DIODE(net1546));
 sky130_fd_sc_hd__diode_2 ANTENNA__6258__B1 (.DIODE(net1235));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__A1 (.DIODE(net1230));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__A2 (.DIODE(net1523));
 sky130_fd_sc_hd__diode_2 ANTENNA__6260__A1 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__6260__S (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA__6261__A (.DIODE(net1576));
 sky130_fd_sc_hd__diode_2 ANTENNA__6261__B (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__A2 (.DIODE(net1522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__A2 (.DIODE(net1545));
 sky130_fd_sc_hd__diode_2 ANTENNA__6264__A1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__6264__S (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__A1 (.DIODE(net1224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__A2 (.DIODE(m1_wbd_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__B1 (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6266__A1 (.DIODE(net1224));
 sky130_fd_sc_hd__diode_2 ANTENNA__6266__B1 (.DIODE(m0_wbd_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6266__B2 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6267__A1 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA__6267__S (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA__6268__A2 (.DIODE(net1544));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__A2 (.DIODE(net1521));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__B1 (.DIODE(net1575));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__B2 (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__A1 (.DIODE(net2029));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__S (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__A (.DIODE(net1573));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__B (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6272__A2 (.DIODE(net1542));
 sky130_fd_sc_hd__diode_2 ANTENNA__6272__B1 (.DIODE(net1237));
 sky130_fd_sc_hd__diode_2 ANTENNA__6273__A2 (.DIODE(net1520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6274__A1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__6274__S (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__A2 (.DIODE(net1541));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__A1 (.DIODE(net1231));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__A2 (.DIODE(net1519));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__B1 (.DIODE(net1572));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__B2 (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__A1 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__S (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA__6278__A0 (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.mem[3][50] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6278__A1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__6278__S (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA__6279__A1 (.DIODE(net1238));
 sky130_fd_sc_hd__diode_2 ANTENNA__6279__A2 (.DIODE(m2_wbd_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6279__B1 (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6279__B2 (.DIODE(m3_wbd_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6279__C1 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6280__A1 (.DIODE(net1883));
 sky130_fd_sc_hd__diode_2 ANTENNA__6281__A1 (.DIODE(net1598));
 sky130_fd_sc_hd__diode_2 ANTENNA__6281__A2 (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6282__A1 (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__6282__S (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA__6283__A (.DIODE(net1410));
 sky130_fd_sc_hd__diode_2 ANTENNA__6283__B (.DIODE(net1408));
 sky130_fd_sc_hd__diode_2 ANTENNA__6283__C (.DIODE(m3_wbd_adr_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__A1 (.DIODE(net1233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__A2 (.DIODE(net1931));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__B1 (.DIODE(m1_wbd_adr_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__B2 (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__C1 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6285__A1 (.DIODE(net1597));
 sky130_fd_sc_hd__diode_2 ANTENNA__6285__A2 (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__A1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__S (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__A (.DIODE(\u_s2.gnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__B (.DIODE(net1408));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__C (.DIODE(m3_wbd_adr_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__A1 (.DIODE(net1238));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__A2 (.DIODE(net1917));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__B1 (.DIODE(m1_wbd_adr_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__C1 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6289__A1 (.DIODE(net1596));
 sky130_fd_sc_hd__diode_2 ANTENNA__6289__A2 (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__A1 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__S (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA__6291__A (.DIODE(m1_wbd_adr_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__A1 (.DIODE(net1233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__A2 (.DIODE(net1887));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__B1 (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__B2 (.DIODE(m3_wbd_adr_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__C1 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6293__A1 (.DIODE(net1595));
 sky130_fd_sc_hd__diode_2 ANTENNA__6293__A2 (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6294__A1 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__6294__S (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__A (.DIODE(net1409));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__B (.DIODE(\u_s2.gnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__C (.DIODE(m3_wbd_adr_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6296__A1 (.DIODE(net1233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6296__A2 (.DIODE(m2_wbd_adr_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6296__B1 (.DIODE(m1_wbd_adr_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6296__B2 (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6296__C1 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__A1 (.DIODE(net1832));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__A2 (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__A1 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__S (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__A (.DIODE(m1_wbd_adr_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6300__A1 (.DIODE(net1238));
 sky130_fd_sc_hd__diode_2 ANTENNA__6300__A2 (.DIODE(m2_wbd_adr_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6300__B1 (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6300__B2 (.DIODE(m3_wbd_adr_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6300__C1 (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__A1 (.DIODE(net1594));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__A2 (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6302__A1 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__6302__S (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__A (.DIODE(m1_wbd_adr_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__B (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6304__A1 (.DIODE(net1233));
 sky130_fd_sc_hd__diode_2 ANTENNA__6304__B1 (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6304__B2 (.DIODE(m3_wbd_adr_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6304__C1 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6305__A1 (.DIODE(net1946));
 sky130_fd_sc_hd__diode_2 ANTENNA__6305__A2 (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6306__A1 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA__6306__S (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA__6307__A (.DIODE(net1409));
 sky130_fd_sc_hd__diode_2 ANTENNA__6307__B (.DIODE(net1407));
 sky130_fd_sc_hd__diode_2 ANTENNA__6307__C (.DIODE(m3_wbd_adr_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6308__A1 (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6308__B1 (.DIODE(net2032));
 sky130_fd_sc_hd__diode_2 ANTENNA__6308__B2 (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6308__C1 (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__A1 (.DIODE(net1954));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__A2 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__A1 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__S (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__A (.DIODE(net1409));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__B (.DIODE(net1407));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__C (.DIODE(m3_wbd_adr_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__A1 (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__A2 (.DIODE(m2_wbd_adr_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__B1 (.DIODE(m1_wbd_adr_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__B2 (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__C1 (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6313__A1 (.DIODE(m0_wbd_adr_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6313__A2 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6314__A1 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__6314__S (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA__6315__A1 (.DIODE(_2426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6315__S (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__6316__A1 (.DIODE(_1912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6316__S (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__6317__A1 (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6317__S (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__6318__A1 (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6318__S (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__6319__A1 (.DIODE(_1909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6319__S (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__6320__A1 (.DIODE(_1908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6320__S (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__A1 (.DIODE(_1907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__S (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__A1 (.DIODE(_1906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__S (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__A1 (.DIODE(_1905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__S (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__6324__A1 (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6324__S (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__6325__A1 (.DIODE(_2427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6325__S (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__A1 (.DIODE(_2428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__S (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__6327__A1 (.DIODE(_2429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6327__S (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__S (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__6330__S (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__S (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__6332__S (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__6333__S (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__6334__A1 (.DIODE(_2436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6334__S (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__S (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__A1 (.DIODE(_2438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__S (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__6337__A1 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6337__S (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__S (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__6339__A1 (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6339__S (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__S (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__6341__S (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__6342__S (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__S (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__A1 (.DIODE(_2446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__S (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__6345__A1 (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6345__S (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__A1 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__S (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__S (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__S (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__6349__S (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__S (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__6351__S (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__A1 (.DIODE(_2454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__S (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__6353__A1 (.DIODE(_2455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6353__S (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__A1 (.DIODE(_2456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__S (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__6355__S (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__6356__A1 (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6356__S (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__S (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__A1 (.DIODE(_2460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__S (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__A1 (.DIODE(_2461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__S (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__A1 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__S (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__A1 (.DIODE(_2007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__S (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__A1 (.DIODE(_2463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__S (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__A1 (.DIODE(_2464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__S (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__A1 (.DIODE(_2465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__S (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__A1 (.DIODE(_2466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__S (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__S (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__A1 (.DIODE(_2469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__S (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__A1 (.DIODE(_2470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__S (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__A1 (.DIODE(_2471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__S (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__A1 (.DIODE(_2472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__S (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__A1 (.DIODE(_2473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__S (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__A1 (.DIODE(_2474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__S (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__A1 (.DIODE(_2475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__S (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__6375__A1 (.DIODE(_2476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__A1 (.DIODE(_2477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__S (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__6377__A1 (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6377__S (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__6378__S (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__A1 (.DIODE(_2481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__S (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__A1 (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__S (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__A1 (.DIODE(_2483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__S (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__6383__A1 (.DIODE(_2484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__A1 (.DIODE(_2485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__S (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__6385__A1 (.DIODE(_2486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6386__A1 (.DIODE(_2487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__A1 (.DIODE(_2488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__S (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__6388__A1 (.DIODE(_2489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6388__S (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__6389__A1 (.DIODE(_2490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6390__A1 (.DIODE(_2491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6391__A1 (.DIODE(_2492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A (.DIODE(_1704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__B (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__C_N (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__6395__S (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__A1 (.DIODE(net1924));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__S (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__A1 (.DIODE(net1929));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__S (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__6398__S (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__6399__A1 (.DIODE(net1911));
 sky130_fd_sc_hd__diode_2 ANTENNA__6399__S (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__A1 (.DIODE(net1936));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__S (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__A1 (.DIODE(net1942));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__S (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__6402__S (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__A1 (.DIODE(net1938));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__S (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__6404__S (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__A1 (.DIODE(net2044));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__S (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__6406__S (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__6407__S (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__6408__S (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__S (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__6410__A1 (.DIODE(net1920));
 sky130_fd_sc_hd__diode_2 ANTENNA__6410__S (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__A1 (.DIODE(net1921));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__S (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__S (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__A1 (.DIODE(net1923));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__S (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__6414__A1 (.DIODE(net1877));
 sky130_fd_sc_hd__diode_2 ANTENNA__6414__S (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__6415__S (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__A1 (.DIODE(net1862));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__S (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__6417__A1 (.DIODE(net1871));
 sky130_fd_sc_hd__diode_2 ANTENNA__6417__S (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__S (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__A1 (.DIODE(net1875));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__S (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__S (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__A1 (.DIODE(net2048));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__S (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__6422__A1 (.DIODE(net1873));
 sky130_fd_sc_hd__diode_2 ANTENNA__6422__S (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__6423__S (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__6424__S (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__A1 (.DIODE(net1872));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__S (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__S (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__S (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__6429__A0 (.DIODE(net1924));
 sky130_fd_sc_hd__diode_2 ANTENNA__6429__S (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__6430__A0 (.DIODE(net1929));
 sky130_fd_sc_hd__diode_2 ANTENNA__6430__S (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__S (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__A0 (.DIODE(net1911));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__S (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__A0 (.DIODE(net1936));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__S (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__A0 (.DIODE(net1942));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__S (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__S (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__A0 (.DIODE(net1938));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__S (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__S (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__6438__S (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__S (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__6440__S (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__6441__S (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__S (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__A0 (.DIODE(net1920));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__S (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__A0 (.DIODE(net1921));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__S (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__6445__S (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__6446__A0 (.DIODE(net1923));
 sky130_fd_sc_hd__diode_2 ANTENNA__6446__S (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__A0 (.DIODE(net1877));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__S (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__S (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__6449__A0 (.DIODE(net1862));
 sky130_fd_sc_hd__diode_2 ANTENNA__6449__S (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__S (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__S (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__6452__A0 (.DIODE(net2045));
 sky130_fd_sc_hd__diode_2 ANTENNA__6452__S (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__6453__S (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__A0 (.DIODE(net2048));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__S (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__6455__A0 (.DIODE(net1873));
 sky130_fd_sc_hd__diode_2 ANTENNA__6455__S (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__6456__S (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__6457__S (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__A0 (.DIODE(net1872));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__S (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__6459__S (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__6461__S (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6462__A0 (.DIODE(net1924));
 sky130_fd_sc_hd__diode_2 ANTENNA__6462__S (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__A0 (.DIODE(net1929));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__S (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6464__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__A0 (.DIODE(net1911));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__S (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6466__A0 (.DIODE(net1936));
 sky130_fd_sc_hd__diode_2 ANTENNA__6466__S (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__6467__A0 (.DIODE(net1942));
 sky130_fd_sc_hd__diode_2 ANTENNA__6467__S (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6468__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__A0 (.DIODE(net1938));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__S (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__6471__A0 (.DIODE(net2044));
 sky130_fd_sc_hd__diode_2 ANTENNA__6471__S (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__6472__S (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__6473__S (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__6474__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__S (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__A0 (.DIODE(net1920));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__S (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6477__A0 (.DIODE(net1921));
 sky130_fd_sc_hd__diode_2 ANTENNA__6477__S (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6478__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__A0 (.DIODE(net1923));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__S (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__A0 (.DIODE(net2042));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__S (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__6482__A0 (.DIODE(net1862));
 sky130_fd_sc_hd__diode_2 ANTENNA__6482__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__A0 (.DIODE(net1871));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__S (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__S (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__6485__A0 (.DIODE(net1875));
 sky130_fd_sc_hd__diode_2 ANTENNA__6485__S (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__6486__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__A0 (.DIODE(net2048));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__S (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__A0 (.DIODE(net1873));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__S (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__6489__S (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__6490__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__6491__A0 (.DIODE(net1872));
 sky130_fd_sc_hd__diode_2 ANTENNA__6491__S (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__6494__S (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__A0 (.DIODE(net1924));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__S (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__6496__A0 (.DIODE(net1929));
 sky130_fd_sc_hd__diode_2 ANTENNA__6496__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__6497__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6498__A0 (.DIODE(net1911));
 sky130_fd_sc_hd__diode_2 ANTENNA__6498__S (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__6499__A0 (.DIODE(net1936));
 sky130_fd_sc_hd__diode_2 ANTENNA__6499__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__6500__A0 (.DIODE(net1942));
 sky130_fd_sc_hd__diode_2 ANTENNA__6500__S (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__S (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__6502__A0 (.DIODE(net1938));
 sky130_fd_sc_hd__diode_2 ANTENNA__6502__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__S (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__6504__A0 (.DIODE(net2044));
 sky130_fd_sc_hd__diode_2 ANTENNA__6504__S (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__6505__S (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__6506__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6507__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__S (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__6509__A0 (.DIODE(net1920));
 sky130_fd_sc_hd__diode_2 ANTENNA__6509__S (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__6510__A0 (.DIODE(net1921));
 sky130_fd_sc_hd__diode_2 ANTENNA__6510__S (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__6511__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__A0 (.DIODE(net1923));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__S (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__A0 (.DIODE(net1877));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__S (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__6514__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__A0 (.DIODE(net1862));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6516__A0 (.DIODE(net1871));
 sky130_fd_sc_hd__diode_2 ANTENNA__6516__S (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__6517__S (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__6518__A0 (.DIODE(net2045));
 sky130_fd_sc_hd__diode_2 ANTENNA__6518__S (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__6519__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__A0 (.DIODE(net2048));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__S (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__6521__A0 (.DIODE(net1873));
 sky130_fd_sc_hd__diode_2 ANTENNA__6521__S (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__6522__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6523__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6524__A0 (.DIODE(net1872));
 sky130_fd_sc_hd__diode_2 ANTENNA__6524__S (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__6525__S (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__6526__A2 (.DIODE(_1781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__A (.DIODE(m1_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__6529__A (.DIODE(m3_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__6530__B1 (.DIODE(_1781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6531__A (.DIODE(_3258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__A2 (.DIODE(_3256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6534__A2_N (.DIODE(_1781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6535__B1 (.DIODE(_3258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6536__A2 (.DIODE(_3256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6538__A (.DIODE(\u_s1.u_sync_wbb.m_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6539__A (.DIODE(\u_s1.u_sync_wbb.m_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6540__A (.DIODE(\u_s1.u_sync_wbb.m_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6540__B (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA__6541__A0 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA__6541__S (.DIODE(\u_s1.u_sync_wbb.m_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6542__A1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__6542__A3 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA__6542__B1 (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6543__A0 (.DIODE(\u_s1.u_sync_wbb.wbm_ack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6545__A (.DIODE(\u_s1.u_sync_wbb.m_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6545__B (.DIODE(_1892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__A1 (.DIODE(\u_s1.u_sync_wbb.m_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__B1 (.DIODE(_1902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__B2 (.DIODE(\u_s1.u_sync_wbb.wbm_lack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6547__A1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__6547__A3 (.DIODE(_3265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6548__A0 (.DIODE(\u_s1.u_sync_wbb.wbm_lack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6549__A (.DIODE(_1903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6549__B (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA__6551__A1 (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6552__A2 (.DIODE(\u_s1.u_sync_wbb.m_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6552__B1_N (.DIODE(_1903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6553__A1 (.DIODE(\u_s1.u_sync_wbb.m_resp_rd_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__A2 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__B1 (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6555__A1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA__6556__A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__6557__A1 (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6557__S (.DIODE(net1799));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__A1 (.DIODE(\u_s2.u_sync_wbb.m_bl_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__S (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__A1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__B1_N (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA__6560__A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA__6560__B (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__6561__C (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA__6562__A (.DIODE(\u_s2.u_sync_wbb.m_bl_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6563__A (.DIODE(\u_s2.u_sync_wbb.m_bl_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__A1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__B1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__6565__A1_N (.DIODE(_3283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6565__B2 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__6566__A (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__6566__B (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA__6566__C (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__6567__B1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__A1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__A1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__B1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__B2 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__6573__B1_N (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__6574__A_N (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__6576__A (.DIODE(\u_s2.u_sync_wbb.m_bl_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__A (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA__6578__A1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA__6578__C1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__A2 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__B (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__A1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__B1 (.DIODE(_3299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__C1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA__6582__B1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA__6584__A (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__A2 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__A1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__A2 (.DIODE(_3299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__B1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__A1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__A2 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__A3 (.DIODE(_3299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__B1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__A (.DIODE(\u_s2.u_sync_wbb.m_bl_cnt[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__B1 (.DIODE(\u_s2.u_sync_wbb.m_bl_cnt[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__A1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__B1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__A1_N (.DIODE(_3306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__B1 (.DIODE(\u_s2.u_sync_wbb.m_bl_cnt[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__B2 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__A1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__A3 (.DIODE(_3299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6594__B (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__6594__D (.DIODE(_3299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6595__A (.DIODE(\u_s2.u_sync_wbb.m_bl_cnt[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6596__A (.DIODE(\u_s2.u_sync_wbb.m_bl_cnt[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6597__A (.DIODE(_2921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6598__A1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA__6598__C1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__6599__A1 (.DIODE(\u_s2.u_sync_wbb.m_bl_cnt[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6599__A2 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__6599__B1_N (.DIODE(_3315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6600__A2 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__6600__A4 (.DIODE(_3299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__C (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__D_N (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__A (.DIODE(\u_s2.u_sync_wbb.m_bl_cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__A (.DIODE(\u_s2.u_sync_wbb.m_bl_cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__A (.DIODE(_2921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__C (.DIODE(_3319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__A1 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__A3 (.DIODE(_3317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__C1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__A1 (.DIODE(\u_s2.u_sync_wbb.m_bl_cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__A2 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__A (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__A1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__A2 (.DIODE(_3322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__B1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__A1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__A2 (.DIODE(_3317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6610__B (.DIODE(_3319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__B (.DIODE(_3319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__A1 (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__B1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__A2 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__B1 (.DIODE(_3324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__A1 (.DIODE(_2921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__B1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__A2 (.DIODE(_3322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__B1_N (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__A_N (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__C (.DIODE(_3322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__A (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__C_N (.DIODE(\u_s2.u_sync_wbb.m_bl_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__A1 (.DIODE(_2921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__A2 (.DIODE(_3329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__A3 (.DIODE(_3330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__A1 (.DIODE(\u_s2.u_sync_wbb.m_bl_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__B2 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__6622__A (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__B (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__A (.DIODE(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__A_N (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__A (.DIODE(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__B (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__A (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__C_N (.DIODE(\u_s2.u_sync_wbb.m_cmd_wr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__A0 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__S (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__A0 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__S (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA__6632__A0 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__6632__S (.DIODE(_3336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__A0 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__S (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__A0 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__S (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__A0 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__S (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__A0 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__S (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__A0 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__S (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__A0 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__S (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__A0 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__S (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__A0 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__S (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__A0 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__S (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__A0 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__S (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__A0 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__S (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA__6644__A0 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__6644__S (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__6645__A0 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA__6645__S (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA__6646__A0 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__6646__S (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA__6647__A0 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA__6647__S (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA__6648__A0 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA__6648__S (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__6649__A0 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__6649__A1 (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.mem[0][24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6649__S (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__6650__A0 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__6650__S (.DIODE(_3336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__A0 (.DIODE(_3164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__S (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__A0 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__S (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA__6653__A0 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__6653__S (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA__6654__A0 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__6654__S (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__A0 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__S (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA__6656__A0 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__6656__S (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__A0 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__S (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__A0 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__S (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__A0 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__S (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA__6660__A0 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA__6660__S (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA__6661__A0 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__6661__S (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__A0 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__S (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__A0 (.DIODE(_3195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__S (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA__6664__A0 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__6664__S (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__A0 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__S (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA__6666__A0 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__6666__S (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA__6667__A0 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__6667__S (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__A0 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__S (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__A0 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__S (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__A0 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__S (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__A0 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__S (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__A0 (.DIODE(_3216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__S (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__A0 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__S (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__A0 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__S (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__A0 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__S (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__A0 (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__A1 (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.mem[0][53] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__S (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__A0 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__S (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__A0 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__S (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__A0 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__S (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__A0 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__S (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__A0 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__S (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__A0 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__S (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__A0 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__S (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__A0 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__S (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__C (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__6688__B (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__A (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__C (.DIODE(_2791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__D_N (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__A (.DIODE(_2796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__C (.DIODE(_2798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__A1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__B1 (.DIODE(_1704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__A (.DIODE(net1361));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__B (.DIODE(net1506));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__A1 (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__A2 (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__B1 (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__A (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__B (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__C (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__B (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__B (.DIODE(_3344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__A (.DIODE(net1350));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__B (.DIODE(\u_s1.u_sync_wbb.m_resp_rd_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__A1 (.DIODE(net1349));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__A2 (.DIODE(\u_s1.u_sync_wbb.m_resp_rd_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__B1 (.DIODE(net1345));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__A (.DIODE(net1346));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__B (.DIODE(net1350));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__C (.DIODE(\u_s1.u_sync_wbb.m_resp_rd_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__A (.DIODE(\u_s1.u_sync_wbb.u_resp_if.rd_ptr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__A (.DIODE(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__B (.DIODE(\u_s0.u_sync_wbb.m_cmd_wr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6703__A (.DIODE(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6703__B (.DIODE(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6703__C (.DIODE(\u_s0.u_sync_wbb.m_cmd_wr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__A1 (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__S (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__A1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__S (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA__6706__A1 (.DIODE(_1792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6706__S (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__A1 (.DIODE(_1794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__S (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA__6708__A1 (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6708__S (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__A1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__S (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__A1 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__S (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__A1 (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__S (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__A1 (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__S (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__A1 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__S (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA__6714__A1 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6714__S (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__S (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__A1 (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__S (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__A1 (.DIODE(_2957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__S (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__S (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__A1 (.DIODE(_2962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__S (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA__6720__A1 (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6720__S (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__A1 (.DIODE(_2966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__S (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__S (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__S (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA__6724__S (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA__6725__A1 (.DIODE(_2976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6725__S (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__6726__S (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__S (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__S (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__S (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__A1 (.DIODE(_2988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__S (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA__6731__A1 (.DIODE(_2991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6731__S (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA__6732__S (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__S (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__A1 (.DIODE(_2998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__S (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__A1 (.DIODE(_3001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__S (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__A1 (.DIODE(_3004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__S (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__S (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__A1 (.DIODE(_3010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__S (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA__6739__A1 (.DIODE(_3012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6739__S (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA__6740__A1 (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6740__S (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__A1 (.DIODE(_3016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__S (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA__6742__S (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA__6743__S (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA__6744__A1 (.DIODE(_3024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6744__S (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__S (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__A1 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__S (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__A1 (.DIODE(_3031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__S (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__6748__S (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA__6749__S (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA__6750__A1 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6750__S (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA__6751__S (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__A1 (.DIODE(_3041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__S (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__A1 (.DIODE(_3044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__S (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__A1 (.DIODE(_3047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__S (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__6755__A1 (.DIODE(_3050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6755__S (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA__6756__A1 (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6756__S (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__S (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__6758__S (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA__6759__S (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__S (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__A1 (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__S (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__S (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__S (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__S (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__A1 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__S (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__A1 (.DIODE(_3083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__S (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA__6767__S (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__S (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__A1 (.DIODE(_3092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__S (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__A1 (.DIODE(_3095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__S (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__A1 (.DIODE(_3098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__S (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__S (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__S (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__S (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__S (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA__6776__S (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA__6777__S (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA__6778__S (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA__6779__S (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__S (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__A_N (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__C (.DIODE(\u_s2.u_sync_wbb.m_cmd_wr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__A0 (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.mem[2][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__S (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__A1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__S (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__S (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__A1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__S (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__A1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__S (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__A1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__S (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__S (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA__6789__A1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__6789__S (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA__6790__A1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__6790__S (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__A1 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__S (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__A1 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__S (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA__6793__A1 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA__6793__S (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__A1 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__S (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA__6795__A1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__6795__S (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__A1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__S (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA__6797__A1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA__6797__S (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA__6798__A1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__6798__S (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__6799__A1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA__6799__S (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA__6800__A1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA__6800__S (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__A1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__S (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__A1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__S (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA__6803__A1 (.DIODE(_3164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6803__S (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA__6804__A1 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA__6804__S (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__A1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__S (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA__6806__A1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__6806__S (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA__6807__A1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__6807__S (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__6808__A1 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__6808__S (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA__6809__A1 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA__6809__S (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA__6810__A1 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA__6810__S (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__A1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__S (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__A1 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__S (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA__6813__A1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__6813__S (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__A1 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__S (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA__6815__A1 (.DIODE(_3195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6815__S (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__A1 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__S (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__A1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__S (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__6818__A1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__6818__S (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA__6819__A1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__6819__S (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__A1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__S (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__6821__A1 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__6821__S (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA__6822__A1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__6822__S (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA__6823__A1 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA__6823__S (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__A1 (.DIODE(net2029));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__S (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA__6825__A1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__6825__S (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA__6826__A1 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__6826__S (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA__6827__A0 (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.mem[2][50] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6827__A1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__6827__S (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA__6828__A1 (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__6828__S (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA__6829__A1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__6829__S (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__6830__A0 (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.mem[2][55] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6830__A1 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__6830__S (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__6831__A1 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__6831__S (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA__6832__A1 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__6832__S (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__6833__A1 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__6833__S (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__A1 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__S (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__A1 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__S (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA__6836__A1 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__6836__S (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA__6837__C (.DIODE(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6838__A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__6838__S (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA__6839__A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__6839__S (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA__6840__A1 (.DIODE(_1860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6840__S (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA__6841__A1 (.DIODE(_1856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6841__S (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA__6842__A1 (.DIODE(_1869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6842__S (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA__6843__A1 (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6843__S (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__6844__A1 (.DIODE(_1867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6844__S (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA__6845__A1 (.DIODE(_1866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6845__S (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__6846__A1 (.DIODE(_1873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6846__S (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA__6847__A1 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA__6847__S (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA__6848__A1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__6848__S (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA__6849__A1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__6849__S (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA__6850__A1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__6850__S (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__6851__A1 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA__6851__S (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__A1 (.DIODE(_2816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__S (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__6853__A1 (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6853__S (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA__6854__A1 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA__6854__S (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__A1 (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__S (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA__6856__A1 (.DIODE(_2825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6856__S (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__S (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__A1 (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__S (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA__6859__A1 (.DIODE(_2832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6859__S (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA__6860__A1 (.DIODE(_2835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6860__S (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__A1 (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__S (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA__6862__A1 (.DIODE(_2841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6862__S (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA__6863__A1 (.DIODE(_2844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6863__S (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__A1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__S (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA__6865__A1 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6865__S (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__6866__A1 (.DIODE(_2851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6866__S (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA__6867__A1 (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6867__S (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__6868__A1 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6868__S (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA__6869__A1 (.DIODE(_2858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6869__S (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA__6870__A1 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6870__S (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__6871__A1 (.DIODE(_2863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6871__S (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__S (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__A1 (.DIODE(_2867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__S (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__A1 (.DIODE(_2869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__S (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__6875__A1 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA__6875__S (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA__6876__A1 (.DIODE(net2080));
 sky130_fd_sc_hd__diode_2 ANTENNA__6876__S (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA__6877__A1 (.DIODE(_2875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6877__S (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__A1 (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__S (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA__6879__A1 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA__6879__S (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__A1 (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__S (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA__6881__S (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA__6882__A1 (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6882__S (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA__6883__A1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__6883__S (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA__6884__A1 (.DIODE(_2888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6884__S (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA__6885__A1 (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6885__S (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA__6886__A1 (.DIODE(_2894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6886__S (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA__6887__A1 (.DIODE(_2897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6887__S (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA__6888__A1 (.DIODE(_2900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6888__S (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA__6889__A1 (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6889__S (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA__6890__A1 (.DIODE(_2906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6890__S (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA__6891__A_N (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__6891__B (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__6891__C (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__6892__A0 (.DIODE(\u_reg.reg_7[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6892__A1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA__6892__S (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6893__A1 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA__6893__S (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6894__A1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA__6894__S (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6895__A1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA__6895__S (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6896__A1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA__6896__S (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6897__A1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__6897__S (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6898__A1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA__6898__S (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6899__A1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA__6901__A (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6901__B (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__A_N (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__B (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__C (.DIODE(_2589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6903__A (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6905__A0 (.DIODE(\u_s0.u_sync_wbb.wbm_ack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6905__S (.DIODE(_3352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6906__B1 (.DIODE(_3352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6907__A1 (.DIODE(\u_s0.u_sync_wbb.m_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6907__B2 (.DIODE(\u_s0.u_sync_wbb.wbm_lack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6909__A0 (.DIODE(\u_s0.u_sync_wbb.wbm_lack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6909__S (.DIODE(_3357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6910__A1 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6910__B2 (.DIODE(\u_s0.u_sync_wbb.m_cmd_wr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6911__A1 (.DIODE(\u_s0.u_sync_wbb.m_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6912__B2 (.DIODE(\u_s0.u_sync_wbb.m_resp_rd_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6913__B1 (.DIODE(_1892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6913__B2 (.DIODE(\u_s1.u_sync_wbb.m_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__A1 (.DIODE(_1902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__A2 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__C1 (.DIODE(_1903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6915__A1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__6915__B1 (.DIODE(_1875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6916__A (.DIODE(_1875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6916__B (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__6917__A (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6917__B (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__A1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__A2 (.DIODE(_3363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6919__A1 (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6919__S (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__6920__B (.DIODE(_3363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6921__A2 (.DIODE(_3363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6921__B1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA__6922__A1 (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6922__B1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA__6923__A1 (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6925__S (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__6926__A2 (.DIODE(_3363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6927__A3 (.DIODE(_3363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6927__B1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA__6928__A1 (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6928__B1 (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__A (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__C (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6931__B2 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA__6932__A1 (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6932__S (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__6933__A3 (.DIODE(_3363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__B (.DIODE(_1860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__C (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__D_N (.DIODE(_3363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6936__A (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6936__D (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6937__A (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA__6938__A1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA__6939__A0 (.DIODE(_3383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6939__S (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__6940__B (.DIODE(_1875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6941__A1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__6942__A1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__6943__A1 (.DIODE(_1856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6943__B1 (.DIODE(_3385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6943__C1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA__6944__B1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA__6946__A (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__6947__A2 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__6947__B1 (.DIODE(_3387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6948__A (.DIODE(_1869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6948__B (.DIODE(_3386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6949__A (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA__6952__A1 (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA__6952__A2 (.DIODE(_3393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6952__B1 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__6953__A1_N (.DIODE(_3392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6953__B2 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__6954__A1 (.DIODE(_1869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6954__A2 (.DIODE(_3386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6954__B1 (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__A1 (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__A2 (.DIODE(_1869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__A3 (.DIODE(_3386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__B1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA__6956__B (.DIODE(_3393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6957__A2 (.DIODE(_3393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6957__B1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA__6959__S (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__6960__A1 (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6960__A2 (.DIODE(_1869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6960__A3 (.DIODE(_3386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6960__B1 (.DIODE(_1867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6961__B (.DIODE(_3386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6962__A (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6963__A (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6963__C (.DIODE(_3393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6964__A (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA__6965__A1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA__6965__C1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__6966__A1 (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6966__A2 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__6967__A2 (.DIODE(_3385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6967__B2 (.DIODE(_1866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6967__C1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA__6968__A (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6969__A (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA__6970__A1 (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6971__A (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__6972__A1 (.DIODE(\u_s1.u_sync_wbb.m_bl_cnt[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6972__A2 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__6973__A_N (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__6974__A (.DIODE(_1872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6974__B (.DIODE(_3386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6974__C_N (.DIODE(_1873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6975__A2 (.DIODE(_3385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6975__B1 (.DIODE(_1873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6976__B1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA__6977__A1 (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA__6977__C1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__6979__A (.DIODE(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6979__B (.DIODE(_2423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6980__A1 (.DIODE(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6981__A (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__6982__B (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__6983__A (.DIODE(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6983__B (.DIODE(\u_s0.u_sync_wbb.m_cmd_wr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6985__A (.DIODE(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6986__A (.DIODE(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6987__B (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__6988__A (.DIODE(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6988__B (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA__6989__B (.DIODE(\u_s2.u_sync_wbb.m_cmd_wr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6989__C (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6990__A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA__6990__S (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA__6991__A1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__6991__S (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA__6992__A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__6992__S (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA__6993__A1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA__6993__S (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA__6994__A1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__6994__S (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA__6995__A1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__6995__S (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__6996__A0 (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.mem[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6996__A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__6996__S (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA__6997__A1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__6997__S (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA__6998__A1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__6998__S (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__6999__A1 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA__6999__S (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__A1 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__S (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA__7001__A1 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA__7001__S (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__7002__A1 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__7002__S (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__A1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__S (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA__7004__A1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__7004__S (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA__7005__A1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA__7005__S (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA__7006__A1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__7006__S (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__7007__A1 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA__7007__S (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA__7008__A1 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA__7008__S (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA__7009__A1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__7009__S (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA__7010__A1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__7010__S (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA__7011__A1 (.DIODE(_3164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7011__S (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__7012__A1 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA__7012__S (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__A1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__S (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__A1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__S (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__7015__A1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__7015__S (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA__7016__A1 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__7016__S (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA__7017__A1 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA__7017__S (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA__7018__A1 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA__7018__S (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__7019__A1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__7019__S (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA__7020__A1 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA__7020__S (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA__7021__A1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__7021__S (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA__7022__A1 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__7022__S (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA__7023__A1 (.DIODE(_3195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7023__S (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA__7024__A1 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__7024__S (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA__7025__A1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__7025__S (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA__7026__A1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__7026__S (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA__7027__A1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__7027__S (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__7028__A1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__7028__S (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA__7029__A1 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__7029__S (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA__7030__A1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__7030__S (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__7031__A1 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA__7031__S (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__7032__A1 (.DIODE(_3216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7032__S (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA__7033__A1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__7033__S (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__7034__A1 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__7034__S (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__7035__A1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__7035__S (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA__7036__A1 (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__7036__S (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA__7037__A1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__7037__S (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__7038__A1 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__7038__S (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA__7039__A1 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__7039__S (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA__7040__A1 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__7040__S (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA__7041__A1 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__7041__S (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA__7042__A1 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA__7042__S (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__7043__A0 (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.mem[1][60] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7043__A1 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__7043__S (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__A1 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__S (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__A (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__B (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__7046__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__7046__B (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__7046__C (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__7046__D (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__7047__A (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA__7047__B (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__7048__A2 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__7049__A (.DIODE(net1337));
 sky130_fd_sc_hd__diode_2 ANTENNA__7049__B (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__7050__A (.DIODE(net1339));
 sky130_fd_sc_hd__diode_2 ANTENNA__7050__B (.DIODE(net1329));
 sky130_fd_sc_hd__diode_2 ANTENNA__7050__C (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__7051__A1 (.DIODE(net1340));
 sky130_fd_sc_hd__diode_2 ANTENNA__7051__A2 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__7051__B1 (.DIODE(net1330));
 sky130_fd_sc_hd__diode_2 ANTENNA__7054__A (.DIODE(net1320));
 sky130_fd_sc_hd__diode_2 ANTENNA__7054__B (.DIODE(\u_s0.u_sync_wbb.m_resp_rd_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7055__A1 (.DIODE(net1320));
 sky130_fd_sc_hd__diode_2 ANTENNA__7055__A2 (.DIODE(\u_s0.u_sync_wbb.m_resp_rd_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7055__B1 (.DIODE(net1315));
 sky130_fd_sc_hd__diode_2 ANTENNA__7056__A (.DIODE(net1315));
 sky130_fd_sc_hd__diode_2 ANTENNA__7056__B (.DIODE(net1320));
 sky130_fd_sc_hd__diode_2 ANTENNA__7056__C (.DIODE(\u_s0.u_sync_wbb.m_resp_rd_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7059__A2 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__7059__B1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7060__A2 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__7060__B1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__7060__B2 (.DIODE(\u_dcg_s0.cfg_mode[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7061__A (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7061__B (.DIODE(_2779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7062__A (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7062__B (.DIODE(_2779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7063__A2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__7063__B1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__7064__A2 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__7065__B (.DIODE(_3431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7065__C (.DIODE(_3434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__A1 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__A2 (.DIODE(_3431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__B1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__7067__A2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__7067__B2 (.DIODE(_3436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7068__A2 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__7068__B1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7069__A2 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__7069__B1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__7069__B2 (.DIODE(\u_dcg_s0.cfg_mode[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7070__A2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__7070__B1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__7071__A2 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__7072__A (.DIODE(_3431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7073__A1 (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7073__A2 (.DIODE(_3431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7073__B1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__7074__A1 (.DIODE(\u_reg.reg_rdata[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7074__A2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__7075__B (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7076__A2 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__7076__B1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__7077__A2 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__7078__A2 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7078__B1 (.DIODE(_2779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7079__A2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__7079__B1 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__7080__A1 (.DIODE(m2_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__7080__A2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__7080__B2 (.DIODE(_3447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7080__C1 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__7081__A1 (.DIODE(\u_reg.reg_rdata[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7081__A2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__7082__A (.DIODE(\u_dcg_s1.cfg_mode[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7082__B (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7083__A2 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__7083__B1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__7084__A2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__7085__A2 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7085__B1 (.DIODE(_2779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7086__A1 (.DIODE(\u_reg.reg_5[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7086__A2 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__7086__B1 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__7087__A1 (.DIODE(m3_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__7087__A2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__7087__B2 (.DIODE(_3453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7087__C1 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__7088__A1 (.DIODE(\u_reg.reg_rdata[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7088__A2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__7089__A2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__7089__B1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__7089__B2 (.DIODE(\u_dcg_s2.cfg_mode[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7090__A2 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__7090__B1 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__7091__A2 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__7091__B1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7092__A2 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__7092__C1 (.DIODE(_3457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7093__A1 (.DIODE(_3458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7093__S (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__7094__A2 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__7094__B1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__7094__B2 (.DIODE(\u_dcg_s2.cfg_mode[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7095__A2 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__7095__B1 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__7096__A2 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__7096__B1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__7097__A2 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__7098__A0 (.DIODE(\u_reg.reg_rdata[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7098__S (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__7099__A2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__7099__B1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__7100__A2 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__7100__B1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7101__A2 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__7101__B1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7102__A2 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__7103__A0 (.DIODE(\u_reg.reg_rdata[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7103__A1 (.DIODE(_3466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7103__S (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__7104__A2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__7104__B1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__7104__B2 (.DIODE(\u_dcg_peri.cfg_mode[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7105__A2 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__7105__B1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7106__A2 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__7106__B1 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__7107__A2 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__7107__C1 (.DIODE(_3469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7108__S (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__7109__A2 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__7109__B1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__7110__A (.DIODE(\u_dcg_riscv.cfg_mode[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7110__B (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7111__A2 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__7112__A2 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__7112__B1 (.DIODE(_2779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7113__A1 (.DIODE(\u_reg.reg_5[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7113__A2 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__7113__B1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__7114__A1 (.DIODE(\u_dsync.out_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7114__A2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__7114__B1 (.DIODE(_3473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7114__C1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__7115__A1 (.DIODE(\u_reg.reg_rdata[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7115__A2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__7115__B1 (.DIODE(_3476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7116__A2 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7116__B1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__7117__A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__7117__B1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__7118__A2 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__7118__B1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7119__A2 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__7120__A (.DIODE(_3431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7120__B (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__7121__A2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__7121__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__7122__A2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__7122__B1 (.DIODE(_3481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7123__A2 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__7123__B1 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__7124__A2 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__7124__B1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__7125__A2 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__7125__B1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7126__A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__7126__B1 (.DIODE(_3431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7127__A1 (.DIODE(\u_dsync.out_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7127__A2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__7128__A0 (.DIODE(\u_reg.reg_rdata[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7128__A1 (.DIODE(_3487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7129__A2 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7129__B1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__7130__A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__7130__B1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__7131__A2 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__7131__B1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__7131__B2 (.DIODE(\u_reg.reg_2[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7132__A1 (.DIODE(\u_reg.reg_5[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7132__A2 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__7133__A (.DIODE(_3431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7133__B (.DIODE(_3489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7134__A1 (.DIODE(\u_dsync.out_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7134__A2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__7134__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__7135__A2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__7135__B1 (.DIODE(_3492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7136__A2 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__7136__B1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__7137__A2 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__7137__B1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__7138__A2 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__7138__B1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__7139__A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__7139__B1 (.DIODE(_3431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7140__A2 (.DIODE(_3432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7140__B1 (.DIODE(_3495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7141__A0 (.DIODE(\u_reg.reg_rdata[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7141__S (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__7142__A2 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__7142__B1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__7143__A2 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__7143__B1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__7144__A2 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__7144__B1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__7145__A2 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__7146__A (.DIODE(_3431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7147__A1 (.DIODE(\u_dsync.out_data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7147__A2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__7147__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__7148__A1 (.DIODE(\u_reg.reg_rdata[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7148__A2 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__7149__A (.DIODE(\u_dsync.out_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7149__B (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__7150__A2 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7150__B1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__7151__A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__7151__B1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__7152__A2 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__7152__B1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__7153__A2 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__7154__A1 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__7154__A2 (.DIODE(_3507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7154__B1 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__7155__B1 (.DIODE(\u_reg.reg_rdata[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7155__B2 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__7156__A2 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7156__B1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__7157__A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__7157__B1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__7157__C1 (.DIODE(_3511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7158__A2 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__7158__B1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__7159__A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__7160__A (.DIODE(_3431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7160__B (.DIODE(_3512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7161__A1 (.DIODE(\u_dsync.out_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7161__A2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__7161__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__7162__A1 (.DIODE(\u_reg.reg_rdata[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7162__A2 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__7163__A2 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__7163__B1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__7164__A1 (.DIODE(\u_reg.reg_4[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7164__A2 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__7164__B1 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__7165__A2 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7165__B1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__7166__A2 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__7167__A0 (.DIODE(\u_reg.reg_rdata[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7167__S (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__7168__A2 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__7168__B1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__7169__A1 (.DIODE(\u_reg.reg_7[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7169__A2 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7169__B1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__7170__A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__7170__B1 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__7171__A2 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__7171__C1 (.DIODE(_3523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7172__A0 (.DIODE(\u_reg.reg_rdata[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7172__S (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__7173__A2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__7173__B1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__7174__A2 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__7174__B1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7175__A2 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__7175__B1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7176__A2 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__7176__C1 (.DIODE(_3527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7177__A0 (.DIODE(\u_reg.reg_rdata[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7177__A1 (.DIODE(_3528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7177__S (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__7178__A2 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__7178__B1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__7179__A2 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__7179__B1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7180__A2 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__7180__B1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7181__A2 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__7182__A0 (.DIODE(\u_reg.reg_rdata[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7182__A1 (.DIODE(_3532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7182__S (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__7183__A2 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__7183__B1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__7184__A1 (.DIODE(\u_reg.reg_6[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7184__A2 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__7184__B1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__7185__A2 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__7185__B1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__7186__A2 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__7187__A0 (.DIODE(\u_reg.reg_rdata[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7187__S (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__7188__A2 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__7188__B1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__7189__A2 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__7189__B1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__7190__A2 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__7190__B1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__7191__A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__7192__A0 (.DIODE(\u_reg.reg_rdata[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7192__S (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__7193__A2 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__7193__B1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7194__A2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__7194__B1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__7195__A2 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__7195__B1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7196__A2 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__7196__B1 (.DIODE(_3542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7196__C1 (.DIODE(_3543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7197__A0 (.DIODE(net1290));
 sky130_fd_sc_hd__diode_2 ANTENNA__7197__A1 (.DIODE(_3544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7197__S (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__7198__B (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__7199__A2 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__7199__B1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__7200__A2 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__7200__B1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__7201__A2 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__7201__B1 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__7202__A (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__7202__C (.DIODE(_3548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7203__A1 (.DIODE(\u_reg.reg_rdata[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7203__A2 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__7203__B1 (.DIODE(_3549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7204__A2 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__7204__B1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__7205__A1 (.DIODE(\u_reg.reg_7[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7205__A2 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7205__B1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__7206__A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__7206__B1 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__7207__A2 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__7207__C1 (.DIODE(_3552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7208__A1 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__7208__S (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__7209__A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__7209__B1 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__7210__A2 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__7210__B1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__7210__B2 (.DIODE(\u_reg.cfg_dcg_ctrl[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7211__A2 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7211__B1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__7211__B2 (.DIODE(\u_reg.reg_3[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7212__A2 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__7212__C1 (.DIODE(_3556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7213__A0 (.DIODE(\u_reg.reg_rdata[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7213__A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__7213__S (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__7214__A2 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__7214__B1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__7215__A2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__7215__B1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__7216__A1 (.DIODE(\u_reg.reg_4[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7216__A2 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__7216__B1 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__7217__A2 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__7218__A0 (.DIODE(\u_reg.reg_rdata[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7218__S (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__7219__A2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__7219__B1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__7220__A2 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__7220__B1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__7221__A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__7221__B1 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__7222__A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__7222__C1 (.DIODE(_3564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7223__A0 (.DIODE(\u_reg.reg_rdata[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7223__A1 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__7223__S (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__7224__A2 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__7224__B1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__7225__A2 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__7225__B1 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__A2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__B1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__7227__A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__7227__C1 (.DIODE(_3568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7228__A0 (.DIODE(\u_reg.reg_rdata[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7228__A1 (.DIODE(_3569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7228__S (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__7229__A2 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__7229__B1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__7230__A2 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__7230__B1 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__7231__A2 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7231__B1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__7232__A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__7233__A1 (.DIODE(_3573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7233__S (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__7234__A2 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__7234__B1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__7235__A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__7235__B1 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__7236__A2 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7236__B1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__7237__A2 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__7237__C1 (.DIODE(_3576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7238__A0 (.DIODE(\u_reg.reg_rdata[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7238__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__7238__S (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__7239__A2 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__7239__B1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__7240__A2 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__7240__B1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__7241__A2 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__7241__B1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__7242__A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__7243__A0 (.DIODE(\u_reg.reg_rdata[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7243__S (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__7244__A_N (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__7244__B (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7244__C (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__7245__A0 (.DIODE(\u_dcg_s0.cfg_mode[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7245__A1 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7245__S (.DIODE(_3582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7246__A0 (.DIODE(\u_dcg_s0.cfg_mode[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7246__A1 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7246__S (.DIODE(_3582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7247__A1 (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7247__S (.DIODE(_3582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7248__A0 (.DIODE(\u_dcg_s1.cfg_mode[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7248__A1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7248__S (.DIODE(_3582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7249__A0 (.DIODE(\u_dcg_s2.cfg_mode[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7249__A1 (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7249__S (.DIODE(_3582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7250__A0 (.DIODE(\u_dcg_s2.cfg_mode[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7250__A1 (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7250__S (.DIODE(_3582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7251__A1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7251__S (.DIODE(_3582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7252__A0 (.DIODE(\u_dcg_peri.cfg_mode[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7252__A1 (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7252__S (.DIODE(_3582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7253__A_N (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__7253__B (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7253__C (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__7254__A1 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7254__S (.DIODE(_3583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7255__A1 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7255__S (.DIODE(_3583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7256__A1 (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7256__S (.DIODE(_3583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7257__A1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7257__S (.DIODE(_3583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7258__A1 (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7258__S (.DIODE(_3583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7259__A1 (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7259__S (.DIODE(_3583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7260__A1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7260__S (.DIODE(_3583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7261__A1 (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7261__S (.DIODE(_3583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7262__A_N (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__7262__B (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__7262__C (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7263__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__7263__S (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__7264__A1 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA__7264__S (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__7265__A1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7265__S (.DIODE(_3584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7266__A1 (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7266__S (.DIODE(_3584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7267__A1 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA__7267__S (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__7268__A1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__7268__S (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__7269__A1 (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7269__S (.DIODE(_3584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7270__A1 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA__7270__S (.DIODE(_3584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7271__A_N (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__7271__B (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__7271__C (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__7272__A1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA__7272__S (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__7273__A1 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA__7273__S (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__7274__A0 (.DIODE(\u_reg.reg_4[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7274__A1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA__7274__S (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__7275__A1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA__7275__S (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__7276__A1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA__7276__S (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__7277__A1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__7277__S (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__7278__A1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA__7278__S (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__7279__A1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA__7280__A_N (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA__7280__B (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__7280__C (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7280__D (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__7281__A1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA__7281__S (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__7282__A1 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA__7282__S (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__7283__A1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA__7283__S (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__7284__A1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA__7284__S (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__7285__A1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA__7285__S (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__7286__A1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__7286__S (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__7287__A1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA__7287__S (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__7288__A1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA__7288__S (.DIODE(_3586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7289__A_N (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__7289__B (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__7289__C (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__7290__A1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA__7290__S (.DIODE(_3587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7291__A1 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA__7291__S (.DIODE(_3587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7292__A1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA__7292__S (.DIODE(_3587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7293__A1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA__7293__S (.DIODE(_3587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7294__A1 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA__7294__S (.DIODE(_3587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7295__A1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__7295__S (.DIODE(_3587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7296__A1 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA__7296__S (.DIODE(_3587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7297__A1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA__7297__S (.DIODE(_3587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7298__A (.DIODE(net1511));
 sky130_fd_sc_hd__diode_2 ANTENNA__7298__B (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__7301__B1 (.DIODE(_3588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7303__B1 (.DIODE(_3588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7305__C1 (.DIODE(_3588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7306__B1 (.DIODE(_3588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7307__A (.DIODE(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7308__A0 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__7308__S (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA__7309__A0 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__7309__S (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA__7310__A0 (.DIODE(_1860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7310__S (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA__7311__A0 (.DIODE(_1856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7311__S (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA__7312__A0 (.DIODE(_1869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7312__S (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA__7313__A0 (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7313__S (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA__7314__A0 (.DIODE(_1867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7314__S (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA__7315__A0 (.DIODE(_1866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7315__S (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA__7316__A0 (.DIODE(_1873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7316__S (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA__7317__A0 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA__7317__S (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA__7318__A0 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__7318__S (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA__7319__A0 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__7319__S (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA__7320__A0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__7320__S (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA__7321__A0 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA__7321__S (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA__7322__A0 (.DIODE(_2816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7322__S (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA__7323__A0 (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7323__S (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA__7324__A0 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA__7324__S (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA__7325__A0 (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7325__S (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA__7326__A0 (.DIODE(_2825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7326__S (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA__7327__S (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA__7328__A0 (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7328__S (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA__7329__A0 (.DIODE(_2832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7329__S (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA__7330__A0 (.DIODE(_2835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7330__S (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA__7331__A0 (.DIODE(_2838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7331__S (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA__7332__A0 (.DIODE(_2841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7332__S (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA__7333__A0 (.DIODE(_2844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7333__S (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA__7334__A0 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7334__S (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA__7335__A0 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7335__S (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA__7336__A0 (.DIODE(_2851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7336__S (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA__7337__A0 (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7337__S (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA__7338__A0 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7338__S (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA__7339__A0 (.DIODE(_2858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7339__S (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA__7340__A0 (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7340__S (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA__7341__A0 (.DIODE(_2863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7341__S (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA__7342__S (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA__7343__A0 (.DIODE(_2867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7343__S (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA__7344__A0 (.DIODE(_2869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7344__S (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA__7345__A0 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA__7345__S (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA__7346__A0 (.DIODE(net2080));
 sky130_fd_sc_hd__diode_2 ANTENNA__7346__S (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA__7347__A0 (.DIODE(_2875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7347__S (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA__7348__A0 (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7348__S (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA__7349__A0 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA__7349__S (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA__7350__A0 (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7350__S (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA__7351__S (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA__7352__A0 (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7352__S (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA__7353__A0 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__7353__S (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA__7354__A0 (.DIODE(_2888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7354__S (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA__7355__A0 (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7355__S (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA__7356__A0 (.DIODE(_2894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7356__S (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA__7357__A0 (.DIODE(_2897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7357__S (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA__7358__A0 (.DIODE(_2900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7358__S (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA__7359__A0 (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7359__S (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA__7360__A0 (.DIODE(_2906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7360__S (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA__7361__A1 (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7361__S (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA__7362__A1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7362__S (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA__7363__A1 (.DIODE(_1792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7363__S (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__7364__A1 (.DIODE(_1794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7364__S (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__7365__A1 (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7365__S (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__7366__A1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA__7366__S (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__7367__A1 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7367__S (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__7368__A1 (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7368__S (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__7369__A1 (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7369__S (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__7370__A1 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7370__S (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA__7371__A1 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7371__S (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__7372__S (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA__7373__A1 (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7373__S (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA__7374__A1 (.DIODE(_2957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7374__S (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA__7375__S (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__7376__A1 (.DIODE(_2962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7376__S (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__7377__A1 (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7377__S (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__7378__A1 (.DIODE(_2966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7378__S (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__7379__S (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA__7380__S (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA__7381__S (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA__7382__A1 (.DIODE(_2976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7382__S (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__7383__S (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA__7384__S (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__7385__S (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__7386__S (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__7387__A1 (.DIODE(_2988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7387__S (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA__7388__A1 (.DIODE(_2991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7388__S (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__7389__S (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__7390__S (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA__7391__A1 (.DIODE(_2998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7391__S (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__7392__A1 (.DIODE(_3001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7392__S (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__7393__A1 (.DIODE(_3004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7393__S (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA__7394__S (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA__7395__A1 (.DIODE(_3010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7395__S (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA__7396__A1 (.DIODE(_3012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7396__S (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA__7397__A1 (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7397__S (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__7398__A1 (.DIODE(_3016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7398__S (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA__7399__S (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__7400__S (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA__7401__A1 (.DIODE(_3024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7401__S (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__7402__S (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__7403__A1 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7403__S (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA__7404__A1 (.DIODE(_3031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7404__S (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__7405__S (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA__7406__S (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA__7407__A1 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7407__S (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA__7408__S (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA__7409__A1 (.DIODE(_3041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7409__S (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__7410__A1 (.DIODE(_3044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7410__S (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA__7411__A1 (.DIODE(_3047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7411__S (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__7412__A1 (.DIODE(_3050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7412__S (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA__7413__A1 (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7413__S (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__7414__S (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__7415__S (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__7416__S (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__7417__S (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA__7418__A1 (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7418__S (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA__7419__S (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__7420__S (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__7421__S (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__7422__A1 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7422__S (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__7423__A1 (.DIODE(_3083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7423__S (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__7424__S (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__7425__S (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__7426__A1 (.DIODE(_3092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7426__S (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__7427__A1 (.DIODE(_3095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7427__S (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA__7428__A1 (.DIODE(_3098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7428__S (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__7429__S (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__7430__S (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA__7431__S (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA__7432__S (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA__7433__S (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__7434__S (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA__7435__S (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__7436__S (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__7437__S (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__7438__A_N (.DIODE(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7438__B (.DIODE(\u_s0.u_sync_wbb.m_cmd_wr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7438__C (.DIODE(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7439__A1 (.DIODE(_1786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7439__S (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA__7440__A1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7440__S (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__7441__A1 (.DIODE(_1792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7441__S (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA__7442__A1 (.DIODE(_1794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7442__S (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__7443__A1 (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7443__S (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA__7444__A1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA__7444__S (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA__7445__A1 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7445__S (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA__7446__A1 (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7446__S (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__7447__A1 (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7447__S (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__7448__A1 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7448__S (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA__7449__A1 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7449__S (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA__7450__S (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__7451__A1 (.DIODE(_2954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7451__S (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA__7452__A1 (.DIODE(_2957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7452__S (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA__7453__S (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA__7454__A1 (.DIODE(_2962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7454__S (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA__7455__A1 (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7455__S (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__7456__A1 (.DIODE(_2966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7456__S (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA__7457__S (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA__7458__S (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA__7459__S (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA__7460__A1 (.DIODE(_2976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7460__S (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA__7461__S (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA__7462__S (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA__7463__S (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA__7464__S (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__7465__A1 (.DIODE(_2988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7465__S (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__7466__A1 (.DIODE(_2991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7466__S (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA__7467__S (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__7468__S (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA__7469__S (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA__7470__A1 (.DIODE(_3001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7470__S (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA__7471__A1 (.DIODE(_3004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7471__S (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA__7472__S (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA__7473__A1 (.DIODE(_3010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7473__S (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA__7474__A1 (.DIODE(_3012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7474__S (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA__7475__A1 (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7475__S (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA__7476__A1 (.DIODE(_3016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7476__S (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA__7477__S (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA__7478__S (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA__7479__A1 (.DIODE(_3024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7479__S (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA__7480__S (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA__7481__A1 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7481__S (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA__7482__A1 (.DIODE(_3031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7482__S (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA__7483__S (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA__7484__S (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA__7485__A1 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7485__S (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA__7486__S (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA__7487__A1 (.DIODE(_3041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7487__S (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA__7488__A1 (.DIODE(_3044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7488__S (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA__7489__A1 (.DIODE(_3047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7489__S (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA__7490__A1 (.DIODE(_3050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7490__S (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA__7491__A1 (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7491__S (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA__7492__S (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA__7493__S (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA__7494__S (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA__7495__S (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__7496__A1 (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7496__S (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA__7497__S (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__7498__S (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA__7499__S (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA__7500__A1 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7500__S (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__7501__A1 (.DIODE(_3083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7501__S (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA__7502__S (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA__7503__S (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA__7504__A1 (.DIODE(_3092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7504__S (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA__7505__A1 (.DIODE(_3095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7505__S (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__7506__A1 (.DIODE(_3098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7506__S (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA__7507__S (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA__7508__S (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__7509__S (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__7510__S (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA__7511__S (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA__7512__S (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__7513__S (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA__7514__S (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA__7515__S (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA__7517__B1 (.DIODE(_3588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7519__A_N (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7519__B (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA__7519__C (.DIODE(m1_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__7520__A (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA__7522__A1 (.DIODE(m2_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__7522__A2 (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA__7522__B1 (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA__7523__A (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7524__A1 (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA__7524__A2 (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA__7525__A1 (.DIODE(m3_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__7525__A2 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA__7526__A1 (.DIODE(net1278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7527__A1 (.DIODE(m0_wbd_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__7527__A2 (.DIODE(net1278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7527__A3 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA__7529__A1 (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA__7530__CLK (.DIODE(\clknet_leaf_30_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7530__RESET_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA__7531__CLK (.DIODE(\clknet_leaf_30_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7531__RESET_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA__7532__CLK (.DIODE(\clknet_leaf_30_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7532__RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA__7533__CLK (.DIODE(\clknet_leaf_29_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7533__RESET_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA__7534__CLK (.DIODE(\clknet_leaf_29_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7534__RESET_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA__7535__CLK (.DIODE(\clknet_leaf_29_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7535__RESET_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA__7536__CLK (.DIODE(\clknet_leaf_29_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7536__RESET_B (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__7537__CLK (.DIODE(\clknet_leaf_29_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7537__RESET_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA__7538__CLK (.DIODE(\clknet_leaf_32_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7538__RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA__7539__CLK (.DIODE(\clknet_leaf_54_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7539__RESET_B (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA__7540__CLK (.DIODE(\clknet_leaf_52_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7540__RESET_B (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA__7541__CLK (.DIODE(\clknet_leaf_51_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7541__RESET_B (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA__7542__CLK (.DIODE(\clknet_leaf_53_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7542__RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__7543__CLK (.DIODE(\clknet_leaf_48_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7543__RESET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA__7544__CLK (.DIODE(\clknet_leaf_47_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7544__RESET_B (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA__7545__CLK (.DIODE(\clknet_leaf_51_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7545__RESET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA__7546__CLK (.DIODE(\clknet_leaf_42_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7546__RESET_B (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA__7547__CLK (.DIODE(\clknet_leaf_47_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7547__RESET_B (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA__7548__CLK (.DIODE(\clknet_leaf_45_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7548__RESET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA__7549__CLK (.DIODE(\clknet_leaf_49_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7549__RESET_B (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA__7550__CLK (.DIODE(\clknet_leaf_49_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7550__RESET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA__7551__CLK (.DIODE(\clknet_leaf_53_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7551__RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__7552__CLK (.DIODE(\clknet_leaf_54_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7552__RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__7553__CLK (.DIODE(\clknet_leaf_47_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7553__RESET_B (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA__7554__CLK (.DIODE(\clknet_leaf_49_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7554__RESET_B (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA__7555__CLK (.DIODE(\clknet_leaf_54_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7555__RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__7556__CLK (.DIODE(\clknet_leaf_56_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7556__RESET_B (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA__7557__CLK (.DIODE(\clknet_leaf_54_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7557__RESET_B (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA__7558__CLK (.DIODE(\clknet_leaf_53_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7558__RESET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA__7559__CLK (.DIODE(\clknet_leaf_51_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7559__RESET_B (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA__7560__CLK (.DIODE(\clknet_leaf_53_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7560__RESET_B (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA__7561__CLK (.DIODE(\clknet_leaf_51_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7561__RESET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA__7562__CLK (.DIODE(\clknet_leaf_50_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7562__RESET_B (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA__7563__CLK (.DIODE(\clknet_leaf_53_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7563__RESET_B (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA__7564__CLK (.DIODE(\clknet_leaf_56_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7565__CLK (.DIODE(\clknet_leaf_56_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7565__RESET_B (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA__7566__CLK (.DIODE(\clknet_leaf_54_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7566__RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__7567__CLK (.DIODE(\clknet_leaf_56_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7567__RESET_B (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA__7568__CLK (.DIODE(\clknet_leaf_53_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7568__RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__7569__CLK (.DIODE(\clknet_leaf_53_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7569__RESET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA__7570__CLK (.DIODE(\clknet_leaf_54_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7570__RESET_B (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA__7571__CLK (.DIODE(\clknet_leaf_57_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7571__RESET_B (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA__7572__CLK (.DIODE(\clknet_leaf_53_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7572__RESET_B (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA__7573__CLK (.DIODE(\clknet_leaf_50_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7573__RESET_B (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA__7574__CLK (.DIODE(\clknet_leaf_54_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7574__RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__7575__CLK (.DIODE(\clknet_leaf_32_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7575__RESET_B (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA__7576__CLK (.DIODE(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7576__RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA__7577__CLK (.DIODE(\clknet_leaf_54_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7577__RESET_B (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA__7578__CLK (.DIODE(\clknet_leaf_44_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7578__RESET_B (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA__7579__CLK (.DIODE(\clknet_leaf_56_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7580__CLK (.DIODE(\clknet_leaf_54_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7580__RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__7581__CLK (.DIODE(\clknet_leaf_41_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7581__RESET_B (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA__7582__CLK (.DIODE(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7582__RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA__7583__CLK (.DIODE(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7583__RESET_B (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA__7584__CLK (.DIODE(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7584__RESET_B (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA__7585__CLK (.DIODE(\clknet_leaf_107_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7585__RESET_B (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA__7586__CLK (.DIODE(\clknet_leaf_107_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7586__RESET_B (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA__7587__CLK (.DIODE(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7587__RESET_B (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__7588__CLK (.DIODE(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7588__RESET_B (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__7589__CLK (.DIODE(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7589__RESET_B (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__7590__CLK (.DIODE(\clknet_leaf_99_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7590__RESET_B (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__7591__CLK (.DIODE(\clknet_leaf_99_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7591__RESET_B (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__7592__CLK (.DIODE(\clknet_leaf_98_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7592__RESET_B (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__7593__CLK (.DIODE(\clknet_leaf_99_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7593__RESET_B (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA__7594__CLK (.DIODE(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7594__RESET_B (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__7595__CLK (.DIODE(\clknet_leaf_97_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7595__RESET_B (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA__7596__CLK (.DIODE(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7596__RESET_B (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA__7597__CLK (.DIODE(\clknet_leaf_26_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7597__RESET_B (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA__7598__CLK (.DIODE(\clknet_leaf_20_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7599__CLK (.DIODE(\clknet_leaf_2_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7600__CLK (.DIODE(\clknet_leaf_3_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7600__RESET_B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__7601__CLK (.DIODE(\clknet_leaf_18_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7601__RESET_B (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__7602__CLK (.DIODE(\clknet_leaf_18_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7602__RESET_B (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__7603__CLK (.DIODE(\clknet_leaf_2_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7603__RESET_B (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__7604__CLK (.DIODE(\clknet_leaf_2_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7604__RESET_B (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA__7605__CLK (.DIODE(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7605__RESET_B (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__7606__CLK (.DIODE(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7606__RESET_B (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__7607__CLK (.DIODE(\clknet_leaf_2_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7608__CLK (.DIODE(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7608__RESET_B (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__7609__CLK (.DIODE(\clknet_leaf_14_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7609__RESET_B (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__7610__CLK (.DIODE(\clknet_leaf_15_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7610__RESET_B (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA__7611__CLK (.DIODE(\clknet_leaf_3_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7611__RESET_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__7612__CLK (.DIODE(\clknet_leaf_4_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7612__RESET_B (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA__7613__CLK (.DIODE(\clknet_leaf_13_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7614__CLK (.DIODE(\clknet_leaf_13_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7615__CLK (.DIODE(\clknet_leaf_13_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7616__CLK (.DIODE(\clknet_leaf_20_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7616__RESET_B (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA__7617__CLK (.DIODE(\clknet_leaf_13_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7618__CLK (.DIODE(\clknet_leaf_19_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7618__RESET_B (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA__7619__CLK (.DIODE(\clknet_leaf_19_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7619__RESET_B (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA__7620__CLK (.DIODE(\clknet_leaf_19_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7621__CLK (.DIODE(\clknet_leaf_26_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7621__RESET_B (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA__7622__CLK (.DIODE(\clknet_leaf_20_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7623__CLK (.DIODE(\clknet_leaf_2_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7623__RESET_B (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA__7624__CLK (.DIODE(\clknet_leaf_3_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7624__RESET_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__7625__CLK (.DIODE(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7625__RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA__7626__CLK (.DIODE(\clknet_leaf_18_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7626__RESET_B (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA__7627__CLK (.DIODE(\clknet_leaf_2_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7627__RESET_B (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA__7628__CLK (.DIODE(\clknet_leaf_16_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7629__CLK (.DIODE(\clknet_leaf_4_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7629__RESET_B (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA__7630__CLK (.DIODE(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7630__RESET_B (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__7631__CLK (.DIODE(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7631__RESET_B (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__7632__CLK (.DIODE(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7632__RESET_B (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__7633__CLK (.DIODE(\clknet_leaf_19_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7633__RESET_B (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__7634__CLK (.DIODE(\clknet_leaf_17_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7634__RESET_B (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__7635__CLK (.DIODE(\clknet_leaf_3_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7635__RESET_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__7636__CLK (.DIODE(\clknet_leaf_15_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7636__RESET_B (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA__7637__CLK (.DIODE(\clknet_leaf_12_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7638__CLK (.DIODE(\clknet_leaf_25_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7639__CLK (.DIODE(\clknet_leaf_14_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7640__CLK (.DIODE(\clknet_leaf_26_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7640__RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA__7641__CLK (.DIODE(\clknet_leaf_20_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7641__RESET_B (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA__7642__CLK (.DIODE(\clknet_leaf_12_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7642__RESET_B (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__7643__CLK (.DIODE(\clknet_leaf_25_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7643__RESET_B (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA__7644__CLK (.DIODE(\clknet_leaf_25_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7644__RESET_B (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA__7645__CLK (.DIODE(\clknet_leaf_25_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7645__RESET_B (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA__7646__CLK (.DIODE(\clknet_leaf_20_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7646__RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA__7647__CLK (.DIODE(\clknet_leaf_16_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7647__RESET_B (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA__7648__CLK (.DIODE(\clknet_leaf_3_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7648__RESET_B (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA__7649__CLK (.DIODE(\clknet_leaf_18_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7649__RESET_B (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__7650__CLK (.DIODE(\clknet_leaf_18_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7650__RESET_B (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__7651__CLK (.DIODE(\clknet_leaf_3_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7651__RESET_B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__7652__CLK (.DIODE(\clknet_leaf_17_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7652__RESET_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA__7653__CLK (.DIODE(\clknet_leaf_4_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7653__RESET_B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__7654__CLK (.DIODE(\clknet_leaf_13_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7654__RESET_B (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__7655__CLK (.DIODE(\clknet_leaf_12_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7656__CLK (.DIODE(\clknet_leaf_26_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7657__CLK (.DIODE(\clknet_leaf_19_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7657__RESET_B (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__7658__CLK (.DIODE(\clknet_leaf_20_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7658__RESET_B (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA__7659__CLK (.DIODE(\clknet_leaf_20_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7659__RESET_B (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA__7660__CLK (.DIODE(\clknet_leaf_12_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7661__CLK (.DIODE(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7661__RESET_B (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__7662__CLK (.DIODE(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7662__RESET_B (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__7663__CLK (.DIODE(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7663__RESET_B (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__7664__CLK (.DIODE(\clknet_leaf_0_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7664__RESET_B (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__7665__CLK (.DIODE(\clknet_leaf_15_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7665__RESET_B (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA__7666__CLK (.DIODE(\clknet_leaf_15_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7666__RESET_B (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA__7667__CLK (.DIODE(\clknet_leaf_3_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7667__RESET_B (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA__7668__CLK (.DIODE(\clknet_leaf_3_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7668__RESET_B (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA__7669__CLK (.DIODE(\clknet_leaf_20_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7669__RESET_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA__7670__CLK (.DIODE(\clknet_leaf_24_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7670__RESET_B (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA__7671__CLK (.DIODE(\clknet_leaf_16_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7671__RESET_B (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA__7672__CLK (.DIODE(\clknet_leaf_3_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7672__RESET_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__7673__CLK (.DIODE(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7674__CLK (.DIODE(\clknet_leaf_18_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7674__RESET_B (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA__7675__CLK (.DIODE(\clknet_leaf_16_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7675__RESET_B (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA__7676__CLK (.DIODE(\clknet_leaf_3_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7676__RESET_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__7677__CLK (.DIODE(\clknet_leaf_14_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7677__RESET_B (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA__7678__CLK (.DIODE(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7678__RESET_B (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA__7679__CLK (.DIODE(\clknet_leaf_13_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7679__RESET_B (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA__7680__CLK (.DIODE(\clknet_leaf_26_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7681__CLK (.DIODE(\clknet_leaf_19_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7682__CLK (.DIODE(\clknet_leaf_12_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7682__RESET_B (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__7683__CLK (.DIODE(\clknet_leaf_25_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7683__RESET_B (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA__7684__CLK (.DIODE(\clknet_leaf_25_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7684__RESET_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__7685__CLK (.DIODE(\clknet_leaf_5_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7685__RESET_B (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA__7686__CLK (.DIODE(\clknet_leaf_5_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7687__CLK (.DIODE(\clknet_leaf_2_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7688__CLK (.DIODE(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7689__CLK (.DIODE(\clknet_leaf_15_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7689__RESET_B (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA__7690__CLK (.DIODE(\clknet_leaf_16_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7690__RESET_B (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA__7691__CLK (.DIODE(\clknet_leaf_15_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7691__RESET_B (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA__7692__CLK (.DIODE(\clknet_leaf_15_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7692__RESET_B (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA__7693__CLK (.DIODE(\clknet_leaf_23_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7694__CLK (.DIODE(\clknet_leaf_23_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7694__RESET_B (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__7695__CLK (.DIODE(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7696__CLK (.DIODE(\clknet_leaf_24_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7696__RESET_B (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA__7697__CLK (.DIODE(\clknet_leaf_18_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7697__RESET_B (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__7698__CLK (.DIODE(\clknet_leaf_22_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7698__RESET_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA__7699__CLK (.DIODE(\clknet_leaf_23_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7700__CLK (.DIODE(\clknet_leaf_17_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7700__RESET_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA__7701__CLK (.DIODE(\clknet_leaf_14_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7702__CLK (.DIODE(\clknet_leaf_24_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7702__RESET_B (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__7703__CLK (.DIODE(\clknet_leaf_14_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7703__RESET_B (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__7704__CLK (.DIODE(\clknet_leaf_26_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7704__RESET_B (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA__7705__CLK (.DIODE(\clknet_leaf_20_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7706__CLK (.DIODE(\clknet_leaf_19_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7707__CLK (.DIODE(\clknet_leaf_25_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7707__RESET_B (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA__7708__CLK (.DIODE(\clknet_leaf_24_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7708__RESET_B (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA__7709__CLK (.DIODE(\clknet_leaf_5_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7709__RESET_B (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA__7710__CLK (.DIODE(\clknet_leaf_2_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7710__RESET_B (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA__7711__CLK (.DIODE(\clknet_leaf_2_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7711__RESET_B (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA__7712__CLK (.DIODE(\clknet_leaf_4_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7712__RESET_B (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA__7713__CLK (.DIODE(\clknet_leaf_18_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7713__RESET_B (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__7714__CLK (.DIODE(\clknet_leaf_17_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7714__RESET_B (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__7715__CLK (.DIODE(\clknet_leaf_3_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7715__RESET_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__7716__CLK (.DIODE(\clknet_leaf_15_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7716__RESET_B (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA__7717__CLK (.DIODE(\clknet_leaf_13_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7718__CLK (.DIODE(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7719__CLK (.DIODE(\clknet_leaf_13_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7720__CLK (.DIODE(\clknet_leaf_12_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7721__CLK (.DIODE(\clknet_leaf_19_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7721__RESET_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA__7722__CLK (.DIODE(\clknet_leaf_12_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7722__RESET_B (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__7723__CLK (.DIODE(\clknet_leaf_19_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7723__RESET_B (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA__7724__CLK (.DIODE(\clknet_leaf_19_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7725__CLK (.DIODE(\clknet_leaf_24_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7725__RESET_B (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA__7726__CLK (.DIODE(\clknet_leaf_24_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7727__CLK (.DIODE(\clknet_leaf_16_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7727__RESET_B (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA__7728__CLK (.DIODE(\clknet_leaf_3_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7728__RESET_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__7729__CLK (.DIODE(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7730__CLK (.DIODE(\clknet_leaf_19_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7730__RESET_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA__7731__CLK (.DIODE(\clknet_leaf_16_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7731__RESET_B (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA__7732__CLK (.DIODE(\clknet_leaf_17_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7732__RESET_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA__7733__CLK (.DIODE(\clknet_leaf_23_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7734__CLK (.DIODE(\clknet_leaf_23_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7735__CLK (.DIODE(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7736__CLK (.DIODE(\clknet_leaf_23_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7736__RESET_B (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__7737__CLK (.DIODE(\clknet_leaf_18_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7737__RESET_B (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__7738__CLK (.DIODE(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7738__RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA__7739__CLK (.DIODE(\clknet_leaf_23_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7739__RESET_B (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__7740__CLK (.DIODE(\clknet_leaf_18_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7740__RESET_B (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__7741__CLK (.DIODE(\clknet_leaf_13_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7742__CLK (.DIODE(\clknet_leaf_25_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7742__RESET_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__7743__CLK (.DIODE(\clknet_leaf_13_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7744__CLK (.DIODE(\clknet_leaf_26_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7745__CLK (.DIODE(\clknet_leaf_19_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7745__RESET_B (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA__7746__CLK (.DIODE(\clknet_leaf_12_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7746__RESET_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA__7747__CLK (.DIODE(\clknet_leaf_25_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7747__RESET_B (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA__7748__CLK (.DIODE(\clknet_leaf_26_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7748__RESET_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA__7749__CLK (.DIODE(\clknet_leaf_20_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7750__CLK (.DIODE(\clknet_leaf_20_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7751__CLK (.DIODE(\clknet_leaf_2_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7751__RESET_B (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA__7752__CLK (.DIODE(\clknet_leaf_3_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7752__RESET_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__7753__CLK (.DIODE(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7753__RESET_B (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA__7754__CLK (.DIODE(\clknet_leaf_18_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7754__RESET_B (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA__7755__CLK (.DIODE(\clknet_leaf_3_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7755__RESET_B (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA__7756__CLK (.DIODE(\clknet_leaf_2_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7756__RESET_B (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA__7757__CLK (.DIODE(\clknet_leaf_22_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7757__RESET_B (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA__7758__CLK (.DIODE(\clknet_leaf_22_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7759__CLK (.DIODE(\clknet_leaf_18_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7759__RESET_B (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA__7760__CLK (.DIODE(\clknet_leaf_23_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7760__RESET_B (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA__7761__CLK (.DIODE(\clknet_leaf_17_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7761__RESET_B (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__7762__CLK (.DIODE(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7762__RESET_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA__7763__CLK (.DIODE(\clknet_leaf_22_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7763__RESET_B (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA__7764__CLK (.DIODE(\clknet_leaf_16_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7765__CLK (.DIODE(\clknet_leaf_42_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7766__CLK (.DIODE(\clknet_leaf_52_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7767__CLK (.DIODE(\clknet_leaf_51_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7768__CLK (.DIODE(\clknet_leaf_53_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7769__CLK (.DIODE(\clknet_leaf_48_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7770__CLK (.DIODE(\clknet_leaf_48_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7771__CLK (.DIODE(\clknet_leaf_48_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7772__CLK (.DIODE(\clknet_leaf_60_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7773__CLK (.DIODE(\clknet_leaf_49_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7774__CLK (.DIODE(\clknet_leaf_50_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7775__CLK (.DIODE(\clknet_leaf_48_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7776__CLK (.DIODE(\clknet_leaf_62_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7777__CLK (.DIODE(\clknet_leaf_51_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7778__CLK (.DIODE(\clknet_leaf_56_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7779__CLK (.DIODE(\clknet_leaf_55_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7780__CLK (.DIODE(\clknet_leaf_50_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7781__CLK (.DIODE(\clknet_leaf_55_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7782__CLK (.DIODE(\clknet_leaf_51_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7783__CLK (.DIODE(\clknet_leaf_51_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7784__CLK (.DIODE(\clknet_leaf_50_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7785__CLK (.DIODE(\clknet_leaf_50_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7786__CLK (.DIODE(\clknet_leaf_55_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7787__CLK (.DIODE(\clknet_leaf_55_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7788__CLK (.DIODE(\clknet_leaf_50_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7789__CLK (.DIODE(\clknet_leaf_62_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7790__CLK (.DIODE(\clknet_leaf_62_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7791__CLK (.DIODE(\clknet_leaf_63_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7792__CLK (.DIODE(\clknet_leaf_54_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7793__CLK (.DIODE(\clknet_leaf_63_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7794__CLK (.DIODE(\clknet_leaf_60_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7795__CLK (.DIODE(\clknet_leaf_61_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7796__CLK (.DIODE(\clknet_leaf_62_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7797__CLK (.DIODE(\clknet_leaf_42_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7798__CLK (.DIODE(\clknet_leaf_52_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7799__CLK (.DIODE(\clknet_leaf_51_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7800__CLK (.DIODE(\clknet_leaf_52_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7801__CLK (.DIODE(\clknet_leaf_48_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7802__CLK (.DIODE(\clknet_leaf_48_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7803__CLK (.DIODE(\clknet_leaf_48_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7804__CLK (.DIODE(\clknet_leaf_61_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7805__CLK (.DIODE(\clknet_leaf_50_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7806__CLK (.DIODE(\clknet_leaf_54_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7807__CLK (.DIODE(\clknet_leaf_48_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7808__CLK (.DIODE(\clknet_leaf_62_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7809__CLK (.DIODE(\clknet_leaf_49_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7810__CLK (.DIODE(\clknet_leaf_62_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7811__CLK (.DIODE(\clknet_leaf_55_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7812__CLK (.DIODE(\clknet_leaf_50_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7813__CLK (.DIODE(\clknet_leaf_54_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7814__CLK (.DIODE(\clknet_leaf_52_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7815__CLK (.DIODE(\clknet_leaf_51_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7816__CLK (.DIODE(\clknet_leaf_42_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7817__CLK (.DIODE(\clknet_leaf_49_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7818__CLK (.DIODE(\clknet_leaf_63_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7819__CLK (.DIODE(\clknet_leaf_42_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7820__CLK (.DIODE(\clknet_leaf_50_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7821__CLK (.DIODE(\clknet_leaf_63_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7822__CLK (.DIODE(\clknet_leaf_62_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7823__CLK (.DIODE(\clknet_leaf_63_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7824__CLK (.DIODE(\clknet_leaf_54_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7825__CLK (.DIODE(\clknet_leaf_63_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7826__CLK (.DIODE(\clknet_leaf_61_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7827__CLK (.DIODE(\clknet_leaf_62_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7828__CLK (.DIODE(\clknet_leaf_61_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7829__CLK (.DIODE(\clknet_leaf_42_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7830__CLK (.DIODE(\clknet_leaf_52_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7831__CLK (.DIODE(\clknet_leaf_52_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7832__CLK (.DIODE(\clknet_leaf_52_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7833__CLK (.DIODE(\clknet_leaf_47_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7834__CLK (.DIODE(\clknet_leaf_48_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7835__CLK (.DIODE(\clknet_leaf_48_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7836__CLK (.DIODE(\clknet_leaf_62_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7837__CLK (.DIODE(\clknet_leaf_50_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7838__CLK (.DIODE(\clknet_leaf_50_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7839__CLK (.DIODE(\clknet_leaf_47_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7840__CLK (.DIODE(\clknet_leaf_55_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7841__CLK (.DIODE(\clknet_leaf_48_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7842__CLK (.DIODE(\clknet_leaf_62_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7843__CLK (.DIODE(\clknet_leaf_55_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7844__CLK (.DIODE(\clknet_leaf_49_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7845__CLK (.DIODE(\clknet_leaf_50_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7846__CLK (.DIODE(\clknet_leaf_52_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7847__CLK (.DIODE(\clknet_leaf_51_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7848__CLK (.DIODE(\clknet_leaf_49_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7849__CLK (.DIODE(\clknet_leaf_49_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7850__CLK (.DIODE(\clknet_leaf_63_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7851__CLK (.DIODE(\clknet_leaf_42_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7852__CLK (.DIODE(\clknet_leaf_50_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7853__CLK (.DIODE(\clknet_leaf_63_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7854__CLK (.DIODE(\clknet_leaf_63_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7855__CLK (.DIODE(\clknet_leaf_64_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7856__CLK (.DIODE(\clknet_leaf_55_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7857__CLK (.DIODE(\clknet_leaf_41_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7858__CLK (.DIODE(\clknet_leaf_60_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7859__CLK (.DIODE(\clknet_leaf_62_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7860__CLK (.DIODE(\clknet_leaf_61_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7861__CLK (.DIODE(\clknet_leaf_42_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7862__CLK (.DIODE(\clknet_leaf_52_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7863__CLK (.DIODE(\clknet_leaf_51_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7864__CLK (.DIODE(\clknet_leaf_54_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7865__CLK (.DIODE(\clknet_leaf_48_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7866__CLK (.DIODE(\clknet_leaf_48_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7867__CLK (.DIODE(\clknet_leaf_49_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7868__CLK (.DIODE(\clknet_leaf_61_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7869__CLK (.DIODE(\clknet_leaf_49_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7870__CLK (.DIODE(\clknet_leaf_54_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7871__CLK (.DIODE(\clknet_leaf_47_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7872__CLK (.DIODE(\clknet_leaf_62_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7873__CLK (.DIODE(\clknet_leaf_48_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7874__CLK (.DIODE(\clknet_leaf_55_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7875__CLK (.DIODE(\clknet_leaf_55_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7876__CLK (.DIODE(\clknet_leaf_55_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7877__CLK (.DIODE(\clknet_leaf_55_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7878__CLK (.DIODE(\clknet_leaf_52_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7879__CLK (.DIODE(\clknet_leaf_50_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7880__CLK (.DIODE(\clknet_leaf_42_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7881__CLK (.DIODE(\clknet_leaf_49_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7882__CLK (.DIODE(\clknet_leaf_55_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7883__CLK (.DIODE(\clknet_leaf_42_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7884__CLK (.DIODE(\clknet_leaf_54_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7885__CLK (.DIODE(\clknet_leaf_63_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7886__CLK (.DIODE(\clknet_leaf_62_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7887__CLK (.DIODE(\clknet_leaf_64_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7888__CLK (.DIODE(\clknet_leaf_54_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7889__CLK (.DIODE(\clknet_leaf_41_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7890__CLK (.DIODE(\clknet_leaf_61_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7891__CLK (.DIODE(\clknet_leaf_61_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7892__CLK (.DIODE(\clknet_leaf_61_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7893__CLK (.DIODE(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7893__RESET_B (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__7894__CLK (.DIODE(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7894__RESET_B (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA__7895__CLK (.DIODE(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7895__RESET_B (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__7896__CLK (.DIODE(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7896__RESET_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__7897__CLK (.DIODE(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7897__RESET_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__7898__CLK (.DIODE(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7898__RESET_B (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA__7899__CLK (.DIODE(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7899__RESET_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__7900__CLK (.DIODE(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7900__RESET_B (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA__7901__CLK (.DIODE(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7901__RESET_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__7902__CLK (.DIODE(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7902__RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__7903__CLK (.DIODE(\clknet_leaf_96_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7903__RESET_B (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA__7904__CLK (.DIODE(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7904__RESET_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__7905__CLK (.DIODE(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7905__RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__7906__CLK (.DIODE(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7906__RESET_B (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__7907__CLK (.DIODE(\clknet_leaf_72_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7907__RESET_B (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA__7908__CLK (.DIODE(\clknet_leaf_64_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7908__RESET_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__7909__CLK (.DIODE(\clknet_leaf_64_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7909__RESET_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__7910__CLK (.DIODE(\clknet_leaf_64_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7910__RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__7911__CLK (.DIODE(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7911__RESET_B (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__7912__CLK (.DIODE(\clknet_leaf_72_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7912__RESET_B (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA__7913__CLK (.DIODE(\clknet_leaf_64_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7913__RESET_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__7914__CLK (.DIODE(\clknet_leaf_64_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7914__RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__7915__CLK (.DIODE(\clknet_leaf_64_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7915__RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__7916__CLK (.DIODE(\clknet_leaf_64_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7916__RESET_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__7917__CLK (.DIODE(\clknet_leaf_61_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7917__RESET_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__7918__CLK (.DIODE(\clknet_leaf_63_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7918__RESET_B (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA__7919__CLK (.DIODE(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7919__RESET_B (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__7920__CLK (.DIODE(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7920__RESET_B (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__7921__CLK (.DIODE(\clknet_leaf_71_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7921__RESET_B (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__7922__CLK (.DIODE(\clknet_leaf_67_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7922__RESET_B (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__7923__CLK (.DIODE(\clknet_leaf_61_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7923__RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__7924__CLK (.DIODE(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7924__RESET_B (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__7925__CLK (.DIODE(\clknet_leaf_71_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7925__RESET_B (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA__7926__CLK (.DIODE(\clknet_leaf_61_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7926__RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__7927__CLK (.DIODE(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7927__RESET_B (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA__7928__CLK (.DIODE(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7928__RESET_B (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA__7929__CLK (.DIODE(\clknet_leaf_64_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7929__RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__7930__CLK (.DIODE(\clknet_leaf_71_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7930__RESET_B (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA__7931__CLK (.DIODE(\clknet_leaf_72_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7931__RESET_B (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA__7932__CLK (.DIODE(\clknet_leaf_71_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7932__RESET_B (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__7933__CLK (.DIODE(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7933__RESET_B (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA__7934__CLK (.DIODE(\clknet_leaf_60_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7934__RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__7935__CLK (.DIODE(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7935__RESET_B (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA__7936__CLK (.DIODE(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7936__RESET_B (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA__7937__CLK (.DIODE(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7937__RESET_B (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA__7938__CLK (.DIODE(\clknet_leaf_66_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7938__RESET_B (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__7939__CLK (.DIODE(\clknet_leaf_96_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7939__RESET_B (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__7940__CLK (.DIODE(\clknet_leaf_96_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7940__RESET_B (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__7941__CLK (.DIODE(\clknet_leaf_96_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7941__RESET_B (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA__7942__CLK (.DIODE(\clknet_leaf_96_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7942__RESET_B (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__7943__CLK (.DIODE(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7943__RESET_B (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA__7944__CLK (.DIODE(\clknet_leaf_96_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7944__RESET_B (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__7945__CLK (.DIODE(\clknet_leaf_95_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7945__RESET_B (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA__7946__CLK (.DIODE(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7947__CLK (.DIODE(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7948__CLK (.DIODE(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7949__CLK (.DIODE(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7950__CLK (.DIODE(\clknet_leaf_11_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7951__CLK (.DIODE(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7952__CLK (.DIODE(\clknet_leaf_99_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7953__CLK (.DIODE(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7954__CLK (.DIODE(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7955__CLK (.DIODE(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7956__CLK (.DIODE(\clknet_leaf_8_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7957__CLK (.DIODE(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7958__CLK (.DIODE(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7959__CLK (.DIODE(\clknet_leaf_63_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7960__CLK (.DIODE(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7961__CLK (.DIODE(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7962__CLK (.DIODE(\clknet_leaf_66_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7963__CLK (.DIODE(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7964__CLK (.DIODE(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7965__CLK (.DIODE(\clknet_leaf_67_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7966__CLK (.DIODE(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7967__CLK (.DIODE(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7968__CLK (.DIODE(\clknet_leaf_64_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7969__CLK (.DIODE(\clknet_leaf_41_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7970__CLK (.DIODE(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7971__CLK (.DIODE(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7972__CLK (.DIODE(\clknet_leaf_67_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7973__CLK (.DIODE(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7974__CLK (.DIODE(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7975__CLK (.DIODE(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7976__CLK (.DIODE(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7977__CLK (.DIODE(\clknet_leaf_67_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7978__CLK (.DIODE(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7979__CLK (.DIODE(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7980__CLK (.DIODE(\clknet_leaf_69_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7981__CLK (.DIODE(\clknet_leaf_66_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7982__CLK (.DIODE(\clknet_leaf_66_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7983__CLK (.DIODE(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7984__CLK (.DIODE(\clknet_leaf_66_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7985__CLK (.DIODE(\clknet_leaf_95_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7986__CLK (.DIODE(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7987__CLK (.DIODE(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7988__CLK (.DIODE(\clknet_leaf_69_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7989__CLK (.DIODE(\clknet_leaf_95_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7990__CLK (.DIODE(\clknet_leaf_95_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7991__CLK (.DIODE(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7992__CLK (.DIODE(\clknet_leaf_8_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7993__CLK (.DIODE(\clknet_leaf_8_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7994__CLK (.DIODE(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7995__CLK (.DIODE(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7996__CLK (.DIODE(\clknet_leaf_96_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7997__CLK (.DIODE(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7998__CLK (.DIODE(\clknet_leaf_8_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7999__CLK (.DIODE(\clknet_leaf_0_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7999__RESET_B (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__8000__CLK (.DIODE(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8000__RESET_B (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__8001__CLK (.DIODE(\clknet_leaf_12_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8001__RESET_B (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA__8002__CLK (.DIODE(\clknet_leaf_12_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8002__RESET_B (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA__8003__CLK (.DIODE(\clknet_leaf_34_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8003__RESET_B (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA__8004__CLK (.DIODE(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8004__D (.DIODE(_0484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8004__RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA__8005__CLK (.DIODE(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8005__D (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA__8005__RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA__8006__CLK (.DIODE(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8006__D (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__8006__RESET_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA__8007__CLK (.DIODE(\clknet_leaf_49_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8007__RESET_B (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA__8008__CLK (.DIODE(\clknet_leaf_47_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8008__RESET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA__8009__CLK (.DIODE(\clknet_leaf_46_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8009__RESET_B (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA__8010__CLK (.DIODE(\clknet_leaf_30_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8010__RESET_B (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__8011__CLK (.DIODE(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8011__RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA__8012__CLK (.DIODE(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8012__RESET_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA__8013__CLK (.DIODE(\clknet_leaf_30_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8013__RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA__8014__CLK (.DIODE(\clknet_leaf_30_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8014__RESET_B (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__8015__CLK (.DIODE(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8015__RESET_B (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__8016__CLK (.DIODE(\clknet_leaf_30_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8016__RESET_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA__8017__CLK (.DIODE(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8018__CLK (.DIODE(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8019__CLK (.DIODE(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8020__CLK (.DIODE(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8021__CLK (.DIODE(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8022__CLK (.DIODE(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8023__CLK (.DIODE(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8024__CLK (.DIODE(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8025__CLK (.DIODE(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8026__CLK (.DIODE(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8027__CLK (.DIODE(\clknet_leaf_8_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8028__CLK (.DIODE(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8029__CLK (.DIODE(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8030__CLK (.DIODE(\clknet_leaf_41_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8031__CLK (.DIODE(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8032__CLK (.DIODE(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8033__CLK (.DIODE(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8034__CLK (.DIODE(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8035__CLK (.DIODE(\clknet_leaf_64_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8036__CLK (.DIODE(\clknet_leaf_67_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8037__CLK (.DIODE(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8038__CLK (.DIODE(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8039__CLK (.DIODE(\clknet_leaf_64_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8040__CLK (.DIODE(\clknet_leaf_41_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8041__CLK (.DIODE(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8042__CLK (.DIODE(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8043__CLK (.DIODE(\clknet_leaf_67_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8044__CLK (.DIODE(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8045__CLK (.DIODE(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8046__CLK (.DIODE(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8047__CLK (.DIODE(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8048__CLK (.DIODE(\clknet_leaf_67_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8049__CLK (.DIODE(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8050__CLK (.DIODE(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8051__CLK (.DIODE(\clknet_leaf_69_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8052__CLK (.DIODE(\clknet_leaf_67_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8053__CLK (.DIODE(\clknet_leaf_67_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8054__CLK (.DIODE(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8055__CLK (.DIODE(\clknet_leaf_66_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8056__CLK (.DIODE(\clknet_leaf_95_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8057__CLK (.DIODE(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8058__CLK (.DIODE(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8059__CLK (.DIODE(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8060__CLK (.DIODE(\clknet_leaf_95_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8061__CLK (.DIODE(\clknet_leaf_67_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8062__CLK (.DIODE(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8063__CLK (.DIODE(\clknet_leaf_96_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8064__CLK (.DIODE(\clknet_leaf_8_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8065__CLK (.DIODE(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8066__CLK (.DIODE(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8067__CLK (.DIODE(\clknet_leaf_96_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8068__CLK (.DIODE(\clknet_leaf_8_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8069__CLK (.DIODE(\clknet_leaf_97_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8070__CLK (.DIODE(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8071__CLK (.DIODE(\clknet_leaf_105_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8072__CLK (.DIODE(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8073__CLK (.DIODE(\clknet_leaf_97_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8074__CLK (.DIODE(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8075__CLK (.DIODE(\clknet_leaf_97_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8076__CLK (.DIODE(\clknet_leaf_97_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8077__CLK (.DIODE(\clknet_leaf_97_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8078__CLK (.DIODE(\clknet_leaf_98_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8079__CLK (.DIODE(\clknet_leaf_101_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8080__CLK (.DIODE(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8081__CLK (.DIODE(\clknet_leaf_90_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8082__CLK (.DIODE(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8083__CLK (.DIODE(\clknet_leaf_89_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8084__CLK (.DIODE(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8085__CLK (.DIODE(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8086__CLK (.DIODE(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8087__CLK (.DIODE(\clknet_leaf_93_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8088__CLK (.DIODE(\clknet_leaf_86_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8089__CLK (.DIODE(\clknet_leaf_93_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8090__CLK (.DIODE(\clknet_leaf_93_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8091__CLK (.DIODE(\clknet_leaf_86_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8092__CLK (.DIODE(\clknet_leaf_86_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8093__CLK (.DIODE(\clknet_leaf_69_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8094__CLK (.DIODE(\clknet_leaf_93_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8095__CLK (.DIODE(\clknet_leaf_69_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8096__CLK (.DIODE(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8097__CLK (.DIODE(\clknet_leaf_87_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8098__CLK (.DIODE(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8099__CLK (.DIODE(\clknet_leaf_92_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8100__CLK (.DIODE(\clknet_leaf_87_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8101__CLK (.DIODE(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8102__CLK (.DIODE(\clknet_leaf_89_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8103__CLK (.DIODE(\clknet_leaf_92_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8104__CLK (.DIODE(\clknet_leaf_87_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8105__CLK (.DIODE(\clknet_leaf_92_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8106__CLK (.DIODE(\clknet_leaf_87_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8107__CLK (.DIODE(\clknet_leaf_91_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8108__CLK (.DIODE(\clknet_leaf_92_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8109__CLK (.DIODE(\clknet_leaf_91_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8110__CLK (.DIODE(\clknet_leaf_90_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8111__CLK (.DIODE(\clknet_leaf_101_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8112__CLK (.DIODE(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8113__CLK (.DIODE(\clknet_leaf_86_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8114__CLK (.DIODE(\clknet_leaf_91_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8115__CLK (.DIODE(\clknet_leaf_90_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8116__CLK (.DIODE(\clknet_leaf_91_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8117__CLK (.DIODE(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8118__CLK (.DIODE(\clknet_leaf_106_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8119__CLK (.DIODE(\clknet_leaf_101_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8120__CLK (.DIODE(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8121__CLK (.DIODE(\clknet_leaf_90_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8122__CLK (.DIODE(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8123__CLK (.DIODE(\clknet_leaf_101_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8124__CLK (.DIODE(\clknet_leaf_105_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8125__CLK (.DIODE(\clknet_leaf_106_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8126__CLK (.DIODE(\clknet_leaf_107_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8127__CLK (.DIODE(\clknet_leaf_107_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8128__CLK (.DIODE(\clknet_leaf_107_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8129__CLK (.DIODE(\clknet_leaf_108_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8130__CLK (.DIODE(\clknet_leaf_107_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8131__CLK (.DIODE(\clknet_leaf_102_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8132__CLK (.DIODE(\clknet_leaf_102_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8133__CLK (.DIODE(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8134__CLK (.DIODE(\clknet_leaf_90_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8135__CLK (.DIODE(\clknet_leaf_106_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8136__CLK (.DIODE(\clknet_leaf_102_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8137__CLK (.DIODE(\clknet_leaf_102_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8138__CLK (.DIODE(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8139__CLK (.DIODE(\clknet_leaf_104_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8140__CLK (.DIODE(\clknet_leaf_104_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8141__CLK (.DIODE(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8142__CLK (.DIODE(\clknet_leaf_104_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8143__CLK (.DIODE(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8144__CLK (.DIODE(\clknet_leaf_105_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8145__CLK (.DIODE(\clknet_leaf_105_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8146__CLK (.DIODE(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8147__CLK (.DIODE(\clknet_leaf_48_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8147__RESET_B (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA__8148__CLK (.DIODE(\clknet_leaf_47_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8148__RESET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA__8149__CLK (.DIODE(\clknet_leaf_46_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8149__RESET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA__8150__CLK (.DIODE(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8151__CLK (.DIODE(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8152__CLK (.DIODE(\clknet_leaf_75_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8153__CLK (.DIODE(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8154__CLK (.DIODE(\clknet_leaf_75_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8155__CLK (.DIODE(\clknet_leaf_75_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8156__CLK (.DIODE(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8157__CLK (.DIODE(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8158__CLK (.DIODE(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8159__CLK (.DIODE(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8160__CLK (.DIODE(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8161__CLK (.DIODE(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8162__CLK (.DIODE(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8163__CLK (.DIODE(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8164__CLK (.DIODE(\clknet_leaf_81_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8165__CLK (.DIODE(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8166__CLK (.DIODE(\clknet_leaf_82_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8167__CLK (.DIODE(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8168__CLK (.DIODE(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8169__CLK (.DIODE(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8170__CLK (.DIODE(\clknet_leaf_81_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8171__CLK (.DIODE(\clknet_leaf_77_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8172__CLK (.DIODE(\clknet_leaf_82_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8173__CLK (.DIODE(\clknet_leaf_85_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8174__CLK (.DIODE(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8175__CLK (.DIODE(\clknet_leaf_85_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8176__CLK (.DIODE(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8177__CLK (.DIODE(\clknet_leaf_82_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8178__CLK (.DIODE(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8179__CLK (.DIODE(\clknet_leaf_81_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8180__CLK (.DIODE(\clknet_leaf_83_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8181__CLK (.DIODE(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8182__CLK (.DIODE(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8183__CLK (.DIODE(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8184__CLK (.DIODE(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8185__CLK (.DIODE(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8186__CLK (.DIODE(\clknet_leaf_75_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8187__CLK (.DIODE(\clknet_leaf_75_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8188__CLK (.DIODE(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8189__CLK (.DIODE(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8190__CLK (.DIODE(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8191__CLK (.DIODE(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8192__CLK (.DIODE(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8193__CLK (.DIODE(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8194__CLK (.DIODE(\clknet_leaf_81_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8195__CLK (.DIODE(\clknet_leaf_85_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8196__CLK (.DIODE(\clknet_leaf_81_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8197__CLK (.DIODE(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8198__CLK (.DIODE(\clknet_leaf_81_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8199__CLK (.DIODE(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8200__CLK (.DIODE(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8201__CLK (.DIODE(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8202__CLK (.DIODE(\clknet_leaf_81_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8203__CLK (.DIODE(\clknet_leaf_71_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8204__CLK (.DIODE(\clknet_leaf_82_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8205__CLK (.DIODE(\clknet_leaf_85_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8206__CLK (.DIODE(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8207__CLK (.DIODE(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8208__CLK (.DIODE(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8209__CLK (.DIODE(\clknet_leaf_82_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8210__CLK (.DIODE(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8211__CLK (.DIODE(\clknet_leaf_81_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8212__CLK (.DIODE(\clknet_leaf_82_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8213__CLK (.DIODE(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8214__CLK (.DIODE(\clknet_leaf_85_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8215__CLK (.DIODE(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8216__CLK (.DIODE(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8217__CLK (.DIODE(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8218__CLK (.DIODE(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8219__CLK (.DIODE(\clknet_leaf_75_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8220__CLK (.DIODE(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8221__CLK (.DIODE(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8222__CLK (.DIODE(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8223__CLK (.DIODE(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8224__CLK (.DIODE(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8225__CLK (.DIODE(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8226__CLK (.DIODE(\clknet_leaf_81_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8227__CLK (.DIODE(\clknet_leaf_85_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8228__CLK (.DIODE(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8229__CLK (.DIODE(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8230__CLK (.DIODE(\clknet_leaf_82_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8231__CLK (.DIODE(\clknet_leaf_77_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8232__CLK (.DIODE(\clknet_leaf_77_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8233__CLK (.DIODE(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8234__CLK (.DIODE(\clknet_leaf_81_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8235__CLK (.DIODE(\clknet_leaf_71_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8236__CLK (.DIODE(\clknet_leaf_82_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8237__CLK (.DIODE(\clknet_leaf_84_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8238__CLK (.DIODE(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8239__CLK (.DIODE(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8240__CLK (.DIODE(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8241__CLK (.DIODE(\clknet_leaf_85_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8242__CLK (.DIODE(\clknet_leaf_82_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8243__CLK (.DIODE(\clknet_leaf_81_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8244__CLK (.DIODE(\clknet_leaf_83_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8245__CLK (.DIODE(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8246__CLK (.DIODE(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8247__CLK (.DIODE(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8248__CLK (.DIODE(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8249__CLK (.DIODE(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8250__CLK (.DIODE(\clknet_leaf_75_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8251__CLK (.DIODE(\clknet_leaf_75_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8252__CLK (.DIODE(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8253__CLK (.DIODE(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8254__CLK (.DIODE(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8255__CLK (.DIODE(\clknet_leaf_77_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8256__CLK (.DIODE(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8257__CLK (.DIODE(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8258__CLK (.DIODE(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8259__CLK (.DIODE(\clknet_leaf_85_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8260__CLK (.DIODE(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8261__CLK (.DIODE(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8262__CLK (.DIODE(\clknet_leaf_82_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8263__CLK (.DIODE(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8264__CLK (.DIODE(\clknet_leaf_77_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8265__CLK (.DIODE(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8266__CLK (.DIODE(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8267__CLK (.DIODE(\clknet_leaf_71_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8268__CLK (.DIODE(\clknet_leaf_82_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8269__CLK (.DIODE(\clknet_leaf_84_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8270__CLK (.DIODE(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8271__CLK (.DIODE(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8272__CLK (.DIODE(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8273__CLK (.DIODE(\clknet_leaf_83_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8274__CLK (.DIODE(\clknet_leaf_82_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8275__CLK (.DIODE(\clknet_leaf_81_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8276__CLK (.DIODE(\clknet_leaf_83_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8277__CLK (.DIODE(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8278__CLK (.DIODE(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8279__CLK (.DIODE(\clknet_leaf_30_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8280__CLK (.DIODE(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8281__CLK (.DIODE(\clknet_leaf_29_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8282__CLK (.DIODE(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8283__CLK (.DIODE(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8284__CLK (.DIODE(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8285__CLK (.DIODE(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8286__CLK (.DIODE(\clknet_leaf_27_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8287__CLK (.DIODE(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8288__CLK (.DIODE(\clknet_leaf_30_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8289__CLK (.DIODE(\clknet_leaf_32_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8290__CLK (.DIODE(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8291__CLK (.DIODE(\clknet_leaf_43_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8292__CLK (.DIODE(\clknet_leaf_43_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8293__CLK (.DIODE(\clknet_leaf_45_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8294__CLK (.DIODE(\clknet_leaf_43_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8295__CLK (.DIODE(\clknet_leaf_48_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8296__CLK (.DIODE(\clknet_leaf_43_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8297__CLK (.DIODE(\clknet_leaf_43_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8298__CLK (.DIODE(\clknet_leaf_46_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8299__CLK (.DIODE(\clknet_leaf_41_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8300__CLK (.DIODE(\clknet_leaf_44_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8301__CLK (.DIODE(\clknet_leaf_47_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8302__CLK (.DIODE(\clknet_leaf_40_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8303__CLK (.DIODE(\clknet_leaf_44_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8304__CLK (.DIODE(\clknet_leaf_40_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8305__CLK (.DIODE(\clknet_leaf_45_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8306__CLK (.DIODE(\clknet_leaf_43_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8307__CLK (.DIODE(\clknet_leaf_45_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8308__CLK (.DIODE(\clknet_leaf_32_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8309__CLK (.DIODE(\clknet_leaf_45_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8310__CLK (.DIODE(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8311__CLK (.DIODE(\clknet_leaf_40_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8312__CLK (.DIODE(\clknet_leaf_41_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8313__CLK (.DIODE(\clknet_leaf_44_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8314__CLK (.DIODE(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8315__CLK (.DIODE(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8316__CLK (.DIODE(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8317__CLK (.DIODE(\clknet_leaf_46_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8318__CLK (.DIODE(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8319__CLK (.DIODE(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8320__CLK (.DIODE(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8321__CLK (.DIODE(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8322__CLK (.DIODE(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8323__CLK (.DIODE(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8324__CLK (.DIODE(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8325__CLK (.DIODE(\clknet_leaf_27_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8326__CLK (.DIODE(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8327__CLK (.DIODE(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8328__CLK (.DIODE(\clknet_leaf_34_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8329__CLK (.DIODE(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8330__CLK (.DIODE(\clknet_leaf_34_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8331__CLK (.DIODE(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8332__CLK (.DIODE(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8333__CLK (.DIODE(\clknet_leaf_86_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8333__RESET_B (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA__8334__CLK (.DIODE(\clknet_leaf_83_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8334__RESET_B (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__8335__CLK (.DIODE(\clknet_leaf_84_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8335__RESET_B (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__8336__CLK (.DIODE(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8336__RESET_B (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA__8337__CLK (.DIODE(\clknet_leaf_87_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8337__RESET_B (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__8338__CLK (.DIODE(\clknet_leaf_77_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8338__RESET_B (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA__8339__CLK (.DIODE(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8339__RESET_B (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__8340__CLK (.DIODE(\clknet_leaf_71_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8340__RESET_B (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA__8341__CLK (.DIODE(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8341__RESET_B (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA__8342__CLK (.DIODE(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8342__RESET_B (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA__8343__CLK (.DIODE(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8343__RESET_B (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA__8344__CLK (.DIODE(\clknet_leaf_89_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8344__RESET_B (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__8345__CLK (.DIODE(\clknet_leaf_83_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8345__RESET_B (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__8346__CLK (.DIODE(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8347__CLK (.DIODE(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8347__RESET_B (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__8348__CLK (.DIODE(\clknet_leaf_77_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8348__RESET_B (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__8349__CLK (.DIODE(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8349__RESET_B (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA__8350__CLK (.DIODE(\clknet_leaf_93_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8350__RESET_B (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__8351__CLK (.DIODE(\clknet_leaf_86_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8351__RESET_B (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA__8352__CLK (.DIODE(\clknet_leaf_86_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8352__RESET_B (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA__8353__CLK (.DIODE(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8353__RESET_B (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA__8354__CLK (.DIODE(\clknet_leaf_84_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8354__RESET_B (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__8355__CLK (.DIODE(\clknet_leaf_85_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8355__RESET_B (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA__8356__CLK (.DIODE(\clknet_leaf_69_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8356__RESET_B (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA__8357__CLK (.DIODE(\clknet_leaf_85_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8357__RESET_B (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA__8358__CLK (.DIODE(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8358__RESET_B (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA__8359__CLK (.DIODE(\clknet_leaf_87_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8359__RESET_B (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__8360__CLK (.DIODE(\clknet_leaf_84_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8360__RESET_B (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__8361__CLK (.DIODE(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8361__RESET_B (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA__8362__CLK (.DIODE(\clknet_leaf_85_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8362__RESET_B (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA__8363__CLK (.DIODE(\clknet_leaf_87_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8363__RESET_B (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__8364__CLK (.DIODE(\clknet_leaf_85_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8364__RESET_B (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA__8365__CLK (.DIODE(\clknet_leaf_87_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8365__RESET_B (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA__8366__CLK (.DIODE(\clknet_leaf_86_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8366__RESET_B (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA__8367__CLK (.DIODE(\clknet_leaf_84_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8367__RESET_B (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__8368__CLK (.DIODE(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8368__RESET_B (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA__8369__CLK (.DIODE(\clknet_leaf_87_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8369__RESET_B (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA__8370__CLK (.DIODE(\clknet_leaf_84_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8370__RESET_B (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__8371__CLK (.DIODE(\clknet_leaf_87_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8371__RESET_B (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA__8372__CLK (.DIODE(\clknet_leaf_86_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8372__RESET_B (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA__8373__CLK (.DIODE(\clknet_leaf_92_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8373__RESET_B (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA__8374__CLK (.DIODE(\clknet_leaf_85_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8374__RESET_B (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA__8375__CLK (.DIODE(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8375__RESET_B (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__8376__CLK (.DIODE(\clknet_leaf_85_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8376__RESET_B (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__8377__CLK (.DIODE(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8377__RESET_B (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA__8378__CLK (.DIODE(\clknet_leaf_84_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8378__RESET_B (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__8379__CLK (.DIODE(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8379__RESET_B (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__8380__CLK (.DIODE(\clknet_leaf_84_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8380__RESET_B (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__8381__CLK (.DIODE(\clknet_leaf_85_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8381__RESET_B (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA__8382__CLK (.DIODE(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8382__RESET_B (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA__8383__CLK (.DIODE(\clknet_leaf_85_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8383__RESET_B (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA__8384__CLK (.DIODE(\clknet_leaf_89_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8384__RESET_B (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__8385__CLK (.DIODE(\clknet_leaf_84_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8386__CLK (.DIODE(\clknet_leaf_85_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8386__RESET_B (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA__8387__CLK (.DIODE(\clknet_leaf_83_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8387__RESET_B (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__8388__CLK (.DIODE(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8389__CLK (.DIODE(\clknet_leaf_82_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8390__CLK (.DIODE(\clknet_leaf_83_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8390__RESET_B (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__8391__CLK (.DIODE(\clknet_leaf_85_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8391__RESET_B (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA__8392__CLK (.DIODE(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8392__RESET_B (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__8393__CLK (.DIODE(\clknet_leaf_83_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8394__CLK (.DIODE(\clknet_leaf_89_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8394__RESET_B (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__8395__CLK (.DIODE(\clknet_leaf_89_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8395__RESET_B (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__8396__CLK (.DIODE(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8396__RESET_B (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__8397__CLK (.DIODE(\clknet_leaf_83_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8398__CLK (.DIODE(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8398__RESET_B (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__8399__CLK (.DIODE(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8399__RESET_B (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__8400__CLK (.DIODE(\clknet_leaf_84_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8400__RESET_B (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA__8401__CLK (.DIODE(\clknet_leaf_83_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8402__CLK (.DIODE(\clknet_leaf_84_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8402__RESET_B (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__8403__CLK (.DIODE(\clknet_leaf_83_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8404__CLK (.DIODE(\clknet_leaf_83_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8405__CLK (.DIODE(\clknet_leaf_83_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8406__CLK (.DIODE(\clknet_leaf_84_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8407__CLK (.DIODE(\clknet_leaf_83_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8408__CLK (.DIODE(\clknet_leaf_84_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8409__CLK (.DIODE(\clknet_leaf_83_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8410__CLK (.DIODE(\clknet_leaf_11_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8410__SET_B (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA__8411__CLK (.DIODE(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8411__RESET_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__8412__CLK (.DIODE(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8412__RESET_B (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__8413__CLK (.DIODE(\clknet_leaf_58_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8414__CLK (.DIODE(\clknet_leaf_62_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8415__CLK (.DIODE(\clknet_leaf_57_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8416__CLK (.DIODE(\clknet_leaf_73_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8417__CLK (.DIODE(\clknet_leaf_60_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8418__CLK (.DIODE(\clknet_leaf_56_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8419__CLK (.DIODE(\clknet_leaf_56_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8420__CLK (.DIODE(\clknet_leaf_60_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8421__CLK (.DIODE(\clknet_leaf_58_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8422__CLK (.DIODE(\clknet_leaf_59_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8423__CLK (.DIODE(\clknet_leaf_75_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8424__CLK (.DIODE(\clknet_leaf_74_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8425__CLK (.DIODE(\clknet_leaf_59_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8426__CLK (.DIODE(\clknet_leaf_72_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8427__CLK (.DIODE(\clknet_leaf_59_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8428__CLK (.DIODE(\clknet_leaf_59_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8429__CLK (.DIODE(\clknet_leaf_59_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8430__CLK (.DIODE(\clknet_leaf_71_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8431__CLK (.DIODE(\clknet_leaf_58_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8432__CLK (.DIODE(\clknet_leaf_77_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8433__CLK (.DIODE(\clknet_leaf_73_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8434__CLK (.DIODE(\clknet_leaf_59_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8435__CLK (.DIODE(\clknet_leaf_73_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8436__CLK (.DIODE(\clknet_leaf_74_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8437__CLK (.DIODE(\clknet_leaf_74_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8438__CLK (.DIODE(\clknet_leaf_73_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8439__CLK (.DIODE(\clknet_leaf_75_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8440__CLK (.DIODE(\clknet_leaf_71_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8441__CLK (.DIODE(\clknet_leaf_71_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8442__CLK (.DIODE(\clknet_leaf_73_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8443__CLK (.DIODE(\clknet_leaf_71_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8444__CLK (.DIODE(\clknet_leaf_72_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8445__CLK (.DIODE(\clknet_leaf_59_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8446__CLK (.DIODE(\clknet_leaf_61_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8447__CLK (.DIODE(\clknet_leaf_56_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8448__CLK (.DIODE(\clknet_leaf_74_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8449__CLK (.DIODE(\clknet_leaf_60_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8450__CLK (.DIODE(\clknet_leaf_62_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8451__CLK (.DIODE(\clknet_leaf_56_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8452__CLK (.DIODE(\clknet_leaf_60_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8453__CLK (.DIODE(\clknet_leaf_57_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8454__CLK (.DIODE(\clknet_leaf_59_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8455__CLK (.DIODE(\clknet_leaf_74_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8456__CLK (.DIODE(\clknet_leaf_73_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8457__CLK (.DIODE(\clknet_leaf_60_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8458__CLK (.DIODE(\clknet_leaf_72_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8459__CLK (.DIODE(\clknet_leaf_59_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8460__CLK (.DIODE(\clknet_leaf_60_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8461__CLK (.DIODE(\clknet_leaf_60_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8462__CLK (.DIODE(\clknet_leaf_72_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8463__CLK (.DIODE(\clknet_leaf_60_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8464__CLK (.DIODE(\clknet_leaf_71_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8465__CLK (.DIODE(\clknet_leaf_72_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8466__CLK (.DIODE(\clknet_leaf_74_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8467__CLK (.DIODE(\clknet_leaf_75_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8468__CLK (.DIODE(\clknet_leaf_73_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8469__CLK (.DIODE(\clknet_leaf_75_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8470__CLK (.DIODE(\clknet_leaf_73_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8471__CLK (.DIODE(\clknet_leaf_75_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8472__CLK (.DIODE(\clknet_leaf_71_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8473__CLK (.DIODE(\clknet_leaf_71_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8474__CLK (.DIODE(\clknet_leaf_73_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8475__CLK (.DIODE(\clknet_leaf_71_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8476__CLK (.DIODE(\clknet_leaf_72_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8477__CLK (.DIODE(\clknet_leaf_58_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8478__CLK (.DIODE(\clknet_leaf_61_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8479__CLK (.DIODE(\clknet_leaf_60_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8480__CLK (.DIODE(\clknet_leaf_74_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8481__CLK (.DIODE(\clknet_leaf_60_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8482__CLK (.DIODE(\clknet_leaf_58_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8483__CLK (.DIODE(\clknet_leaf_56_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8484__CLK (.DIODE(\clknet_leaf_60_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8485__CLK (.DIODE(\clknet_leaf_58_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8486__CLK (.DIODE(\clknet_leaf_59_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8487__CLK (.DIODE(\clknet_leaf_75_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8488__CLK (.DIODE(\clknet_leaf_74_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8489__CLK (.DIODE(\clknet_leaf_60_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8490__CLK (.DIODE(\clknet_leaf_72_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8491__CLK (.DIODE(\clknet_leaf_59_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8492__CLK (.DIODE(\clknet_leaf_59_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8493__CLK (.DIODE(\clknet_leaf_59_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8494__CLK (.DIODE(\clknet_leaf_71_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8495__CLK (.DIODE(\clknet_leaf_58_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8496__CLK (.DIODE(\clknet_leaf_75_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8497__CLK (.DIODE(\clknet_leaf_73_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8498__CLK (.DIODE(\clknet_leaf_74_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8499__CLK (.DIODE(\clknet_leaf_74_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8500__CLK (.DIODE(\clknet_leaf_74_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8501__CLK (.DIODE(\clknet_leaf_74_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8502__CLK (.DIODE(\clknet_leaf_73_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8503__CLK (.DIODE(\clknet_leaf_75_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8504__CLK (.DIODE(\clknet_leaf_72_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8505__CLK (.DIODE(\clknet_leaf_72_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8506__CLK (.DIODE(\clknet_leaf_73_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8507__CLK (.DIODE(\clknet_leaf_71_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8508__CLK (.DIODE(\clknet_leaf_72_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8509__CLK (.DIODE(\clknet_leaf_58_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8510__CLK (.DIODE(\clknet_leaf_60_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8511__CLK (.DIODE(\clknet_leaf_57_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8512__CLK (.DIODE(\clknet_leaf_74_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8513__CLK (.DIODE(\clknet_leaf_59_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8514__CLK (.DIODE(\clknet_leaf_58_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8515__CLK (.DIODE(\clknet_leaf_57_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8516__CLK (.DIODE(\clknet_leaf_60_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8517__CLK (.DIODE(\clknet_leaf_58_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8518__CLK (.DIODE(\clknet_leaf_59_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8519__CLK (.DIODE(\clknet_leaf_75_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8520__CLK (.DIODE(\clknet_leaf_74_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8521__CLK (.DIODE(\clknet_leaf_59_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8522__CLK (.DIODE(\clknet_leaf_72_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8523__CLK (.DIODE(\clknet_leaf_59_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8524__CLK (.DIODE(\clknet_leaf_60_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8525__CLK (.DIODE(\clknet_leaf_59_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8526__CLK (.DIODE(\clknet_leaf_72_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8527__CLK (.DIODE(\clknet_leaf_58_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8528__CLK (.DIODE(\clknet_leaf_74_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8529__CLK (.DIODE(\clknet_leaf_73_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8530__CLK (.DIODE(\clknet_leaf_74_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8531__CLK (.DIODE(\clknet_leaf_74_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8532__CLK (.DIODE(\clknet_leaf_74_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8533__CLK (.DIODE(\clknet_leaf_75_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8534__CLK (.DIODE(\clknet_leaf_73_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8535__CLK (.DIODE(\clknet_leaf_75_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8536__CLK (.DIODE(\clknet_leaf_73_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8537__CLK (.DIODE(\clknet_leaf_72_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8538__CLK (.DIODE(\clknet_leaf_74_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8539__CLK (.DIODE(\clknet_leaf_72_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8540__CLK (.DIODE(\clknet_leaf_73_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8541__CLK (.DIODE(\clknet_leaf_107_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8541__RESET_B (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__8542__CLK (.DIODE(\clknet_leaf_109_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8542__RESET_B (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__8543__CLK (.DIODE(\clknet_leaf_14_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8543__RESET_B (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA__8544__CLK (.DIODE(\clknet_leaf_14_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8544__RESET_B (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA__8545__CLK (.DIODE(\clknet_leaf_11_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8545__RESET_B (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__8546__CLK (.DIODE(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8546__RESET_B (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__8547__CLK (.DIODE(\clknet_leaf_27_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8547__RESET_B (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA__8548__CLK (.DIODE(\clknet_leaf_26_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8548__RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA__8549__CLK (.DIODE(\clknet_leaf_27_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8549__RESET_B (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA__8550__CLK (.DIODE(\clknet_leaf_34_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8550__RESET_B (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA__8551__CLK (.DIODE(\clknet_leaf_34_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8551__RESET_B (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA__8552__CLK (.DIODE(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8552__RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA__8553__CLK (.DIODE(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8553__RESET_B (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA__8554__CLK (.DIODE(\clknet_leaf_27_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8554__RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA__8555__CLK (.DIODE(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8555__RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA__8556__CLK (.DIODE(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8556__RESET_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA__8557__CLK (.DIODE(\clknet_leaf_8_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8557__D (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__8557__RESET_B (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA__8558__CLK (.DIODE(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8558__D (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__8558__RESET_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__8559__CLK (.DIODE(\clknet_leaf_61_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8559__RESET_B (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__8560__CLK (.DIODE(\clknet_leaf_72_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8560__RESET_B (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA__8561__CLK (.DIODE(\clknet_leaf_61_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8561__RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__8562__CLK (.DIODE(\clknet_leaf_11_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8562__RESET_B (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__8563__CLK (.DIODE(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8563__RESET_B (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__8564__CLK (.DIODE(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8564__RESET_B (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__8565__CLK (.DIODE(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8566__CLK (.DIODE(\clknet_leaf_32_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8567__CLK (.DIODE(\clknet_leaf_29_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8568__CLK (.DIODE(\clknet_leaf_29_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8569__CLK (.DIODE(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8570__CLK (.DIODE(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8571__CLK (.DIODE(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8572__CLK (.DIODE(\clknet_leaf_34_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8573__CLK (.DIODE(\clknet_leaf_34_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8574__CLK (.DIODE(\clknet_leaf_45_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8575__CLK (.DIODE(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8576__CLK (.DIODE(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8577__CLK (.DIODE(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8578__CLK (.DIODE(\clknet_leaf_42_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8579__CLK (.DIODE(\clknet_leaf_42_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8580__CLK (.DIODE(\clknet_leaf_46_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8581__CLK (.DIODE(\clknet_leaf_49_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8582__CLK (.DIODE(\clknet_leaf_47_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8583__CLK (.DIODE(\clknet_leaf_40_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8584__CLK (.DIODE(\clknet_leaf_41_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8585__CLK (.DIODE(\clknet_leaf_46_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8586__CLK (.DIODE(\clknet_leaf_41_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8587__CLK (.DIODE(\clknet_leaf_43_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8588__CLK (.DIODE(\clknet_leaf_47_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8589__CLK (.DIODE(\clknet_leaf_40_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8590__CLK (.DIODE(\clknet_leaf_44_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8591__CLK (.DIODE(\clknet_leaf_40_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8592__CLK (.DIODE(\clknet_leaf_47_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8593__CLK (.DIODE(\clknet_leaf_43_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8594__CLK (.DIODE(\clknet_leaf_45_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8595__CLK (.DIODE(\clknet_leaf_44_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8596__CLK (.DIODE(\clknet_leaf_46_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8597__CLK (.DIODE(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8598__CLK (.DIODE(\clknet_leaf_40_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8599__CLK (.DIODE(\clknet_leaf_41_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8600__CLK (.DIODE(\clknet_leaf_40_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8601__CLK (.DIODE(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8602__CLK (.DIODE(\clknet_leaf_40_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8603__CLK (.DIODE(\clknet_leaf_44_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8604__CLK (.DIODE(\clknet_leaf_46_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8605__CLK (.DIODE(\clknet_leaf_32_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8606__CLK (.DIODE(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8607__CLK (.DIODE(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8608__CLK (.DIODE(\clknet_leaf_32_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8609__CLK (.DIODE(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8610__CLK (.DIODE(\clknet_leaf_32_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8611__CLK (.DIODE(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8612__CLK (.DIODE(\clknet_leaf_34_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8613__CLK (.DIODE(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8614__CLK (.DIODE(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8615__CLK (.DIODE(\clknet_leaf_34_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8616__CLK (.DIODE(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8617__CLK (.DIODE(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8618__CLK (.DIODE(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8619__CLK (.DIODE(\clknet_leaf_11_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8620__CLK (.DIODE(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8620__RESET_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__8621__CLK (.DIODE(\clknet_leaf_67_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8621__RESET_B (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__8622__CLK (.DIODE(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8622__RESET_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__8623__CLK (.DIODE(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8623__RESET_B (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA__8624__CLK (.DIODE(\clknet_leaf_64_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8624__RESET_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__8625__CLK (.DIODE(\clknet_leaf_64_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8625__RESET_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__8626__CLK (.DIODE(\clknet_leaf_61_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8626__RESET_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__8627__CLK (.DIODE(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8628__CLK (.DIODE(\clknet_leaf_105_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8629__CLK (.DIODE(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8630__CLK (.DIODE(\clknet_leaf_97_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8631__CLK (.DIODE(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8632__CLK (.DIODE(\clknet_leaf_98_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8633__CLK (.DIODE(\clknet_leaf_98_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8634__CLK (.DIODE(\clknet_leaf_97_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8635__CLK (.DIODE(\clknet_leaf_97_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8636__CLK (.DIODE(\clknet_leaf_98_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8637__CLK (.DIODE(\clknet_leaf_106_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8638__CLK (.DIODE(\clknet_leaf_102_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8639__CLK (.DIODE(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8640__CLK (.DIODE(\clknet_leaf_90_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8641__CLK (.DIODE(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8642__CLK (.DIODE(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8643__CLK (.DIODE(\clknet_leaf_69_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8644__CLK (.DIODE(\clknet_leaf_93_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8645__CLK (.DIODE(\clknet_leaf_92_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8646__CLK (.DIODE(\clknet_leaf_93_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8647__CLK (.DIODE(\clknet_leaf_93_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8648__CLK (.DIODE(\clknet_leaf_86_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8649__CLK (.DIODE(\clknet_leaf_93_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8650__CLK (.DIODE(\clknet_leaf_93_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8651__CLK (.DIODE(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8652__CLK (.DIODE(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8653__CLK (.DIODE(\clknet_leaf_89_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8654__CLK (.DIODE(\clknet_leaf_87_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8655__CLK (.DIODE(\clknet_leaf_95_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8656__CLK (.DIODE(\clknet_leaf_92_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8657__CLK (.DIODE(\clknet_leaf_87_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8658__CLK (.DIODE(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8659__CLK (.DIODE(\clknet_leaf_89_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8660__CLK (.DIODE(\clknet_leaf_91_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8661__CLK (.DIODE(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8662__CLK (.DIODE(\clknet_leaf_92_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8663__CLK (.DIODE(\clknet_leaf_89_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8664__CLK (.DIODE(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8665__CLK (.DIODE(\clknet_leaf_91_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8666__CLK (.DIODE(\clknet_leaf_91_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8667__CLK (.DIODE(\clknet_leaf_90_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8668__CLK (.DIODE(\clknet_leaf_101_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8669__CLK (.DIODE(\clknet_leaf_89_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8670__CLK (.DIODE(\clknet_leaf_92_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8671__CLK (.DIODE(\clknet_leaf_91_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8672__CLK (.DIODE(\clknet_leaf_90_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8673__CLK (.DIODE(\clknet_leaf_101_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8674__CLK (.DIODE(\clknet_leaf_106_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8675__CLK (.DIODE(\clknet_leaf_106_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8676__CLK (.DIODE(\clknet_leaf_101_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8677__CLK (.DIODE(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8678__CLK (.DIODE(\clknet_leaf_102_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8679__CLK (.DIODE(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8680__CLK (.DIODE(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8681__CLK (.DIODE(\clknet_leaf_105_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8682__CLK (.DIODE(\clknet_leaf_106_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8683__CLK (.DIODE(\clknet_leaf_107_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8684__CLK (.DIODE(\clknet_leaf_107_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8685__CLK (.DIODE(\clknet_leaf_107_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8686__CLK (.DIODE(\clknet_leaf_108_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8687__CLK (.DIODE(\clknet_leaf_108_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8688__CLK (.DIODE(\clknet_leaf_102_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8689__CLK (.DIODE(\clknet_leaf_102_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8690__CLK (.DIODE(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8691__CLK (.DIODE(\clknet_leaf_90_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8692__CLK (.DIODE(\clknet_leaf_105_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8693__CLK (.DIODE(\clknet_leaf_104_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8694__CLK (.DIODE(\clknet_leaf_104_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8695__CLK (.DIODE(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8696__CLK (.DIODE(\clknet_leaf_104_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8697__CLK (.DIODE(\clknet_leaf_104_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8698__CLK (.DIODE(\clknet_leaf_104_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8699__CLK (.DIODE(\clknet_leaf_104_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8700__CLK (.DIODE(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8701__CLK (.DIODE(\clknet_leaf_105_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8702__CLK (.DIODE(\clknet_leaf_108_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8703__CLK (.DIODE(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8704__CLK (.DIODE(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8705__CLK (.DIODE(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8706__CLK (.DIODE(\clknet_leaf_29_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8707__CLK (.DIODE(\clknet_leaf_25_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8708__CLK (.DIODE(\clknet_leaf_11_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8709__CLK (.DIODE(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8710__CLK (.DIODE(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8711__CLK (.DIODE(\clknet_leaf_34_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8712__CLK (.DIODE(\clknet_leaf_27_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8713__CLK (.DIODE(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8714__CLK (.DIODE(\clknet_leaf_30_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8715__CLK (.DIODE(\clknet_leaf_32_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8716__CLK (.DIODE(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8717__CLK (.DIODE(\clknet_leaf_43_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8718__CLK (.DIODE(\clknet_leaf_40_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8719__CLK (.DIODE(\clknet_leaf_46_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8720__CLK (.DIODE(\clknet_leaf_42_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8721__CLK (.DIODE(\clknet_leaf_46_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8722__CLK (.DIODE(\clknet_leaf_40_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8723__CLK (.DIODE(\clknet_leaf_43_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8724__CLK (.DIODE(\clknet_leaf_46_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8725__CLK (.DIODE(\clknet_leaf_41_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8726__CLK (.DIODE(\clknet_leaf_44_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8727__CLK (.DIODE(\clknet_leaf_45_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8728__CLK (.DIODE(\clknet_leaf_40_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8729__CLK (.DIODE(\clknet_leaf_44_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8730__CLK (.DIODE(\clknet_leaf_40_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8731__CLK (.DIODE(\clknet_leaf_44_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8732__CLK (.DIODE(\clknet_leaf_44_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8733__CLK (.DIODE(\clknet_leaf_45_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8734__CLK (.DIODE(\clknet_leaf_32_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8735__CLK (.DIODE(\clknet_leaf_45_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8736__CLK (.DIODE(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8737__CLK (.DIODE(\clknet_leaf_40_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8738__CLK (.DIODE(\clknet_leaf_41_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8739__CLK (.DIODE(\clknet_leaf_44_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8740__CLK (.DIODE(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8741__CLK (.DIODE(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8742__CLK (.DIODE(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8743__CLK (.DIODE(\clknet_leaf_46_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8744__CLK (.DIODE(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8745__CLK (.DIODE(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8746__CLK (.DIODE(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8747__CLK (.DIODE(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8748__CLK (.DIODE(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8749__CLK (.DIODE(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8750__CLK (.DIODE(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8751__CLK (.DIODE(\clknet_leaf_34_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8752__CLK (.DIODE(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8753__CLK (.DIODE(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8754__CLK (.DIODE(\clknet_leaf_34_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8755__CLK (.DIODE(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8756__CLK (.DIODE(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8757__CLK (.DIODE(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8758__CLK (.DIODE(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8759__CLK (.DIODE(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8759__SET_B (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA__8760__CLK (.DIODE(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8760__RESET_B (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA__8761__CLK (.DIODE(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8761__RESET_B (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA__8762__CLK (.DIODE(net1743));
 sky130_fd_sc_hd__diode_2 ANTENNA__8762__RESET_B (.DIODE(rst_n));
 sky130_fd_sc_hd__diode_2 ANTENNA__8763__CLK (.DIODE(\clknet_leaf_109_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8763__RESET_B (.DIODE(rst_n));
 sky130_fd_sc_hd__diode_2 ANTENNA__8764__CLK (.DIODE(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8765__CLK (.DIODE(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8766__CLK (.DIODE(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8767__CLK (.DIODE(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8768__CLK (.DIODE(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8769__CLK (.DIODE(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8770__CLK (.DIODE(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8771__CLK (.DIODE(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8772__CLK (.DIODE(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8773__CLK (.DIODE(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8774__CLK (.DIODE(\clknet_leaf_8_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8775__CLK (.DIODE(\clknet_leaf_8_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8776__CLK (.DIODE(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8777__CLK (.DIODE(\clknet_leaf_63_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8778__CLK (.DIODE(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8779__CLK (.DIODE(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8780__CLK (.DIODE(\clknet_leaf_66_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8781__CLK (.DIODE(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8782__CLK (.DIODE(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8783__CLK (.DIODE(\clknet_leaf_67_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8784__CLK (.DIODE(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8785__CLK (.DIODE(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8786__CLK (.DIODE(\clknet_leaf_63_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8787__CLK (.DIODE(\clknet_leaf_41_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8788__CLK (.DIODE(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8789__CLK (.DIODE(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8790__CLK (.DIODE(\clknet_leaf_66_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8791__CLK (.DIODE(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8792__CLK (.DIODE(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8793__CLK (.DIODE(\clknet_leaf_66_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8794__CLK (.DIODE(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8795__CLK (.DIODE(\clknet_leaf_67_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8796__CLK (.DIODE(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8797__CLK (.DIODE(\clknet_leaf_66_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8798__CLK (.DIODE(\clknet_leaf_69_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8799__CLK (.DIODE(\clknet_leaf_66_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8800__CLK (.DIODE(\clknet_leaf_66_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8801__CLK (.DIODE(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8802__CLK (.DIODE(\clknet_leaf_66_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8803__CLK (.DIODE(\clknet_leaf_95_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8804__CLK (.DIODE(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8805__CLK (.DIODE(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8806__CLK (.DIODE(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8807__CLK (.DIODE(\clknet_leaf_95_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8808__CLK (.DIODE(\clknet_leaf_67_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8809__CLK (.DIODE(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8810__CLK (.DIODE(\clknet_leaf_8_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8811__CLK (.DIODE(\clknet_leaf_8_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8812__CLK (.DIODE(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8813__CLK (.DIODE(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8814__CLK (.DIODE(\clknet_leaf_96_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8815__CLK (.DIODE(\clknet_leaf_8_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8816__CLK (.DIODE(\clknet_leaf_8_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8817__CLK (.DIODE(\clknet_leaf_22_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8817__RESET_B (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA__8818__CLK (.DIODE(\clknet_leaf_24_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8818__RESET_B (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA__8819__CLK (.DIODE(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8819__RESET_B (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA__8820__CLK (.DIODE(\clknet_leaf_24_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8820__RESET_B (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA__8821__CLK (.DIODE(\clknet_leaf_18_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8821__RESET_B (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__8822__CLK (.DIODE(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8823__CLK (.DIODE(\clknet_leaf_23_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8823__RESET_B (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__8824__CLK (.DIODE(\clknet_leaf_17_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8824__RESET_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA__8825__CLK (.DIODE(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8825__RESET_B (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__8826__CLK (.DIODE(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8826__RESET_B (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__8827__CLK (.DIODE(\clknet_leaf_98_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8827__RESET_B (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__8828__CLK (.DIODE(\clknet_leaf_98_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8828__RESET_B (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA__8829__CLK (.DIODE(\clknet_leaf_13_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8829__RESET_B (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA__8830__CLK (.DIODE(\clknet_leaf_12_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8830__RESET_B (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__8831__CLK (.DIODE(\clknet_leaf_12_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8831__RESET_B (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA__8832__CLK (.DIODE(\clknet_leaf_12_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8832__RESET_B (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA__8833__CLK (.DIODE(\clknet_leaf_11_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8833__RESET_B (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA__8834__CLK (.DIODE(\clknet_leaf_11_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8834__RESET_B (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA__8835__CLK (.DIODE(\clknet_leaf_14_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8835__RESET_B (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__8836__CLK (.DIODE(\clknet_leaf_5_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8836__RESET_B (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA__8837__CLK (.DIODE(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8837__RESET_B (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__8838__CLK (.DIODE(\clknet_leaf_5_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8838__RESET_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__8839__CLK (.DIODE(\clknet_leaf_81_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8839__D (.DIODE(s0_wbd_lack_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8839__RESET_B (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__8840__CLK (.DIODE(\clknet_leaf_81_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8840__D (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__8841__CLK (.DIODE(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8841__RESET_B (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA__8842__CLK (.DIODE(\clknet_leaf_77_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8842__RESET_B (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__8843__CLK (.DIODE(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8843__RESET_B (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA__8844__CLK (.DIODE(\clknet_leaf_96_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8844__RESET_B (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA__8845__CLK (.DIODE(\clknet_leaf_97_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8845__RESET_B (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA__8846__CLK (.DIODE(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8846__RESET_B (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA__8847__CLK (.DIODE(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8848__CLK (.DIODE(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8849__CLK (.DIODE(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8850__CLK (.DIODE(\clknet_leaf_29_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8851__CLK (.DIODE(\clknet_leaf_11_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8852__CLK (.DIODE(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8853__CLK (.DIODE(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8854__CLK (.DIODE(\clknet_leaf_34_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8855__CLK (.DIODE(\clknet_leaf_27_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8856__CLK (.DIODE(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8857__CLK (.DIODE(\clknet_leaf_30_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8858__CLK (.DIODE(\clknet_leaf_32_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8859__CLK (.DIODE(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8860__CLK (.DIODE(\clknet_leaf_42_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8861__CLK (.DIODE(\clknet_leaf_42_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8862__CLK (.DIODE(\clknet_leaf_46_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8863__CLK (.DIODE(\clknet_leaf_49_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8864__CLK (.DIODE(\clknet_leaf_47_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8865__CLK (.DIODE(\clknet_leaf_43_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8866__CLK (.DIODE(\clknet_leaf_43_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8867__CLK (.DIODE(\clknet_leaf_45_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8868__CLK (.DIODE(\clknet_leaf_41_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8869__CLK (.DIODE(\clknet_leaf_44_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8870__CLK (.DIODE(\clknet_leaf_45_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8871__CLK (.DIODE(\clknet_leaf_40_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8872__CLK (.DIODE(\clknet_leaf_44_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8873__CLK (.DIODE(\clknet_leaf_40_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8874__CLK (.DIODE(\clknet_leaf_45_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8875__CLK (.DIODE(\clknet_leaf_43_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8876__CLK (.DIODE(\clknet_leaf_45_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8877__CLK (.DIODE(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8878__CLK (.DIODE(\clknet_leaf_45_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8879__CLK (.DIODE(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8880__CLK (.DIODE(\clknet_leaf_40_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8881__CLK (.DIODE(\clknet_leaf_63_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8882__CLK (.DIODE(\clknet_leaf_40_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8883__CLK (.DIODE(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8884__CLK (.DIODE(\clknet_leaf_40_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8885__CLK (.DIODE(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8886__CLK (.DIODE(\clknet_leaf_46_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8887__CLK (.DIODE(\clknet_leaf_32_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8888__CLK (.DIODE(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8889__CLK (.DIODE(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8890__CLK (.DIODE(\clknet_leaf_32_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8891__CLK (.DIODE(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8892__CLK (.DIODE(\clknet_leaf_32_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8893__CLK (.DIODE(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8894__CLK (.DIODE(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8895__CLK (.DIODE(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8896__CLK (.DIODE(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8897__CLK (.DIODE(\clknet_leaf_34_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8898__CLK (.DIODE(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8899__CLK (.DIODE(\clknet_leaf_32_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8900__CLK (.DIODE(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8901__CLK (.DIODE(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8902__CLK (.DIODE(\clknet_leaf_82_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8902__RESET_B (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__8903__CLK (.DIODE(\clknet_leaf_86_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8903__RESET_B (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA__8904__CLK (.DIODE(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8904__RESET_B (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__8905__CLK (.DIODE(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8905__RESET_B (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__8906__CLK (.DIODE(\clknet_leaf_77_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8906__RESET_B (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__8907__CLK (.DIODE(\clknet_leaf_77_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8907__RESET_B (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__8908__CLK (.DIODE(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8908__RESET_B (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA__8909__CLK (.DIODE(\clknet_leaf_5_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8910__CLK (.DIODE(\clknet_leaf_107_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8910__D (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8910__RESET_B (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA__8911__CLK (.DIODE(\clknet_leaf_0_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8911__RESET_B (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__8912__CLK (.DIODE(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8912__RESET_B (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__8913__CLK (.DIODE(\clknet_leaf_3_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8913__RESET_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__8914__CLK (.DIODE(\clknet_leaf_15_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8914__RESET_B (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA__8915__CLK (.DIODE(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8915__RESET_B (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__8916__CLK (.DIODE(\clknet_leaf_5_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8916__RESET_B (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA__8917__CLK (.DIODE(\clknet_leaf_5_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8917__RESET_B (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA__8918__CLK (.DIODE(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8918__RESET_B (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA__8919__CLK (.DIODE(\clknet_leaf_5_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8919__RESET_B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__8920__CLK (.DIODE(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8921__CLK (.DIODE(\clknet_leaf_19_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8921__RESET_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA__8922__CLK (.DIODE(\clknet_leaf_12_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8922__RESET_B (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA__8923__CLK (.DIODE(\clknet_leaf_20_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8923__RESET_B (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA__8924__CLK (.DIODE(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8924__RESET_B (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA__8925__CLK (.DIODE(\clknet_leaf_27_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8925__RESET_B (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA__8926__CLK (.DIODE(\clknet_leaf_27_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8926__RESET_B (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA__8927__CLK (.DIODE(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8927__RESET_B (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__8928__CLK (.DIODE(\clknet_leaf_2_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8928__RESET_B (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__8929__CLK (.DIODE(\clknet_leaf_20_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8929__RESET_B (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA__8930__CLK (.DIODE(\clknet_leaf_19_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8930__RESET_B (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA__8931__CLK (.DIODE(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8931__RESET_B (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__8932__CLK (.DIODE(\clknet_leaf_0_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8932__RESET_B (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__8933__CLK (.DIODE(\clknet_leaf_15_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8933__RESET_B (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA__8934__CLK (.DIODE(\clknet_leaf_16_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8934__RESET_B (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA__8935__CLK (.DIODE(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8935__RESET_B (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA__8936__CLK (.DIODE(\clknet_leaf_15_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8936__RESET_B (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA__8937__CLK (.DIODE(\clknet_leaf_15_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8937__RESET_B (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA__8938__CLK (.DIODE(\clknet_leaf_17_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8938__RESET_B (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__8939__CLK (.DIODE(\clknet_leaf_16_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8939__RESET_B (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA__8940__CLK (.DIODE(\clknet_leaf_17_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8940__RESET_B (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__8941__CLK (.DIODE(\clknet_leaf_5_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8941__RESET_B (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__8942__CLK (.DIODE(\clknet_leaf_5_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8942__RESET_B (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA__8943__CLK (.DIODE(\clknet_leaf_5_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8944__CLK (.DIODE(\clknet_leaf_5_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8944__RESET_B (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA__8945__CLK (.DIODE(\clknet_leaf_3_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8945__RESET_B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__8946__CLK (.DIODE(\clknet_leaf_15_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8946__RESET_B (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA__8947__CLK (.DIODE(\clknet_leaf_3_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8947__RESET_B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__8948__CLK (.DIODE(\clknet_leaf_5_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8948__RESET_B (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA__8949__CLK (.DIODE(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8949__RESET_B (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__8950__CLK (.DIODE(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8950__RESET_B (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__8951__CLK (.DIODE(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8951__RESET_B (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__8952__CLK (.DIODE(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8952__RESET_B (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__8953__CLK (.DIODE(\clknet_leaf_17_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8953__RESET_B (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__8954__CLK (.DIODE(\clknet_leaf_15_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8954__RESET_B (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA__8955__CLK (.DIODE(\clknet_leaf_15_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8955__RESET_B (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA__8956__CLK (.DIODE(\clknet_leaf_15_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8956__RESET_B (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA__8957__CLK (.DIODE(\clknet_leaf_22_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8957__RESET_B (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA__8958__CLK (.DIODE(\clknet_leaf_24_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8959__CLK (.DIODE(\clknet_leaf_16_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8959__RESET_B (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA__8960__CLK (.DIODE(\clknet_leaf_16_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8960__RESET_B (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA__8961__CLK (.DIODE(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8961__RESET_B (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA__8962__CLK (.DIODE(\clknet_leaf_18_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8962__RESET_B (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA__8963__CLK (.DIODE(\clknet_leaf_3_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8963__RESET_B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__8964__CLK (.DIODE(\clknet_leaf_16_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8965__CLK (.DIODE(\clknet_leaf_23_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8965__RESET_B (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__8966__CLK (.DIODE(\clknet_leaf_23_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8966__RESET_B (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA__8967__CLK (.DIODE(\clknet_leaf_22_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8967__RESET_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA__8968__CLK (.DIODE(\clknet_leaf_25_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8968__RESET_B (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA__8969__CLK (.DIODE(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8969__RESET_B (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA__8970__CLK (.DIODE(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8970__RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA__8971__CLK (.DIODE(\clknet_leaf_23_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8971__RESET_B (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__8972__CLK (.DIODE(\clknet_leaf_18_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8972__RESET_B (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__8973__CLK (.DIODE(\clknet_leaf_22_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8973__RESET_B (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA__8974__CLK (.DIODE(\clknet_leaf_22_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8974__RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA__8975__CLK (.DIODE(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8976__CLK (.DIODE(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8976__RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA__8977__CLK (.DIODE(\clknet_leaf_17_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8977__RESET_B (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA__8978__CLK (.DIODE(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8979__CLK (.DIODE(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8979__RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA__8980__CLK (.DIODE(\clknet_leaf_16_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8981__CLK (.DIODE(\clknet_leaf_22_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8981__RESET_B (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA__8982__CLK (.DIODE(\clknet_leaf_22_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8982__RESET_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA__8983__CLK (.DIODE(\clknet_leaf_18_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8983__RESET_B (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA__8984__CLK (.DIODE(\clknet_leaf_26_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8984__RESET_B (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA__8985__CLK (.DIODE(\clknet_leaf_17_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8985__RESET_B (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 ANTENNA__8986__CLK (.DIODE(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8986__RESET_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA__8987__CLK (.DIODE(\clknet_leaf_22_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8987__RESET_B (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA__8988__CLK (.DIODE(\clknet_leaf_16_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8989__CLK (.DIODE(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8989__D (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__8989__RESET_B (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__8990__CLK (.DIODE(net1773));
 sky130_fd_sc_hd__diode_2 ANTENNA__8991__CLK (.DIODE(net1773));
 sky130_fd_sc_hd__diode_2 ANTENNA__8992__CLK (.DIODE(net1773));
 sky130_fd_sc_hd__diode_2 ANTENNA__8993__CLK (.DIODE(net1773));
 sky130_fd_sc_hd__diode_2 ANTENNA__8993__RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__8994__CLK (.DIODE(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8995__CLK (.DIODE(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8996__CLK (.DIODE(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8997__CLK (.DIODE(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8998__CLK (.DIODE(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8999__CLK (.DIODE(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9000__CLK (.DIODE(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9001__CLK (.DIODE(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9002__CLK (.DIODE(\clknet_leaf_99_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9003__CLK (.DIODE(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9004__CLK (.DIODE(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9005__CLK (.DIODE(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9006__CLK (.DIODE(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9007__CLK (.DIODE(\clknet_leaf_63_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9008__CLK (.DIODE(\clknet_leaf_64_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9009__CLK (.DIODE(\clknet_leaf_64_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9010__CLK (.DIODE(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9011__CLK (.DIODE(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9012__CLK (.DIODE(\clknet_leaf_64_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9013__CLK (.DIODE(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9014__CLK (.DIODE(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9015__CLK (.DIODE(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9016__CLK (.DIODE(\clknet_leaf_64_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9017__CLK (.DIODE(\clknet_leaf_41_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9018__CLK (.DIODE(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9019__CLK (.DIODE(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9020__CLK (.DIODE(\clknet_leaf_67_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9021__CLK (.DIODE(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9022__CLK (.DIODE(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9023__CLK (.DIODE(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9024__CLK (.DIODE(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9025__CLK (.DIODE(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9026__CLK (.DIODE(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9027__CLK (.DIODE(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9028__CLK (.DIODE(\clknet_leaf_69_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9029__CLK (.DIODE(\clknet_leaf_66_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9030__CLK (.DIODE(\clknet_leaf_66_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9031__CLK (.DIODE(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9032__CLK (.DIODE(\clknet_leaf_67_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9033__CLK (.DIODE(\clknet_leaf_95_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9034__CLK (.DIODE(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9035__CLK (.DIODE(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9036__CLK (.DIODE(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9037__CLK (.DIODE(\clknet_leaf_95_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9038__CLK (.DIODE(\clknet_leaf_67_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9039__CLK (.DIODE(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9040__CLK (.DIODE(\clknet_leaf_8_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9041__CLK (.DIODE(\clknet_leaf_96_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9042__CLK (.DIODE(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9043__CLK (.DIODE(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9044__CLK (.DIODE(\clknet_leaf_96_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9045__CLK (.DIODE(\clknet_leaf_8_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9046__CLK (.DIODE(\clknet_leaf_8_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9047__CLK (.DIODE(net1766));
 sky130_fd_sc_hd__diode_2 ANTENNA__9047__D (.DIODE(\u_dcg_s2.cfg_mode[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9048__CLK (.DIODE(net1770));
 sky130_fd_sc_hd__diode_2 ANTENNA__9048__D (.DIODE(\u_dcg_s2.cfg_mode[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9049__CLK (.DIODE(net1766));
 sky130_fd_sc_hd__diode_2 ANTENNA__9050__CLK (.DIODE(net1770));
 sky130_fd_sc_hd__diode_2 ANTENNA__9051__CLK (.DIODE(net1770));
 sky130_fd_sc_hd__diode_2 ANTENNA__9051__RESET_B (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__9052__CLK (.DIODE(net1770));
 sky130_fd_sc_hd__diode_2 ANTENNA__9052__RESET_B (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA__9053__CLK (.DIODE(net1766));
 sky130_fd_sc_hd__diode_2 ANTENNA__9053__RESET_B (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA__9054__CLK (.DIODE(clknet_2_1__leaf_mclk_raw));
 sky130_fd_sc_hd__diode_2 ANTENNA__9054__D (.DIODE(\u_dcg_s1.cfg_mode[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9054__RESET_B (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__9055__CLK (.DIODE(net1767));
 sky130_fd_sc_hd__diode_2 ANTENNA__9055__RESET_B (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA__9056__CLK (.DIODE(clknet_2_1__leaf_mclk_raw));
 sky130_fd_sc_hd__diode_2 ANTENNA__9056__RESET_B (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__9057__CLK (.DIODE(clknet_2_1__leaf_mclk_raw));
 sky130_fd_sc_hd__diode_2 ANTENNA__9057__RESET_B (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA__9058__CLK (.DIODE(clknet_2_1__leaf_mclk_raw));
 sky130_fd_sc_hd__diode_2 ANTENNA__9058__RESET_B (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA__9059__CLK (.DIODE(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9059__SET_B (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__9060__CLK (.DIODE(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9060__RESET_B (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA__9061__CLK (.DIODE(\clknet_leaf_98_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9061__RESET_B (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__9062__CLK (.DIODE(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9063__CLK (.DIODE(\clknet_leaf_105_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9064__CLK (.DIODE(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9065__CLK (.DIODE(\clknet_leaf_97_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9066__CLK (.DIODE(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9067__CLK (.DIODE(\clknet_leaf_98_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9068__CLK (.DIODE(\clknet_leaf_97_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9069__CLK (.DIODE(\clknet_leaf_97_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9070__CLK (.DIODE(\clknet_leaf_98_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9071__CLK (.DIODE(\clknet_leaf_101_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9072__CLK (.DIODE(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9073__CLK (.DIODE(\clknet_leaf_102_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9074__CLK (.DIODE(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9075__CLK (.DIODE(\clknet_leaf_89_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9076__CLK (.DIODE(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9077__CLK (.DIODE(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9078__CLK (.DIODE(\clknet_leaf_69_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9079__CLK (.DIODE(\clknet_leaf_93_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9080__CLK (.DIODE(\clknet_leaf_86_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9081__CLK (.DIODE(\clknet_leaf_93_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9082__CLK (.DIODE(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9083__CLK (.DIODE(\clknet_leaf_86_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9084__CLK (.DIODE(\clknet_leaf_86_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9085__CLK (.DIODE(\clknet_leaf_93_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9086__CLK (.DIODE(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9087__CLK (.DIODE(\clknet_leaf_69_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9088__CLK (.DIODE(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9089__CLK (.DIODE(\clknet_leaf_87_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9090__CLK (.DIODE(\clknet_leaf_95_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9091__CLK (.DIODE(\clknet_leaf_92_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9092__CLK (.DIODE(\clknet_leaf_87_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9093__CLK (.DIODE(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9094__CLK (.DIODE(\clknet_leaf_89_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9095__CLK (.DIODE(\clknet_leaf_92_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9096__CLK (.DIODE(\clknet_leaf_87_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9097__CLK (.DIODE(\clknet_leaf_92_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9098__CLK (.DIODE(\clknet_leaf_87_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9099__CLK (.DIODE(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9100__CLK (.DIODE(\clknet_leaf_92_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9101__CLK (.DIODE(\clknet_leaf_91_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9102__CLK (.DIODE(\clknet_leaf_90_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9103__CLK (.DIODE(\clknet_leaf_101_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9104__CLK (.DIODE(\clknet_leaf_89_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9105__CLK (.DIODE(\clknet_leaf_86_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9106__CLK (.DIODE(\clknet_leaf_91_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9107__CLK (.DIODE(\clknet_leaf_90_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9108__CLK (.DIODE(\clknet_leaf_101_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9109__CLK (.DIODE(\clknet_leaf_106_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9110__CLK (.DIODE(\clknet_leaf_106_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9111__CLK (.DIODE(\clknet_leaf_101_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9112__CLK (.DIODE(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9113__CLK (.DIODE(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9114__CLK (.DIODE(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9115__CLK (.DIODE(\clknet_leaf_101_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9116__CLK (.DIODE(\clknet_leaf_105_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9117__CLK (.DIODE(\clknet_leaf_106_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9118__CLK (.DIODE(\clknet_leaf_107_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9119__CLK (.DIODE(\clknet_leaf_107_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9120__CLK (.DIODE(\clknet_leaf_107_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9121__CLK (.DIODE(\clknet_leaf_108_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9122__CLK (.DIODE(\clknet_leaf_108_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9123__CLK (.DIODE(\clknet_leaf_102_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9124__CLK (.DIODE(\clknet_leaf_102_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9125__CLK (.DIODE(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9126__CLK (.DIODE(\clknet_leaf_90_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9127__CLK (.DIODE(\clknet_leaf_106_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9128__CLK (.DIODE(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9129__CLK (.DIODE(\clknet_leaf_102_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9130__CLK (.DIODE(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9131__CLK (.DIODE(\clknet_leaf_104_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9132__CLK (.DIODE(\clknet_leaf_104_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9133__CLK (.DIODE(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9134__CLK (.DIODE(\clknet_leaf_104_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9135__CLK (.DIODE(\clknet_leaf_102_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9136__CLK (.DIODE(\clknet_leaf_105_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9137__CLK (.DIODE(\clknet_leaf_105_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9138__CLK (.DIODE(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9139__CLK (.DIODE(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9140__CLK (.DIODE(\clknet_leaf_105_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9141__CLK (.DIODE(\clknet_leaf_99_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9142__CLK (.DIODE(\clknet_leaf_97_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9143__CLK (.DIODE(\clknet_leaf_98_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9144__CLK (.DIODE(\clknet_leaf_98_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9145__CLK (.DIODE(\clknet_leaf_98_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9146__CLK (.DIODE(\clknet_leaf_97_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9147__CLK (.DIODE(\clknet_leaf_99_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9148__CLK (.DIODE(\clknet_leaf_101_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9149__CLK (.DIODE(\clknet_leaf_106_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9150__CLK (.DIODE(\clknet_leaf_102_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9151__CLK (.DIODE(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9152__CLK (.DIODE(\clknet_leaf_90_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9153__CLK (.DIODE(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9154__CLK (.DIODE(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9155__CLK (.DIODE(\clknet_leaf_69_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9156__CLK (.DIODE(\clknet_leaf_93_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9157__CLK (.DIODE(\clknet_leaf_92_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9158__CLK (.DIODE(\clknet_leaf_93_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9159__CLK (.DIODE(\clknet_leaf_93_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9160__CLK (.DIODE(\clknet_leaf_86_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9161__CLK (.DIODE(\clknet_leaf_93_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9162__CLK (.DIODE(\clknet_leaf_93_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9163__CLK (.DIODE(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9164__CLK (.DIODE(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9165__CLK (.DIODE(\clknet_leaf_89_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9166__CLK (.DIODE(\clknet_leaf_86_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9167__CLK (.DIODE(\clknet_leaf_95_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9168__CLK (.DIODE(\clknet_leaf_92_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9169__CLK (.DIODE(\clknet_leaf_92_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9170__CLK (.DIODE(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9171__CLK (.DIODE(\clknet_leaf_89_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9172__CLK (.DIODE(\clknet_leaf_91_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9173__CLK (.DIODE(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9174__CLK (.DIODE(\clknet_leaf_92_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9175__CLK (.DIODE(\clknet_leaf_89_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9176__CLK (.DIODE(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9177__CLK (.DIODE(\clknet_leaf_91_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9178__CLK (.DIODE(\clknet_leaf_91_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9179__CLK (.DIODE(\clknet_leaf_90_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9180__CLK (.DIODE(\clknet_leaf_101_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9181__CLK (.DIODE(\clknet_leaf_89_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9182__CLK (.DIODE(\clknet_leaf_92_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9183__CLK (.DIODE(\clknet_leaf_91_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9184__CLK (.DIODE(\clknet_leaf_90_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9185__CLK (.DIODE(\clknet_leaf_98_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9186__CLK (.DIODE(\clknet_leaf_106_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9187__CLK (.DIODE(\clknet_leaf_106_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9188__CLK (.DIODE(\clknet_leaf_101_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9189__CLK (.DIODE(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9190__CLK (.DIODE(\clknet_leaf_102_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9191__CLK (.DIODE(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9192__CLK (.DIODE(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9193__CLK (.DIODE(\clknet_leaf_105_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9194__CLK (.DIODE(\clknet_leaf_106_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9195__CLK (.DIODE(\clknet_leaf_107_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9196__CLK (.DIODE(\clknet_leaf_107_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9197__CLK (.DIODE(\clknet_leaf_108_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9198__CLK (.DIODE(\clknet_leaf_108_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9199__CLK (.DIODE(\clknet_leaf_108_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9200__CLK (.DIODE(\clknet_leaf_102_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9201__CLK (.DIODE(\clknet_leaf_102_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9202__CLK (.DIODE(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9203__CLK (.DIODE(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9204__CLK (.DIODE(\clknet_leaf_106_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9205__CLK (.DIODE(\clknet_leaf_104_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9206__CLK (.DIODE(\clknet_leaf_106_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9207__CLK (.DIODE(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9208__CLK (.DIODE(\clknet_leaf_104_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9209__CLK (.DIODE(\clknet_leaf_104_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9210__CLK (.DIODE(\clknet_leaf_104_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9211__CLK (.DIODE(\clknet_leaf_104_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9212__CLK (.DIODE(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9213__CLK (.DIODE(\clknet_leaf_105_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9214__CLK (.DIODE(\clknet_leaf_108_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9215__CLK (.DIODE(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9216__CLK (.DIODE(net1770));
 sky130_fd_sc_hd__diode_2 ANTENNA__9216__D (.DIODE(\u_dcg_s0.cfg_mode[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9216__RESET_B (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__9217__CLK (.DIODE(clknet_2_2__leaf_mclk_raw));
 sky130_fd_sc_hd__diode_2 ANTENNA__9217__D (.DIODE(net1279));
 sky130_fd_sc_hd__diode_2 ANTENNA__9217__RESET_B (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA__9218__CLK (.DIODE(clknet_2_2__leaf_mclk_raw));
 sky130_fd_sc_hd__diode_2 ANTENNA__9218__D (.DIODE(\u_dcg_s0.u_dsync.in_data_s[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9218__RESET_B (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA__9219__CLK (.DIODE(clknet_2_2__leaf_mclk_raw));
 sky130_fd_sc_hd__diode_2 ANTENNA__9219__RESET_B (.DIODE(net890));
 sky130_fd_sc_hd__diode_2 ANTENNA__9220__CLK (.DIODE(net1773));
 sky130_fd_sc_hd__diode_2 ANTENNA__9220__D (.DIODE(net1922));
 sky130_fd_sc_hd__diode_2 ANTENNA__9220__RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__9221__CLK (.DIODE(net1773));
 sky130_fd_sc_hd__diode_2 ANTENNA__9221__RESET_B (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA__9222__CLK (.DIODE(clknet_2_3__leaf_mclk_raw));
 sky130_fd_sc_hd__diode_2 ANTENNA__9222__D (.DIODE(net1511));
 sky130_fd_sc_hd__diode_2 ANTENNA__9222__RESET_B (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA__9223__CLK (.DIODE(clknet_2_3__leaf_mclk_raw));
 sky130_fd_sc_hd__diode_2 ANTENNA__9223__SET_B (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA__9224__CLK (.DIODE(\clknet_leaf_0_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9224__RESET_B (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA__9225__CLK (.DIODE(\clknet_leaf_107_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9225__RESET_B (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA__9226__CLK (.DIODE(net1770));
 sky130_fd_sc_hd__diode_2 ANTENNA__9226__D (.DIODE(\u_dcg_riscv.cfg_mode[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9227__CLK (.DIODE(net1771));
 sky130_fd_sc_hd__diode_2 ANTENNA__9227__RESET_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__9228__CLK (.DIODE(net1770));
 sky130_fd_sc_hd__diode_2 ANTENNA__9229__CLK (.DIODE(net1771));
 sky130_fd_sc_hd__diode_2 ANTENNA__9229__RESET_B (.DIODE(net907));
 sky130_fd_sc_hd__diode_2 ANTENNA__9230__CLK (.DIODE(net1770));
 sky130_fd_sc_hd__diode_2 ANTENNA__9231__CLK (.DIODE(net1771));
 sky130_fd_sc_hd__diode_2 ANTENNA__9231__RESET_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__9232__CLK (.DIODE(net1766));
 sky130_fd_sc_hd__diode_2 ANTENNA__9233__CLK (.DIODE(net1766));
 sky130_fd_sc_hd__diode_2 ANTENNA__9233__D (.DIODE(\u_dcg_peri.cfg_mode[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__9233__RESET_B (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA__9234__CLK (.DIODE(net1766));
 sky130_fd_sc_hd__diode_2 ANTENNA__9235__CLK (.DIODE(net1766));
 sky130_fd_sc_hd__diode_2 ANTENNA__9236__CLK (.DIODE(net1766));
 sky130_fd_sc_hd__diode_2 ANTENNA__9237__CLK (.DIODE(net1766));
 sky130_fd_sc_hd__diode_2 ANTENNA__9237__RESET_B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__9254__A (.DIODE(ch_clk_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9255__A (.DIODE(net1716));
 sky130_fd_sc_hd__diode_2 ANTENNA__9256__A (.DIODE(net1715));
 sky130_fd_sc_hd__diode_2 ANTENNA__9257__A (.DIODE(ch_data_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9258__A (.DIODE(ch_data_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9259__A (.DIODE(ch_data_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9260__A (.DIODE(ch_data_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9261__A (.DIODE(ch_data_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9262__A (.DIODE(ch_data_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9263__A (.DIODE(ch_data_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9264__A (.DIODE(ch_data_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9265__A (.DIODE(ch_data_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9266__A (.DIODE(ch_data_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9267__A (.DIODE(ch_data_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9268__A (.DIODE(ch_data_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9269__A (.DIODE(net1689));
 sky130_fd_sc_hd__diode_2 ANTENNA__9270__A (.DIODE(net1686));
 sky130_fd_sc_hd__diode_2 ANTENNA__9271__A (.DIODE(net1680));
 sky130_fd_sc_hd__diode_2 ANTENNA__9272__A (.DIODE(net1663));
 sky130_fd_sc_hd__diode_2 ANTENNA__9273__A (.DIODE(ch_data_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9274__A (.DIODE(ch_data_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9275__A (.DIODE(ch_data_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9276__A (.DIODE(ch_data_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9277__A (.DIODE(ch_data_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9278__A (.DIODE(ch_data_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9279__A (.DIODE(ch_data_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9280__A (.DIODE(ch_data_in[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9281__A (.DIODE(net1662));
 sky130_fd_sc_hd__diode_2 ANTENNA__9282__A (.DIODE(net1661));
 sky130_fd_sc_hd__diode_2 ANTENNA__9283__A (.DIODE(net1660));
 sky130_fd_sc_hd__diode_2 ANTENNA__9284__A (.DIODE(net1659));
 sky130_fd_sc_hd__diode_2 ANTENNA__9285__A (.DIODE(net1658));
 sky130_fd_sc_hd__diode_2 ANTENNA__9286__A (.DIODE(net1657));
 sky130_fd_sc_hd__diode_2 ANTENNA__9287__A (.DIODE(net1656));
 sky130_fd_sc_hd__diode_2 ANTENNA__9288__A (.DIODE(net1655));
 sky130_fd_sc_hd__diode_2 ANTENNA__9289__A (.DIODE(net1654));
 sky130_fd_sc_hd__diode_2 ANTENNA__9290__A (.DIODE(net1653));
 sky130_fd_sc_hd__diode_2 ANTENNA__9291__A (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__9292__A (.DIODE(net1651));
 sky130_fd_sc_hd__diode_2 ANTENNA__9293__A (.DIODE(net1650));
 sky130_fd_sc_hd__diode_2 ANTENNA__9294__A (.DIODE(net1649));
 sky130_fd_sc_hd__diode_2 ANTENNA__9295__A (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA__9296__A (.DIODE(net1647));
 sky130_fd_sc_hd__diode_2 ANTENNA__9297__A (.DIODE(net1646));
 sky130_fd_sc_hd__diode_2 ANTENNA__9298__A (.DIODE(net1645));
 sky130_fd_sc_hd__diode_2 ANTENNA__9299__A (.DIODE(net1644));
 sky130_fd_sc_hd__diode_2 ANTENNA__9300__A (.DIODE(net1643));
 sky130_fd_sc_hd__diode_2 ANTENNA__9301__A (.DIODE(ch_data_in[44]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9302__A (.DIODE(ch_data_in[45]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9303__A (.DIODE(ch_data_in[46]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9304__A (.DIODE(ch_data_in[47]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9305__A (.DIODE(ch_data_in[48]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9306__A (.DIODE(ch_data_in[49]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9307__A (.DIODE(ch_data_in[50]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9308__A (.DIODE(ch_data_in[51]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9309__A (.DIODE(ch_data_in[52]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9310__A (.DIODE(ch_data_in[53]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9311__A (.DIODE(ch_data_in[54]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9312__A (.DIODE(ch_data_in[55]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9313__A (.DIODE(ch_data_in[56]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9314__A (.DIODE(ch_data_in[57]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9315__A (.DIODE(ch_data_in[58]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9316__A (.DIODE(ch_data_in[59]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9317__A (.DIODE(ch_data_in[60]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9318__A (.DIODE(ch_data_in[61]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9319__A (.DIODE(ch_data_in[62]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9320__A (.DIODE(ch_data_in[63]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9321__A (.DIODE(ch_data_in[64]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9322__A (.DIODE(ch_data_in[65]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9323__A (.DIODE(ch_data_in[66]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9324__A (.DIODE(ch_data_in[67]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9325__A (.DIODE(ch_data_in[68]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9326__A (.DIODE(ch_data_in[69]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9327__A (.DIODE(ch_data_in[70]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9328__A (.DIODE(ch_data_in[71]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9329__A (.DIODE(ch_data_in[72]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9330__A (.DIODE(ch_data_in[73]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9331__A (.DIODE(ch_data_in[74]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9332__A (.DIODE(ch_data_in[75]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9333__A (.DIODE(ch_data_in[76]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9334__A (.DIODE(net1641));
 sky130_fd_sc_hd__diode_2 ANTENNA__9335__A (.DIODE(net1639));
 sky130_fd_sc_hd__diode_2 ANTENNA__9336__A (.DIODE(net1637));
 sky130_fd_sc_hd__diode_2 ANTENNA__9337__A (.DIODE(net1635));
 sky130_fd_sc_hd__diode_2 ANTENNA__9338__A (.DIODE(net1633));
 sky130_fd_sc_hd__diode_2 ANTENNA__9339__A (.DIODE(net1631));
 sky130_fd_sc_hd__diode_2 ANTENNA__9340__A (.DIODE(net1629));
 sky130_fd_sc_hd__diode_2 ANTENNA__9341__A (.DIODE(net1627));
 sky130_fd_sc_hd__diode_2 ANTENNA__9342__A (.DIODE(net1625));
 sky130_fd_sc_hd__diode_2 ANTENNA__9343__A (.DIODE(net1623));
 sky130_fd_sc_hd__diode_2 ANTENNA__9344__A (.DIODE(net1621));
 sky130_fd_sc_hd__diode_2 ANTENNA__9345__A (.DIODE(net1619));
 sky130_fd_sc_hd__diode_2 ANTENNA__9346__A (.DIODE(net1617));
 sky130_fd_sc_hd__diode_2 ANTENNA__9347__A (.DIODE(net1615));
 sky130_fd_sc_hd__diode_2 ANTENNA__9348__A (.DIODE(net1613));
 sky130_fd_sc_hd__diode_2 ANTENNA__9349__A (.DIODE(net1611));
 sky130_fd_sc_hd__diode_2 ANTENNA__9350__A (.DIODE(net1609));
 sky130_fd_sc_hd__diode_2 ANTENNA__9351__A (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__9352__A (.DIODE(net1605));
 sky130_fd_sc_hd__diode_2 ANTENNA__9353__A (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__9354__A (.DIODE(net1601));
 sky130_fd_sc_hd__diode_2 ANTENNA__9355__A (.DIODE(net1600));
 sky130_fd_sc_hd__diode_2 ANTENNA__9356__A (.DIODE(net1599));
 sky130_fd_sc_hd__diode_2 ANTENNA__9357__A (.DIODE(net1713));
 sky130_fd_sc_hd__diode_2 ANTENNA__9358__A (.DIODE(net1711));
 sky130_fd_sc_hd__diode_2 ANTENNA__9359__A (.DIODE(net1709));
 sky130_fd_sc_hd__diode_2 ANTENNA__9360__A (.DIODE(net1707));
 sky130_fd_sc_hd__diode_2 ANTENNA__9361__A (.DIODE(net1705));
 sky130_fd_sc_hd__diode_2 ANTENNA__9362__A (.DIODE(net1703));
 sky130_fd_sc_hd__diode_2 ANTENNA__9363__A (.DIODE(net1701));
 sky130_fd_sc_hd__diode_2 ANTENNA__9364__A (.DIODE(net1699));
 sky130_fd_sc_hd__diode_2 ANTENNA__9365__A (.DIODE(net1697));
 sky130_fd_sc_hd__diode_2 ANTENNA__9366__A (.DIODE(net1695));
 sky130_fd_sc_hd__diode_2 ANTENNA__9367__A (.DIODE(net1693));
 sky130_fd_sc_hd__diode_2 ANTENNA__9368__A (.DIODE(net1691));
 sky130_fd_sc_hd__diode_2 ANTENNA__9369__A (.DIODE(ch_data_in[112]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9370__A (.DIODE(ch_data_in[113]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9371__A (.DIODE(ch_data_in[114]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9372__A (.DIODE(ch_data_in[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9373__A (.DIODE(ch_data_in[116]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9374__A (.DIODE(ch_data_in[117]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9375__A (.DIODE(ch_data_in[118]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9376__A (.DIODE(ch_data_in[119]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9377__A (.DIODE(ch_data_in[120]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9378__A (.DIODE(ch_data_in[121]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9379__A (.DIODE(ch_data_in[122]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9380__A (.DIODE(ch_data_in[123]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9381__A (.DIODE(ch_data_in[124]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9382__A (.DIODE(ch_data_in[125]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9383__A (.DIODE(ch_data_in[126]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9384__A (.DIODE(ch_data_in[127]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9385__A (.DIODE(ch_data_in[128]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9386__A (.DIODE(ch_data_in[129]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9387__A (.DIODE(ch_data_in[130]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9388__A (.DIODE(ch_data_in[131]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9389__A (.DIODE(ch_data_in[132]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9390__A (.DIODE(ch_data_in[133]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9391__A (.DIODE(ch_data_in[134]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9392__A (.DIODE(ch_data_in[135]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9393__A (.DIODE(ch_data_in[136]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9394__A (.DIODE(ch_data_in[137]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9395__A (.DIODE(ch_data_in[138]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9396__A (.DIODE(net1688));
 sky130_fd_sc_hd__diode_2 ANTENNA__9397__A (.DIODE(net1685));
 sky130_fd_sc_hd__diode_2 ANTENNA__9398__A (.DIODE(net1684));
 sky130_fd_sc_hd__diode_2 ANTENNA__9399__A (.DIODE(net1683));
 sky130_fd_sc_hd__diode_2 ANTENNA__9400__A (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA__9401__A (.DIODE(ch_data_in[144]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9402__A (.DIODE(ch_data_in[145]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9403__A (.DIODE(ch_data_in[146]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9404__A (.DIODE(ch_data_in[147]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9405__A (.DIODE(ch_data_in[148]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9406__A (.DIODE(ch_data_in[149]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9407__A (.DIODE(net1677));
 sky130_fd_sc_hd__diode_2 ANTENNA__9408__A (.DIODE(net1674));
 sky130_fd_sc_hd__diode_2 ANTENNA__9409__A (.DIODE(ch_data_in[152]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9410__A (.DIODE(ch_data_in[153]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9411__A (.DIODE(ch_data_in[154]));
 sky130_fd_sc_hd__diode_2 ANTENNA__9412__A (.DIODE(net1671));
 sky130_fd_sc_hd__diode_2 ANTENNA__9413__A (.DIODE(net1668));
 sky130_fd_sc_hd__diode_2 ANTENNA__9414__A (.DIODE(net1665));
 sky130_fd_sc_hd__diode_2 ANTENNA__9415__A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__9416__A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__9417__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_mclk_raw_A (.DIODE(net1761));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_0_u_dsync.out_clk_A  (.DIODE(net1733));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0_0_mclk_raw_A (.DIODE(net1764));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_1_0_0_u_dsync.out_clk_A  (.DIODE(net1737));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1_0_mclk_raw_A (.DIODE(net1765));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_1_1_0_u_dsync.out_clk_A  (.DIODE(net1736));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_mclk_raw_A (.DIODE(clknet_1_0_0_mclk_raw));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_mclk_raw_A (.DIODE(clknet_1_0_0_mclk_raw));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_mclk_raw_A (.DIODE(clknet_1_1_0_mclk_raw));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_mclk_raw_A (.DIODE(clknet_1_1_0_mclk_raw));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_3_0__f_u_dsync.out_clk_A  (.DIODE(net1738));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_3_1__f_u_dsync.out_clk_A  (.DIODE(net1739));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_3_2__f_u_dsync.out_clk_A  (.DIODE(net1738));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_3_3__f_u_dsync.out_clk_A  (.DIODE(net1739));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_3_4__f_u_dsync.out_clk_A  (.DIODE(\clknet_1_1_0_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_3_5__f_u_dsync.out_clk_A  (.DIODE(net1740));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_3_6__f_u_dsync.out_clk_A  (.DIODE(net1741));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_3_7__f_u_dsync.out_clk_A  (.DIODE(net1740));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_0_u_dsync.out_clk_A  (.DIODE(net1742));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_100_u_dsync.out_clk_A  (.DIODE(net1742));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_101_u_dsync.out_clk_A  (.DIODE(net1742));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_102_u_dsync.out_clk_A  (.DIODE(\clknet_3_0__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_103_u_dsync.out_clk_A  (.DIODE(net1743));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_104_u_dsync.out_clk_A  (.DIODE(net1744));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_105_u_dsync.out_clk_A  (.DIODE(net1744));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_106_u_dsync.out_clk_A  (.DIODE(\clknet_3_0__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_107_u_dsync.out_clk_A  (.DIODE(\clknet_3_0__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_108_u_dsync.out_clk_A  (.DIODE(net1743));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_109_u_dsync.out_clk_A  (.DIODE(net1744));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_10_u_dsync.out_clk_A  (.DIODE(net1753));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_11_u_dsync.out_clk_A  (.DIODE(net1754));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_12_u_dsync.out_clk_A  (.DIODE(\clknet_3_4__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_13_u_dsync.out_clk_A  (.DIODE(net1754));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_14_u_dsync.out_clk_A  (.DIODE(net1753));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_15_u_dsync.out_clk_A  (.DIODE(net1753));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_16_u_dsync.out_clk_A  (.DIODE(net1753));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_17_u_dsync.out_clk_A  (.DIODE(net1754));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_18_u_dsync.out_clk_A  (.DIODE(net1752));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_19_u_dsync.out_clk_A  (.DIODE(net1752));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_1_u_dsync.out_clk_A  (.DIODE(net1746));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_20_u_dsync.out_clk_A  (.DIODE(net1752));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_21_u_dsync.out_clk_A  (.DIODE(net1755));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_22_u_dsync.out_clk_A  (.DIODE(\clknet_3_5__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_23_u_dsync.out_clk_A  (.DIODE(net1757));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_24_u_dsync.out_clk_A  (.DIODE(net1757));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_25_u_dsync.out_clk_A  (.DIODE(net1757));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_26_u_dsync.out_clk_A  (.DIODE(net1755));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_27_u_dsync.out_clk_A  (.DIODE(net1755));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_28_u_dsync.out_clk_A  (.DIODE(net1757));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_29_u_dsync.out_clk_A  (.DIODE(net1756));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_2_u_dsync.out_clk_A  (.DIODE(\clknet_3_1__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_30_u_dsync.out_clk_A  (.DIODE(net1756));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_31_u_dsync.out_clk_A  (.DIODE(net1756));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_32_u_dsync.out_clk_A  (.DIODE(net1758));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_33_u_dsync.out_clk_A  (.DIODE(net1755));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_34_u_dsync.out_clk_A  (.DIODE(net1755));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_35_u_dsync.out_clk_A  (.DIODE(\clknet_3_4__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_36_u_dsync.out_clk_A  (.DIODE(net1759));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_37_u_dsync.out_clk_A  (.DIODE(\clknet_3_6__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_38_u_dsync.out_clk_A  (.DIODE(\clknet_3_6__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_39_u_dsync.out_clk_A  (.DIODE(\clknet_3_6__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_3_u_dsync.out_clk_A  (.DIODE(net1745));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_40_u_dsync.out_clk_A  (.DIODE(net1759));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_41_u_dsync.out_clk_A  (.DIODE(\clknet_3_6__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_42_u_dsync.out_clk_A  (.DIODE(net1759));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_43_u_dsync.out_clk_A  (.DIODE(net1758));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_44_u_dsync.out_clk_A  (.DIODE(net1758));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_45_u_dsync.out_clk_A  (.DIODE(net1757));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_46_u_dsync.out_clk_A  (.DIODE(net1756));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_47_u_dsync.out_clk_A  (.DIODE(net1756));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_48_u_dsync.out_clk_A  (.DIODE(net1760));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_49_u_dsync.out_clk_A  (.DIODE(\clknet_3_7__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_4_u_dsync.out_clk_A  (.DIODE(net1745));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_50_u_dsync.out_clk_A  (.DIODE(\clknet_3_7__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_51_u_dsync.out_clk_A  (.DIODE(net1760));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_52_u_dsync.out_clk_A  (.DIODE(net1760));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_53_u_dsync.out_clk_A  (.DIODE(\clknet_3_7__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_54_u_dsync.out_clk_A  (.DIODE(\clknet_3_7__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_55_u_dsync.out_clk_A  (.DIODE(net1759));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_56_u_dsync.out_clk_A  (.DIODE(\clknet_3_6__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_57_u_dsync.out_clk_A  (.DIODE(\clknet_3_6__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_58_u_dsync.out_clk_A  (.DIODE(\clknet_3_6__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_59_u_dsync.out_clk_A  (.DIODE(\clknet_3_6__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_5_u_dsync.out_clk_A  (.DIODE(\clknet_3_1__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_60_u_dsync.out_clk_A  (.DIODE(\clknet_3_6__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_61_u_dsync.out_clk_A  (.DIODE(\clknet_3_6__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_62_u_dsync.out_clk_A  (.DIODE(\clknet_3_6__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_63_u_dsync.out_clk_A  (.DIODE(\clknet_3_6__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_64_u_dsync.out_clk_A  (.DIODE(\clknet_3_6__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_65_u_dsync.out_clk_A  (.DIODE(\clknet_3_6__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_66_u_dsync.out_clk_A  (.DIODE(net1750));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_67_u_dsync.out_clk_A  (.DIODE(net1750));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_68_u_dsync.out_clk_A  (.DIODE(net1750));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_69_u_dsync.out_clk_A  (.DIODE(\clknet_3_3__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_6_u_dsync.out_clk_A  (.DIODE(\clknet_3_1__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_70_u_dsync.out_clk_A  (.DIODE(net1749));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_71_u_dsync.out_clk_A  (.DIODE(net1751));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_72_u_dsync.out_clk_A  (.DIODE(net1751));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_73_u_dsync.out_clk_A  (.DIODE(net1751));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_74_u_dsync.out_clk_A  (.DIODE(net1751));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_75_u_dsync.out_clk_A  (.DIODE(\clknet_3_3__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_76_u_dsync.out_clk_A  (.DIODE(net1749));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_77_u_dsync.out_clk_A  (.DIODE(net1749));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_78_u_dsync.out_clk_A  (.DIODE(net1748));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_79_u_dsync.out_clk_A  (.DIODE(net1748));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_7_u_dsync.out_clk_A  (.DIODE(net1745));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_80_u_dsync.out_clk_A  (.DIODE(\clknet_3_2__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_81_u_dsync.out_clk_A  (.DIODE(net1747));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_82_u_dsync.out_clk_A  (.DIODE(net1747));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_83_u_dsync.out_clk_A  (.DIODE(net1747));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_84_u_dsync.out_clk_A  (.DIODE(net1747));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_85_u_dsync.out_clk_A  (.DIODE(\clknet_3_2__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_86_u_dsync.out_clk_A  (.DIODE(net1748));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_87_u_dsync.out_clk_A  (.DIODE(\clknet_3_2__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_88_u_dsync.out_clk_A  (.DIODE(net1747));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_89_u_dsync.out_clk_A  (.DIODE(net1744));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_8_u_dsync.out_clk_A  (.DIODE(net1745));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_90_u_dsync.out_clk_A  (.DIODE(net1744));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_91_u_dsync.out_clk_A  (.DIODE(net1742));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_92_u_dsync.out_clk_A  (.DIODE(net1742));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_93_u_dsync.out_clk_A  (.DIODE(net1749));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_94_u_dsync.out_clk_A  (.DIODE(net1749));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_95_u_dsync.out_clk_A  (.DIODE(\clknet_3_3__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_96_u_dsync.out_clk_A  (.DIODE(net1745));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_97_u_dsync.out_clk_A  (.DIODE(\clknet_3_1__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_98_u_dsync.out_clk_A  (.DIODE(net1746));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_99_u_dsync.out_clk_A  (.DIODE(net1746));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_9_u_dsync.out_clk_A  (.DIODE(net1753));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1000_A (.DIODE(_2800_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1001_A (.DIODE(_2800_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1002_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1003_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1143_A (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1144_A (.DIODE(_2021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1145_A (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1146_A (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1147_A (.DIODE(_2021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1148_A (.DIODE(net1152));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1149_A (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1150_A (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1151_A (.DIODE(net1152));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1153_A (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1154_A (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1155_A (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1156_A (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1158_A (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1159_A (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1162_A (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1163_A (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1164_A (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1165_A (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1166_A (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1167_A (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1168_A (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1169_A (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1170_A (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1172_A (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1174_A (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1175_A (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1177_A (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1178_A (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1182_A (.DIODE(_1851_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1183_A (.DIODE(_1833_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1184_A (.DIODE(_1833_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1185_A (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1186_A (.DIODE(_1832_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1187_A (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1188_A (.DIODE(_1831_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1189_A (.DIODE(net1190));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1190_A (.DIODE(net1191));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1191_A (.DIODE(_1831_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1192_A (.DIODE(_1830_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1193_A (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1194_A (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1195_A (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1196_A (.DIODE(net1198));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1197_A (.DIODE(net1198));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1198_A (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1199_A (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1200_A (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1201_A (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1202_A (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1203_A (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1204_A (.DIODE(net1205));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1205_A (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1206_A (.DIODE(net1209));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1207_A (.DIODE(net1208));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1208_A (.DIODE(net1209));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1210_A (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1211_A (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1212_A (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1214_A (.DIODE(net1217));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1215_A (.DIODE(net1217));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1216_A (.DIODE(net1217));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1217_A (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1219_A (.DIODE(net1223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1220_A (.DIODE(net1223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1221_A (.DIODE(net1223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1222_A (.DIODE(net1223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1224_A (.DIODE(_1677_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1225_A (.DIODE(_1677_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1226_A (.DIODE(net1231));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1227_A (.DIODE(net1231));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1228_A (.DIODE(net1231));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1229_A (.DIODE(net1230));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1230_A (.DIODE(net1231));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1231_A (.DIODE(_1677_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1232_A (.DIODE(net1233));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1233_A (.DIODE(net1238));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1234_A (.DIODE(net1235));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1236_A (.DIODE(net1237));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1237_A (.DIODE(net1238));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1239_A (.DIODE(net1240));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1240_A (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1242_A (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1243_A (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1244_A (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1245_A (.DIODE(net1246));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1246_A (.DIODE(net1252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1247_A (.DIODE(net1252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1248_A (.DIODE(net1252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1249_A (.DIODE(net1250));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1250_A (.DIODE(net1251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1251_A (.DIODE(net1252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1253_A (.DIODE(net1254));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1254_A (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1257_A (.DIODE(net1258));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1258_A (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1259_A (.DIODE(net1263));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1260_A (.DIODE(net1263));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1261_A (.DIODE(net1263));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1262_A (.DIODE(net1263));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1263_A (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1264_A (.DIODE(net1268));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1266_A (.DIODE(net1267));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1267_A (.DIODE(net1268));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1268_A (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1269_A (.DIODE(net1271));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1270_A (.DIODE(net1271));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1271_A (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1272_A (.DIODE(net1273));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1273_A (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1274_A (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1275_A (.DIODE(\u_wbi_arb.gnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1276_A (.DIODE(net1277));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1277_A (.DIODE(net1278));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1313_A (.DIODE(net1317));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1314_A (.DIODE(net1317));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1315_A (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1316_A (.DIODE(net1317));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1318_A (.DIODE(net1322));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1319_A (.DIODE(net1322));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1320_A (.DIODE(net1321));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1321_A (.DIODE(net1322));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1323_A (.DIODE(net1325));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1324_A (.DIODE(net1325));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1325_A (.DIODE(net1332));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1326_A (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1327_A (.DIODE(net1332));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1328_A (.DIODE(net1332));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1329_A (.DIODE(net1332));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1330_A (.DIODE(net1332));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1331_A (.DIODE(net1332));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1333_A (.DIODE(net1335));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1334_A (.DIODE(net1335));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1335_A (.DIODE(net1342));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1336_A (.DIODE(net1337));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1337_A (.DIODE(net1342));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1338_A (.DIODE(net1342));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1339_A (.DIODE(net1342));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1340_A (.DIODE(net1342));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1341_A (.DIODE(net1342));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1343_A (.DIODE(net1344));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1344_A (.DIODE(\u_s1.u_sync_wbb.u_resp_if.rd_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1345_A (.DIODE(\u_s1.u_sync_wbb.u_resp_if.rd_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1346_A (.DIODE(\u_s1.u_sync_wbb.u_resp_if.rd_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1347_A (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1348_A (.DIODE(net1351));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1349_A (.DIODE(net1351));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1350_A (.DIODE(net1351));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1352_A (.DIODE(net1354));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1353_A (.DIODE(net1354));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1354_A (.DIODE(\u_s1.u_sync_wbb.u_cmd_if.rd_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1355_A (.DIODE(net1358));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1356_A (.DIODE(net1358));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1357_A (.DIODE(net1358));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1358_A (.DIODE(\u_s1.u_sync_wbb.u_cmd_if.rd_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1359_A (.DIODE(net1361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1360_A (.DIODE(net1361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1361_A (.DIODE(\u_s1.u_sync_wbb.u_cmd_if.rd_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1362_A (.DIODE(net1365));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1363_A (.DIODE(net1365));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1364_A (.DIODE(net1365));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1365_A (.DIODE(\u_s1.u_sync_wbb.u_cmd_if.rd_ptr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1368_A (.DIODE(net1370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1369_A (.DIODE(net1370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1370_A (.DIODE(net1371));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1372_A (.DIODE(net1374));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1373_A (.DIODE(net1374));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1374_A (.DIODE(\u_s0.gnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1375_A (.DIODE(\u_s0.gnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1376_A (.DIODE(\u_s2.u_sync_wbb.u_resp_if.rd_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1377_A (.DIODE(\u_s2.u_sync_wbb.u_resp_if.rd_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1378_A (.DIODE(net1379));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1379_A (.DIODE(\u_s2.u_sync_wbb.u_resp_if.rd_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1380_A (.DIODE(net1384));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1381_A (.DIODE(net1384));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1382_A (.DIODE(net1383));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1383_A (.DIODE(net1384));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1385_A (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.rd_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1386_A (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.rd_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1387_A (.DIODE(net1388));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1388_A (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.rd_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1389_A (.DIODE(net1391));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1390_A (.DIODE(net1391));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1391_A (.DIODE(\u_s2.u_sync_wbb.u_cmd_if.rd_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1392_A (.DIODE(net1399));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1393_A (.DIODE(net1399));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1394_A (.DIODE(net1395));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1395_A (.DIODE(net1399));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1396_A (.DIODE(net1399));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1397_A (.DIODE(net1399));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1398_A (.DIODE(net1399));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1404_A (.DIODE(\u_s1.gnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1405_A (.DIODE(\u_s1.gnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1406_A (.DIODE(\u_s1.gnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1407_A (.DIODE(net1408));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1408_A (.DIODE(\u_s2.gnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1409_A (.DIODE(net1410));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1410_A (.DIODE(\u_s2.gnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1495_A (.DIODE(net1498));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1496_A (.DIODE(net1498));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1497_A (.DIODE(net1498));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1498_A (.DIODE(net1784));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1499_A (.DIODE(net1784));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1500_A (.DIODE(net1784));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1501_A (.DIODE(net1502));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1502_A (.DIODE(net1784));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1503_A (.DIODE(net1504));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1504_A (.DIODE(net1510));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1505_A (.DIODE(net1510));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1506_A (.DIODE(net1510));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1507_A (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1508_A (.DIODE(net1509));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1509_A (.DIODE(net1510));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout481_A (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout482_A (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout483_A (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout484_A (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout488_A (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout490_A (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout491_A (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout492_A (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout494_A (.DIODE(_3131_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout495_A (.DIODE(_3131_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout496_A (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout497_A (.DIODE(_3131_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout498_A (.DIODE(_2788_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout499_A (.DIODE(_2788_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout500_A (.DIODE(_2788_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout501_A (.DIODE(_2788_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout502_A (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout503_A (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout504_A (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout505_A (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout506_A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout507_A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout508_A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout513_A (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout514_A (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout518_A (.DIODE(_3432_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout521_A (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout522_A (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout523_A (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout525_A (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout526_A (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout527_A (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout529_A (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout530_A (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout531_A (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout533_A (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout534_A (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout535_A (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout537_A (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout538_A (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout539_A (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout541_A (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout542_A (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout543_A (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout544_A (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout546_A (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout547_A (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout548_A (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout562_A (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout563_A (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout564_A (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout565_A (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout566_A (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout567_A (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout568_A (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout569_A (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout570_A (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout574_A (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout580_A (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout581_A (.DIODE(_1998_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout583_A (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout586_A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout587_A (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout589_A (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout594_A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout595_A (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout596_A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout599_A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout600_A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout601_A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout603_A (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout605_A (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout606_A (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout612_A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout618_A (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout619_A (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout622_A (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout623_A (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout624_A (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout626_A (.DIODE(_2024_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout627_A (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout713_A (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout714_A (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout715_A (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout716_A (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout717_A (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout721_A (.DIODE(_1960_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout722_A (.DIODE(_1960_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout723_A (.DIODE(_1960_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout724_A (.DIODE(_1960_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout733_A (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout734_A (.DIODE(_1769_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout735_A (.DIODE(_1769_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout736_A (.DIODE(_1769_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout739_A (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout740_A (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout741_A (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout742_A (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout743_A (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout744_A (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout745_A (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout746_A (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout747_A (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout749_A (.DIODE(net750));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout750_A (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout751_A (.DIODE(_2944_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout752_A (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout753_A (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout754_A (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout755_A (.DIODE(_2944_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout756_A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout757_A (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout758_A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout760_A (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout761_A (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout762_A (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout766_A (.DIODE(net1776));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout767_A (.DIODE(net1776));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout768_A (.DIODE(_2189_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout769_A (.DIODE(_2189_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout770_A (.DIODE(_2189_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout771_A (.DIODE(_2189_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout772_A (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout773_A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout774_A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout775_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout776_A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout777_A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout779_A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout781_A (.DIODE(net1775));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout782_A (.DIODE(net1775));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout799_A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout801_A (.DIODE(net1774));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout802_A (.DIODE(net1774));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout803_A (.DIODE(_1852_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout804_A (.DIODE(_1852_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout805_A (.DIODE(_1852_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout806_A (.DIODE(_1852_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout809_A (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout810_A (.DIODE(_1780_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout811_A (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout812_A (.DIODE(_1780_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout813_A (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout814_A (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout815_A (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout816_A (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout817_A (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout818_A (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout819_A (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout820_A (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout821_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout822_A (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout823_A (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout824_A (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout826_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout827_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout828_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout829_A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout830_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout831_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout832_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout834_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout835_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout836_A (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout837_A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout838_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout839_A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout840_A (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout841_A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout842_A (.DIODE(net843));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout843_A (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout844_A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout846_A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout847_A (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout848_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout849_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout850_A (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout851_A (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout852_A (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout853_A (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout854_A (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout855_A (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout856_A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout857_A (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout858_A (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout859_A (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout860_A (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout861_A (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout862_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout863_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout864_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout865_A (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout866_A (.DIODE(\u_dcg_peri.reset_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout868_A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout869_A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout870_A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout871_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout872_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout873_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout874_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout875_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout876_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout877_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout878_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout879_A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout880_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout881_A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout882_A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout883_A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout884_A (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout885_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout886_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout887_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout888_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout889_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout890_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout891_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout892_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout893_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout894_A (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout895_A (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout896_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout897_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout898_A (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout899_A (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout900_A (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout901_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout902_A (.DIODE(net903));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout903_A (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout904_A (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout905_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout906_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout907_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout908_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout909_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout910_A (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout911_A (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout912_A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout913_A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout914_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout915_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout916_A (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout917_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout918_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout919_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout921_A (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout922_A (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout923_A (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout924_A (.DIODE(_3594_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout925_A (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout926_A (.DIODE(_3594_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout927_A (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout928_A (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout929_A (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout930_A (.DIODE(_3594_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout931_A (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout932_A (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout933_A (.DIODE(_3593_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout934_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout935_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout936_A (.DIODE(_3593_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout937_A (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout938_A (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout939_A (.DIODE(net940));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout940_A (.DIODE(_3421_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout941_A (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout942_A (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout943_A (.DIODE(_3421_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout944_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout945_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout946_A (.DIODE(_3350_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout947_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout948_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout949_A (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout950_A (.DIODE(_3350_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout951_A (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout952_A (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout953_A (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout954_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout955_A (.DIODE(net956));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout956_A (.DIODE(net957));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout958_A (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout959_A (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout960_A (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout961_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout962_A (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout963_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout964_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout965_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout966_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout967_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout969_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout970_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout971_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout972_A (.DIODE(_3336_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout973_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout974_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout975_A (.DIODE(_3336_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout976_A (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout978_A (.DIODE(_3265_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout979_A (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout980_A (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout981_A (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout982_A (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout983_A (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout984_A (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout985_A (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout986_A (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout987_A (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout989_A (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout990_A (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout991_A (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout992_A (.DIODE(_2934_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout993_A (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout994_A (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout995_A (.DIODE(_2934_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout996_A (.DIODE(_2921_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout997_A (.DIODE(net1799));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout998_A (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout999_A (.DIODE(_2800_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold100_A (.DIODE(s1_wbd_dat_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold102_A (.DIODE(s1_wbd_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold103_A (.DIODE(s1_wbd_dat_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold104_A (.DIODE(s1_wbd_dat_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold106_A (.DIODE(s0_wbd_dat_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold107_A (.DIODE(s0_wbd_dat_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold108_A (.DIODE(s0_wbd_dat_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold109_A (.DIODE(s0_wbd_dat_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold10_A (.DIODE(s2_wbd_dat_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold110_A (.DIODE(m1_wbd_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold112_A (.DIODE(_3224_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold113_A (.DIODE(s0_wbd_dat_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold114_A (.DIODE(m2_wbd_adr_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold115_A (.DIODE(_3233_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold116_A (.DIODE(s0_wbd_dat_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold117_A (.DIODE(s0_wbd_dat_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold118_A (.DIODE(s0_wbd_dat_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold119_A (.DIODE(s0_wbd_dat_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold120_A (.DIODE(s0_wbd_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold121_A (.DIODE(m0_wbd_adr_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold122_A (.DIODE(m2_wbd_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold123_A (.DIODE(_2764_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold124_A (.DIODE(s0_wbd_dat_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold125_A (.DIODE(s0_wbd_dat_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold126_A (.DIODE(s0_wbd_dat_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold127_A (.DIODE(m0_wbd_adr_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold129_A (.DIODE(s0_wbd_dat_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold130_A (.DIODE(s0_wbd_dat_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold131_A (.DIODE(s0_wbd_dat_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold132_A (.DIODE(s1_wbd_dat_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold133_A (.DIODE(s1_wbd_dat_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold134_A (.DIODE(s0_wbd_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold135_A (.DIODE(m0_wbd_adr_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold137_A (.DIODE(s1_wbd_dat_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold138_A (.DIODE(s1_wbd_dat_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold139_A (.DIODE(s0_wbd_dat_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold13_A (.DIODE(_2373_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold140_A (.DIODE(s1_wbd_dat_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold141_A (.DIODE(s1_wbd_dat_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold142_A (.DIODE(m0_wbd_sel_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold143_A (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold144_A (.DIODE(m2_wbd_adr_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold146_A (.DIODE(_3230_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold147_A (.DIODE(s1_wbd_dat_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold148_A (.DIODE(s1_wbd_dat_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold149_A (.DIODE(\u_dcg_s0.u_dsync.in_data_2s[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold150_A (.DIODE(s1_wbd_dat_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold151_A (.DIODE(s1_wbd_dat_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold152_A (.DIODE(\u_s1.u_sync_wbb.m_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold154_A (.DIODE(s2_wbd_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold155_A (.DIODE(m2_wbd_dat_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold156_A (.DIODE(s1_wbd_dat_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold157_A (.DIODE(s2_wbd_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold158_A (.DIODE(m2_wbd_adr_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold160_A (.DIODE(_3227_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold161_A (.DIODE(m2_wbd_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold163_A (.DIODE(s1_wbd_dat_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold164_A (.DIODE(s2_wbd_dat_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold165_A (.DIODE(s1_wbd_dat_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold166_A (.DIODE(s2_wbd_dat_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold168_A (.DIODE(s2_wbd_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold169_A (.DIODE(s1_wbd_dat_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold16_A (.DIODE(_2372_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold170_A (.DIODE(s2_wbd_dat_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold172_A (.DIODE(m1_wbd_dat_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold173_A (.DIODE(m0_wbd_adr_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold174_A (.DIODE(m2_wbd_dat_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold176_A (.DIODE(m1_wbd_dat_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold177_A (.DIODE(m2_wbd_dat_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold17_A (.DIODE(s2_wbd_dat_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold180_A (.DIODE(_2800_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold181_A (.DIODE(m0_wbd_adr_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold182_A (.DIODE(m2_wbd_dat_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold18_A (.DIODE(s2_wbd_dat_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold191_A (.DIODE(m2_wbd_dat_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold194_A (.DIODE(m0_wbd_dat_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold195_A (.DIODE(_3162_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold197_A (.DIODE(m0_wbd_sel_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold19_A (.DIODE(s2_wbd_dat_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold200_A (.DIODE(m2_wbd_dat_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold201_A (.DIODE(m0_wbd_sel_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold203_A (.DIODE(m0_wbd_dat_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold205_A (.DIODE(s0_wbd_dat_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold206_A (.DIODE(s0_wbd_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold207_A (.DIODE(s0_wbd_dat_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold208_A (.DIODE(m0_wbd_dat_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold209_A (.DIODE(_2769_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold210_A (.DIODE(s0_wbd_dat_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold211_A (.DIODE(s0_wbd_dat_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold212_A (.DIODE(s0_wbd_dat_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold213_A (.DIODE(m0_wbd_adr_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold214_A (.DIODE(m1_wbd_adr_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold216_A (.DIODE(s0_wbd_dat_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold217_A (.DIODE(m0_wbd_adr_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold218_A (.DIODE(m1_wbd_adr_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold219_A (.DIODE(s0_wbd_dat_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold220_A (.DIODE(m2_wbd_adr_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold222_A (.DIODE(s0_wbd_dat_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold223_A (.DIODE(m1_wbd_adr_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold225_A (.DIODE(s0_wbd_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold226_A (.DIODE(s0_wbd_dat_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold227_A (.DIODE(m1_wbd_adr_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold229_A (.DIODE(m1_wbd_dat_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold22_A (.DIODE(s2_wbd_dat_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold231_A (.DIODE(m1_wbd_dat_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold233_A (.DIODE(m0_wbd_dat_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold235_A (.DIODE(m0_wbd_adr_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold236_A (.DIODE(m2_wbd_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold237_A (.DIODE(_3214_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold238_A (.DIODE(m0_wbd_adr_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold239_A (.DIODE(m1_wbd_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold23_A (.DIODE(s2_wbd_dat_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold241_A (.DIODE(m0_wbd_dat_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold242_A (.DIODE(m2_wbd_dat_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold243_A (.DIODE(_3188_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold244_A (.DIODE(m0_wbd_adr_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold246_A (.DIODE(m1_wbd_dat_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold248_A (.DIODE(m2_wbd_adr_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold24_A (.DIODE(s2_wbd_dat_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold250_A (.DIODE(m0_wbd_sel_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold251_A (.DIODE(m0_wbd_dat_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold252_A (.DIODE(_3216_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold253_A (.DIODE(m0_wbd_sel_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold254_A (.DIODE(m0_wbd_adr_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold255_A (.DIODE(m1_wbd_adr_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold256_A (.DIODE(s1_wbd_dat_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold257_A (.DIODE(m0_wbd_adr_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold258_A (.DIODE(m0_wbd_adr_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold259_A (.DIODE(m2_wbd_dat_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold260_A (.DIODE(m1_wbd_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold262_A (.DIODE(m1_wbd_dat_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold263_A (.DIODE(_2998_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold264_A (.DIODE(m2_wbd_dat_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold265_A (.DIODE(s1_wbd_dat_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold266_A (.DIODE(m1_wbd_dat_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold267_A (.DIODE(s1_wbd_dat_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold268_A (.DIODE(s1_wbd_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold269_A (.DIODE(m0_wbd_sel_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold26_A (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold270_A (.DIODE(s1_wbd_ack_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold271_A (.DIODE(s1_wbd_dat_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold272_A (.DIODE(s0_wbd_ack_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold273_A (.DIODE(m2_wbd_dat_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold274_A (.DIODE(m2_wbd_dat_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold275_A (.DIODE(m1_wbd_dat_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold276_A (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold277_A (.DIODE(m2_wbd_dat_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold278_A (.DIODE(m1_wbd_dat_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold279_A (.DIODE(m2_wbd_dat_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold280_A (.DIODE(m0_wbd_dat_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold282_A (.DIODE(m1_wbd_sel_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold283_A (.DIODE(s0_wbd_dat_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold284_A (.DIODE(m2_wbd_dat_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold285_A (.DIODE(m0_wbd_dat_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold286_A (.DIODE(s0_wbd_dat_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold287_A (.DIODE(m1_wbd_dat_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold288_A (.DIODE(s0_wbd_dat_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold289_A (.DIODE(m2_wbd_dat_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold28_A (.DIODE(s2_wbd_dat_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold290_A (.DIODE(m2_wbd_dat_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold291_A (.DIODE(m1_wbd_dat_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold292_A (.DIODE(_3170_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold293_A (.DIODE(s2_wbd_dat_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold294_A (.DIODE(m1_wbd_dat_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold295_A (.DIODE(m2_wbd_dat_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold296_A (.DIODE(_3179_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold297_A (.DIODE(m2_wbd_adr_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold298_A (.DIODE(m0_wbd_dat_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold299_A (.DIODE(m2_wbd_dat_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold29_A (.DIODE(s2_wbd_dat_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2_A (.DIODE(s0_wbd_dat_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold300_A (.DIODE(m1_wbd_dat_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold301_A (.DIODE(m2_wbd_dat_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold302_A (.DIODE(m2_wbd_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold303_A (.DIODE(_2873_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold304_A (.DIODE(s2_wbd_dat_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold305_A (.DIODE(m2_wbd_sel_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold306_A (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold307_A (.DIODE(m1_wbd_dat_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold308_A (.DIODE(m1_wbd_sel_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold309_A (.DIODE(m1_wbd_adr_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold310_A (.DIODE(m2_wbd_sel_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold311_A (.DIODE(m2_wbd_dat_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold312_A (.DIODE(s2_wbd_ack_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold313_A (.DIODE(m1_wbd_adr_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold314_A (.DIODE(m1_wbd_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold315_A (.DIODE(m2_wbd_adr_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold316_A (.DIODE(m0_wbd_adr_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold31_A (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold32_A (.DIODE(s2_wbd_dat_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold33_A (.DIODE(s2_wbd_dat_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold34_A (.DIODE(s2_wbd_dat_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold35_A (.DIODE(s2_wbd_dat_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold36_A (.DIODE(s2_wbd_dat_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold37_A (.DIODE(s2_wbd_dat_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold38_A (.DIODE(s2_wbd_dat_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold39_A (.DIODE(s2_wbd_dat_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3_A (.DIODE(m0_wbd_adr_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold40_A (.DIODE(s2_wbd_dat_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold41_A (.DIODE(s2_wbd_dat_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold43_A (.DIODE(_2572_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold4_A (.DIODE(s0_wbd_dat_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold55_A (.DIODE(s2_wbd_dat_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold56_A (.DIODE(s2_wbd_dat_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold57_A (.DIODE(s2_wbd_dat_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold58_A (.DIODE(s2_wbd_dat_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold59_A (.DIODE(m0_wbd_adr_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold5_A (.DIODE(m1_wbd_adr_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold60_A (.DIODE(_3236_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold61_A (.DIODE(s0_wbd_dat_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold62_A (.DIODE(s0_wbd_dat_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold63_A (.DIODE(s0_wbd_dat_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold64_A (.DIODE(s0_wbd_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold65_A (.DIODE(s0_wbd_dat_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold66_A (.DIODE(m2_wbd_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold67_A (.DIODE(_3204_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold68_A (.DIODE(s0_wbd_dat_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold69_A (.DIODE(m0_wbd_adr_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold6_A (.DIODE(s2_wbd_dat_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold70_A (.DIODE(m0_wbd_adr_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold71_A (.DIODE(s0_wbd_dat_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold72_A (.DIODE(s0_wbd_dat_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold73_A (.DIODE(s0_wbd_dat_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold74_A (.DIODE(m0_wbd_adr_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold77_A (.DIODE(s1_wbd_dat_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold78_A (.DIODE(s0_wbd_dat_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold79_A (.DIODE(m0_wbd_adr_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold81_A (.DIODE(m0_wbd_adr_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold82_A (.DIODE(m2_wbd_dat_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold83_A (.DIODE(s1_wbd_dat_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold84_A (.DIODE(s1_wbd_dat_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold85_A (.DIODE(m0_wbd_adr_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold86_A (.DIODE(s1_wbd_dat_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold87_A (.DIODE(s1_wbd_dat_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold88_A (.DIODE(s1_wbd_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold89_A (.DIODE(s1_wbd_dat_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold90_A (.DIODE(s1_wbd_dat_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold91_A (.DIODE(s1_wbd_dat_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold92_A (.DIODE(s1_wbd_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold93_A (.DIODE(m0_wbd_adr_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold95_A (.DIODE(m0_wbd_adr_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold97_A (.DIODE(s1_wbd_dat_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold98_A (.DIODE(s1_wbd_dat_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold99_A (.DIODE(s1_wbd_dat_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1036_A (.DIODE(_2152_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1050_A (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1097_A (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1101_A (.DIODE(_2076_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1119_A (.DIODE(_2056_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length11_A (.DIODE(net1744));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length12_A (.DIODE(\clknet_3_0__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1403_A (.DIODE(\u_s2.u_sync_wbb.wbm_ack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length14_A (.DIODE(\clknet_3_1__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1521_A (.DIODE(m2_wbd_dat_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1530_A (.DIODE(m2_wbd_dat_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length15_A (.DIODE(\clknet_3_2__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length16_A (.DIODE(\clknet_3_2__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length17_A (.DIODE(\clknet_3_3__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length18_A (.DIODE(net1751));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length19_A (.DIODE(\clknet_3_3__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length20_A (.DIODE(\clknet_3_4__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length22_A (.DIODE(\clknet_3_4__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length26_A (.DIODE(\clknet_3_5__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length37_A (.DIODE(clknet_2_1__leaf_mclk_raw));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length554_A (.DIODE(_2746_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length9_A (.DIODE(\clknet_1_1_0_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_output129_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_output130_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_output133_A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_output134_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_output139_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_output150_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_output155_A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_output156_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_output157_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_output158_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_output159_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_output15_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_output160_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_output161_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_output162_A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_output163_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_output164_A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_output165_A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_output166_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_output167_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_output168_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_output169_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_output170_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_output171_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_output172_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_output173_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_output174_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_output175_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_output176_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_output177_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_output178_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_output179_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_output180_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_output181_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_output182_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_output183_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_output184_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_output185_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_output186_A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_output187_A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_output188_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_output189_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_output18_A (.DIODE(net1489));
 sky130_fd_sc_hd__diode_2 ANTENNA_output190_A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_output191_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_output192_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_output193_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_output194_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_output195_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_output19_A (.DIODE(net1487));
 sky130_fd_sc_hd__diode_2 ANTENNA_output203_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_output205_A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_output207_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_output20_A (.DIODE(net1485));
 sky130_fd_sc_hd__diode_2 ANTENNA_output213_A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_output214_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_output21_A (.DIODE(net1483));
 sky130_fd_sc_hd__diode_2 ANTENNA_output225_A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_output22_A (.DIODE(net1481));
 sky130_fd_sc_hd__diode_2 ANTENNA_output23_A (.DIODE(net1479));
 sky130_fd_sc_hd__diode_2 ANTENNA_output24_A (.DIODE(net1477));
 sky130_fd_sc_hd__diode_2 ANTENNA_output25_A (.DIODE(net1475));
 sky130_fd_sc_hd__diode_2 ANTENNA_output268_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_output26_A (.DIODE(net1491));
 sky130_fd_sc_hd__diode_2 ANTENNA_output270_A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_output271_A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_output276_A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_output27_A (.DIODE(net1473));
 sky130_fd_sc_hd__diode_2 ANTENNA_output281_A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_output282_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_output28_A (.DIODE(net1471));
 sky130_fd_sc_hd__diode_2 ANTENNA_output292_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_output294_A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_output296_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_output297_A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_output298_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_output29_A (.DIODE(net1469));
 sky130_fd_sc_hd__diode_2 ANTENNA_output304_A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_output307_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_output308_A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_output30_A (.DIODE(net1467));
 sky130_fd_sc_hd__diode_2 ANTENNA_output312_A (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_output313_A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_output31_A (.DIODE(net1465));
 sky130_fd_sc_hd__diode_2 ANTENNA_output321_A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_output324_A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_output325_A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_output326_A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_output327_A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_output328_A (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_output329_A (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_output32_A (.DIODE(net1463));
 sky130_fd_sc_hd__diode_2 ANTENNA_output331_A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_output333_A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_output334_A (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_output335_A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_output336_A (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_output337_A (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_output338_A (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_output339_A (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_output33_A (.DIODE(net1461));
 sky130_fd_sc_hd__diode_2 ANTENNA_output340_A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_output341_A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_output342_A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_output343_A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_output344_A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_output345_A (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_output346_A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_output347_A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_output348_A (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_output349_A (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_output34_A (.DIODE(net1459));
 sky130_fd_sc_hd__diode_2 ANTENNA_output351_A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_output353_A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_output354_A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_output356_A (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_output357_A (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_output358_A (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_output359_A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_A (.DIODE(net1457));
 sky130_fd_sc_hd__diode_2 ANTENNA_output360_A (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_output361_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_output362_A (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_output364_A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_output365_A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_output366_A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_output368_A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_output369_A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA_output36_A (.DIODE(net1455));
 sky130_fd_sc_hd__diode_2 ANTENNA_output370_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_output371_A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_output373_A (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_output374_A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_output375_A (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_output376_A (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_output378_A (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_output37_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_output380_A (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_output382_A (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_output383_A (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_output384_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_output385_A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_output387_A (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_output388_A (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_output389_A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_output38_A (.DIODE(net1453));
 sky130_fd_sc_hd__diode_2 ANTENNA_output390_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_output391_A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_output392_A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_output393_A (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_output394_A (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_output396_A (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_output397_A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_output398_A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_output39_A (.DIODE(net1451));
 sky130_fd_sc_hd__diode_2 ANTENNA_output402_A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_output405_A (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_output406_A (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_output407_A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_output408_A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_output409_A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_output40_A (.DIODE(net1450));
 sky130_fd_sc_hd__diode_2 ANTENNA_output410_A (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_output411_A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_output412_A (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_output414_A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_output415_A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_output416_A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_output417_A (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_output419_A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_output41_A (.DIODE(net1449));
 sky130_fd_sc_hd__diode_2 ANTENNA_output420_A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_output421_A (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_output422_A (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_output423_A (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_output424_A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_output425_A (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_output427_A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_output429_A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_output42_A (.DIODE(net1448));
 sky130_fd_sc_hd__diode_2 ANTENNA_output430_A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_output432_A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_output433_A (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_output434_A (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_output435_A (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_output436_A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_output437_A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_output438_A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_output439_A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_output43_A (.DIODE(net1447));
 sky130_fd_sc_hd__diode_2 ANTENNA_output440_A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_output443_A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_output445_A (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_output446_A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_output448_A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_output44_A (.DIODE(net1446));
 sky130_fd_sc_hd__diode_2 ANTENNA_output450_A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_output452_A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_output453_A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_output455_A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_output456_A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_output457_A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_output459_A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_A (.DIODE(net1445));
 sky130_fd_sc_hd__diode_2 ANTENNA_output461_A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_output464_A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_output465_A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_output466_A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_output467_A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_output468_A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_output469_A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_output46_A (.DIODE(net1444));
 sky130_fd_sc_hd__diode_2 ANTENNA_output472_A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_output473_A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_output474_A (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_output476_A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_output47_A (.DIODE(net1443));
 sky130_fd_sc_hd__diode_2 ANTENNA_output48_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_output49_A (.DIODE(net1442));
 sky130_fd_sc_hd__diode_2 ANTENNA_output50_A (.DIODE(net1441));
 sky130_fd_sc_hd__diode_2 ANTENNA_output51_A (.DIODE(net1440));
 sky130_fd_sc_hd__diode_2 ANTENNA_output52_A (.DIODE(net1439));
 sky130_fd_sc_hd__diode_2 ANTENNA_output53_A (.DIODE(net1438));
 sky130_fd_sc_hd__diode_2 ANTENNA_output54_A (.DIODE(net1437));
 sky130_fd_sc_hd__diode_2 ANTENNA_output55_A (.DIODE(net1434));
 sky130_fd_sc_hd__diode_2 ANTENNA_output56_A (.DIODE(net1431));
 sky130_fd_sc_hd__diode_2 ANTENNA_output57_A (.DIODE(net1428));
 sky130_fd_sc_hd__diode_2 ANTENNA_output58_A (.DIODE(net1425));
 sky130_fd_sc_hd__diode_2 ANTENNA_output59_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_output5_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_output60_A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_output61_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_output62_A (.DIODE(net1422));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net1419));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net1416));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_output6_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_split4_A (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dcg_peri.u_clkgate.u_gate_CLK  (.DIODE(net1772));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dcg_peri.u_clkgate.u_gate_GATE  (.DIODE(net1411));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dcg_riscv.u_clkgate.u_gate_CLK  (.DIODE(net1768));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dcg_riscv.u_clkgate.u_gate_GATE  (.DIODE(net1413));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dcg_s0.u_clkgate.u_gate_CLK  (.DIODE(net1768));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dcg_s0.u_clkgate.u_gate_GATE  (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dcg_s1.u_clkgate.u_gate_CLK  (.DIODE(net1767));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dcg_s1.u_clkgate.u_gate_GATE  (.DIODE(\u_dcg_s1.clk_enb ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dcg_s2.u_clkgate.u_gate_CLK  (.DIODE(net1773));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dcg_s2.u_clkgate.u_gate_GATE  (.DIODE(net1415));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[0].u_dsync0_CLK  (.DIODE(\clknet_leaf_58_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[0].u_dsync0_D  (.DIODE(\u_dcg_s0.clk_enb ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[0].u_dsync0_RESET_B  (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[0].u_dsync1_CLK  (.DIODE(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[0].u_dsync1_D  (.DIODE(\u_dsync.in_data_s[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[0].u_dsync1_RESET_B  (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[0].u_dsync2_CLK  (.DIODE(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[0].u_dsync2_RESET_B  (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[1].u_dsync0_CLK  (.DIODE(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[1].u_dsync0_D  (.DIODE(\u_dcg_s1.clk_enb ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[1].u_dsync0_RESET_B  (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[1].u_dsync1_CLK  (.DIODE(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[1].u_dsync1_RESET_B  (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[1].u_dsync2_CLK  (.DIODE(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[1].u_dsync2_RESET_B  (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[2].u_dsync0_CLK  (.DIODE(\clknet_leaf_12_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[2].u_dsync0_D  (.DIODE(net1415));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[2].u_dsync0_RESET_B  (.DIODE(net886));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[2].u_dsync1_CLK  (.DIODE(\clknet_leaf_12_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[2].u_dsync1_RESET_B  (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[2].u_dsync2_CLK  (.DIODE(\clknet_leaf_12_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[3].u_dsync0_CLK  (.DIODE(\clknet_leaf_14_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[3].u_dsync0_D  (.DIODE(net1412));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[3].u_dsync0_RESET_B  (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[3].u_dsync1_CLK  (.DIODE(\clknet_leaf_14_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[3].u_dsync2_CLK  (.DIODE(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[4].u_dsync0_CLK  (.DIODE(\clknet_leaf_15_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[4].u_dsync0_D  (.DIODE(\u_dcg_riscv.clk_enb ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[4].u_dsync1_CLK  (.DIODE(\clknet_leaf_17_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[4].u_dsync2_CLK  (.DIODE(\clknet_leaf_19_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[4].u_dsync2_RESET_B  (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[5].u_dsync0_CLK  (.DIODE(\clknet_leaf_24_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[5].u_dsync0_RESET_B  (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[5].u_dsync1_CLK  (.DIODE(\clknet_leaf_24_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[5].u_dsync1_RESET_B  (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[5].u_dsync2_CLK  (.DIODE(\clknet_leaf_24_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[6].u_dsync0_CLK  (.DIODE(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[6].u_dsync0_RESET_B  (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[6].u_dsync1_CLK  (.DIODE(\clknet_leaf_26_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[6].u_dsync1_RESET_B  (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[6].u_dsync2_CLK  (.DIODE(\clknet_leaf_26_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[6].u_dsync2_RESET_B  (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[7].u_dsync0_CLK  (.DIODE(\clknet_leaf_24_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[7].u_dsync1_CLK  (.DIODE(\clknet_leaf_25_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[7].u_dsync1_RESET_B  (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[7].u_dsync2_CLK  (.DIODE(\clknet_leaf_29_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_dsync.bus_.bit_[7].u_dsync2_RESET_B  (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rst_sync.u_buf.genblk1.u_mux_A1  (.DIODE(rst_n));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wi.clkbuf_2.u_dly0_A  (.DIODE(\u_skew_wi.clk_d1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wi.u_clkbuf_in.u_buf_A  (.DIODE(wbd_clk_int));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wi.u_mux_level_00.genblk1.u_mux_S  (.DIODE(cfg_cska_wi[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wi.u_mux_level_01.genblk1.u_mux_S  (.DIODE(cfg_cska_wi[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wi.u_mux_level_02.genblk1.u_mux_S  (.DIODE(cfg_cska_wi[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wi.u_mux_level_03.genblk1.u_mux_S  (.DIODE(cfg_cska_wi[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wi.u_mux_level_04.genblk1.u_mux_S  (.DIODE(cfg_cska_wi[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wi.u_mux_level_05.genblk1.u_mux_S  (.DIODE(cfg_cska_wi[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wi.u_mux_level_06.genblk1.u_mux_S  (.DIODE(cfg_cska_wi[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wi.u_mux_level_07.genblk1.u_mux_S  (.DIODE(cfg_cska_wi[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wi.u_mux_level_10.genblk1.u_mux_S  (.DIODE(cfg_cska_wi[1]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wi.u_mux_level_11.genblk1.u_mux_S  (.DIODE(cfg_cska_wi[1]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wi.u_mux_level_12.genblk1.u_mux_S  (.DIODE(cfg_cska_wi[1]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wi.u_mux_level_13.genblk1.u_mux_S  (.DIODE(cfg_cska_wi[1]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wi.u_mux_level_20.genblk1.u_mux_S  (.DIODE(cfg_cska_wi[2]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wi.u_mux_level_21.genblk1.u_mux_S  (.DIODE(cfg_cska_wi[2]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wi.u_mux_level_30.genblk1.u_mux_S  (.DIODE(cfg_cska_wi[3]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wi.u_tap_1.u_buf_A  (.DIODE(\u_skew_wi.clk_d1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_wbi_clkgate.u_gate_CLK  (.DIODE(clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1007_A (.DIODE(_2187_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1008_A (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1009_A (.DIODE(_2186_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1011_A (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1012_A (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1013_A (.DIODE(_2181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1014_A (.DIODE(_2179_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1015_A (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1016_A (.DIODE(_2177_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1017_A (.DIODE(_2176_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1018_A (.DIODE(_2174_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1019_A (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1020_A (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1021_A (.DIODE(_2171_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1022_A (.DIODE(_2169_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1023_A (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1024_A (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1026_A (.DIODE(_2166_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1027_A (.DIODE(_2164_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1028_A (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1029_A (.DIODE(_2162_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1030_A (.DIODE(_2161_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1031_A (.DIODE(_2159_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1032_A (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1033_A (.DIODE(_2157_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1034_A (.DIODE(_2156_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1035_A (.DIODE(_2154_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1037_A (.DIODE(_2151_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1039_A (.DIODE(_2147_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1040_A (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1041_A (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1043_A (.DIODE(_2142_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1044_A (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1045_A (.DIODE(_2141_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1046_A (.DIODE(_2139_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1047_A (.DIODE(_2137_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1048_A (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1049_A (.DIODE(_2136_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1051_A (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1052_A (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1053_A (.DIODE(_2132_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1054_A (.DIODE(_2131_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1055_A (.DIODE(_2129_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1056_A (.DIODE(_2127_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1058_A (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1059_A (.DIODE(_2122_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1060_A (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1061_A (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1062_A (.DIODE(_2121_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1064_A (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1065_A (.DIODE(_2117_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1068_A (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1069_A (.DIODE(_2112_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1070_A (.DIODE(_2111_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1071_A (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1072_A (.DIODE(_2109_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1073_A (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1075_A (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1076_A (.DIODE(_2106_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1077_A (.DIODE(_2104_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1078_A (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1079_A (.DIODE(_2102_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1080_A (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1081_A (.DIODE(_2099_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1082_A (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1083_A (.DIODE(_2097_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1084_A (.DIODE(_2096_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1085_A (.DIODE(_2094_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1086_A (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1087_A (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1089_A (.DIODE(_2091_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1090_A (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1092_A (.DIODE(_2086_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1094_A (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1095_A (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1096_A (.DIODE(_2082_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1098_A (.DIODE(_2079_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1099_A (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire10_A (.DIODE(\clknet_3_0__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1100_A (.DIODE(_2077_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1102_A (.DIODE(_2074_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1103_A (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1104_A (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1106_A (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1107_A (.DIODE(_2069_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1108_A (.DIODE(_2067_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1109_A (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1111_A (.DIODE(_2064_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1112_A (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1113_A (.DIODE(_2062_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1115_A (.DIODE(_2059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1116_A (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1117_A (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1118_A (.DIODE(_2057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1120_A (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1121_A (.DIODE(_2054_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1123_A (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1124_A (.DIODE(_2051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1126_A (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1127_A (.DIODE(_2047_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1129_A (.DIODE(net1130));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1130_A (.DIODE(_2042_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1131_A (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1132_A (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1133_A (.DIODE(_2041_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1135_A (.DIODE(net1136));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1136_A (.DIODE(_2037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1137_A (.DIODE(_2034_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1138_A (.DIODE(net1139));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1139_A (.DIODE(_2032_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1140_A (.DIODE(net1141));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1141_A (.DIODE(_2031_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1279_A (.DIODE(\u_dcg_s0.cfg_mode[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1280_A (.DIODE(\u_reg.reg_rdata[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1281_A (.DIODE(\u_reg.reg_rdata[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1282_A (.DIODE(net1283));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1284_A (.DIODE(\u_reg.reg_rdata[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1285_A (.DIODE(\u_reg.reg_rdata[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1286_A (.DIODE(net1287));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1287_A (.DIODE(\u_reg.reg_rdata[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1288_A (.DIODE(\u_reg.reg_rdata[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1291_A (.DIODE(net1292));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1292_A (.DIODE(\u_reg.reg_rdata[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1293_A (.DIODE(net1294));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1294_A (.DIODE(\u_reg.reg_rdata[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1295_A (.DIODE(\u_reg.reg_rdata[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1296_A (.DIODE(net1297));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1297_A (.DIODE(\u_reg.reg_rdata[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1298_A (.DIODE(net1299));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1299_A (.DIODE(\u_reg.reg_rdata[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1300_A (.DIODE(net1301));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1301_A (.DIODE(\u_reg.reg_rdata[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1302_A (.DIODE(net1303));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1303_A (.DIODE(\u_reg.reg_rdata[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1304_A (.DIODE(\u_reg.reg_rdata[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1306_A (.DIODE(\u_reg.reg_rdata[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1308_A (.DIODE(\u_reg.reg_rdata[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1310_A (.DIODE(\u_reg.reg_rdata[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1366_A (.DIODE(\u_s1.u_sync_wbb.wbm_lack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1367_A (.DIODE(\u_s1.u_sync_wbb.wbm_ack_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire13_A (.DIODE(\clknet_3_1__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1401_A (.DIODE(net1400));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1402_A (.DIODE(net1403));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1411_A (.DIODE(net1412));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1413_A (.DIODE(net1414));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1414_A (.DIODE(\u_dcg_riscv.clk_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1416_A (.DIODE(net1417));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1417_A (.DIODE(net1418));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1418_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1419_A (.DIODE(net1420));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1420_A (.DIODE(net1421));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1421_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1422_A (.DIODE(net1423));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1423_A (.DIODE(net1424));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1424_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1425_A (.DIODE(net1426));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1426_A (.DIODE(net1427));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1427_A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1428_A (.DIODE(net1429));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1429_A (.DIODE(net1430));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1430_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1431_A (.DIODE(net1432));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1432_A (.DIODE(net1433));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1433_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1434_A (.DIODE(net1435));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1435_A (.DIODE(net1436));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1436_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1437_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1438_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1439_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1440_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1441_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1442_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1443_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1444_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1445_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1446_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1447_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1448_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1449_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1450_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1451_A (.DIODE(net1452));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1452_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1453_A (.DIODE(net1454));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1454_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1455_A (.DIODE(net1456));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1456_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1457_A (.DIODE(net1458));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1458_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1459_A (.DIODE(net1460));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1460_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1461_A (.DIODE(net1462));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1462_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1463_A (.DIODE(net1464));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1464_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1465_A (.DIODE(net1466));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1466_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1467_A (.DIODE(net1468));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1468_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1469_A (.DIODE(net1470));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1470_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1471_A (.DIODE(net1472));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1472_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1473_A (.DIODE(net1474));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1474_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1475_A (.DIODE(net1476));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1476_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1477_A (.DIODE(net1478));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1478_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1479_A (.DIODE(net1480));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1480_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1481_A (.DIODE(net1482));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1482_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1483_A (.DIODE(net1484));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1484_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1485_A (.DIODE(net1486));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1486_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1487_A (.DIODE(net1488));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1488_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1489_A (.DIODE(net1490));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1490_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1491_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1511_A (.DIODE(net1512));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1512_A (.DIODE(s0_idle));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1513_A (.DIODE(m2_wbd_dat_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1514_A (.DIODE(m2_wbd_dat_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1515_A (.DIODE(m2_wbd_dat_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1516_A (.DIODE(m2_wbd_dat_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1517_A (.DIODE(m2_wbd_dat_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1519_A (.DIODE(m2_wbd_dat_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1522_A (.DIODE(net2041));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1524_A (.DIODE(m2_wbd_dat_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1525_A (.DIODE(m2_wbd_dat_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1532_A (.DIODE(m2_wbd_dat_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1534_A (.DIODE(m2_wbd_dat_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1535_A (.DIODE(m1_wbd_dat_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1536_A (.DIODE(m1_wbd_dat_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1537_A (.DIODE(m1_wbd_dat_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1538_A (.DIODE(m1_wbd_dat_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1539_A (.DIODE(m1_wbd_dat_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1540_A (.DIODE(m1_wbd_dat_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1541_A (.DIODE(m1_wbd_dat_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1544_A (.DIODE(net2023));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1545_A (.DIODE(net1945));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1546_A (.DIODE(m1_wbd_dat_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1547_A (.DIODE(m1_wbd_dat_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1548_A (.DIODE(m1_wbd_dat_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1549_A (.DIODE(m1_wbd_dat_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1550_A (.DIODE(net2064));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1551_A (.DIODE(m1_wbd_dat_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1552_A (.DIODE(net2008));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1553_A (.DIODE(m1_wbd_dat_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1555_A (.DIODE(m1_wbd_dat_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1556_A (.DIODE(m1_wbd_dat_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1557_A (.DIODE(m1_wbd_dat_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1558_A (.DIODE(m1_wbd_dat_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1559_A (.DIODE(m1_wbd_dat_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1560_A (.DIODE(m1_wbd_dat_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1562_A (.DIODE(m1_wbd_dat_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1563_A (.DIODE(m1_wbd_bry_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1564_A (.DIODE(m1_wbd_bl_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1565_A (.DIODE(m0_wbd_sel_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1566_A (.DIODE(m0_wbd_dat_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1567_A (.DIODE(m0_wbd_dat_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1568_A (.DIODE(net1967));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1569_A (.DIODE(m0_wbd_dat_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1570_A (.DIODE(m0_wbd_dat_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1571_A (.DIODE(net2062));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1572_A (.DIODE(m0_wbd_dat_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1574_A (.DIODE(m0_wbd_dat_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1576_A (.DIODE(net2010));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1577_A (.DIODE(net2018));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1578_A (.DIODE(m0_wbd_dat_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1579_A (.DIODE(m0_wbd_dat_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1580_A (.DIODE(m0_wbd_dat_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1581_A (.DIODE(net2075));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1582_A (.DIODE(m0_wbd_dat_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1584_A (.DIODE(m0_wbd_dat_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1585_A (.DIODE(m0_wbd_dat_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1586_A (.DIODE(m0_wbd_dat_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1587_A (.DIODE(m0_wbd_dat_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1588_A (.DIODE(m0_wbd_dat_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1589_A (.DIODE(m0_wbd_dat_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1590_A (.DIODE(m0_wbd_dat_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1591_A (.DIODE(m0_wbd_dat_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1592_A (.DIODE(m0_wbd_dat_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1593_A (.DIODE(m0_wbd_dat_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1594_A (.DIODE(m0_wbd_adr_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1595_A (.DIODE(m0_wbd_adr_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1596_A (.DIODE(m0_wbd_adr_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1598_A (.DIODE(m0_wbd_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1599_A (.DIODE(ch_data_in[99]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1600_A (.DIODE(ch_data_in[98]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1601_A (.DIODE(net1602));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1602_A (.DIODE(ch_data_in[97]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1603_A (.DIODE(net1604));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1604_A (.DIODE(ch_data_in[96]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1605_A (.DIODE(net1606));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1606_A (.DIODE(ch_data_in[95]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1607_A (.DIODE(net1608));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1608_A (.DIODE(ch_data_in[94]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1609_A (.DIODE(net1610));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1610_A (.DIODE(ch_data_in[93]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1611_A (.DIODE(net1612));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1612_A (.DIODE(ch_data_in[92]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1613_A (.DIODE(net1614));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1614_A (.DIODE(ch_data_in[91]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1615_A (.DIODE(net1616));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1616_A (.DIODE(ch_data_in[90]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1617_A (.DIODE(net1618));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1618_A (.DIODE(ch_data_in[89]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1619_A (.DIODE(net1620));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1620_A (.DIODE(ch_data_in[88]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1621_A (.DIODE(net1622));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1622_A (.DIODE(ch_data_in[87]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1623_A (.DIODE(net1624));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1624_A (.DIODE(ch_data_in[86]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1625_A (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1626_A (.DIODE(ch_data_in[85]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1627_A (.DIODE(net1628));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1628_A (.DIODE(ch_data_in[84]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1629_A (.DIODE(net1630));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1630_A (.DIODE(ch_data_in[83]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1631_A (.DIODE(net1632));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1632_A (.DIODE(ch_data_in[82]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1633_A (.DIODE(net1634));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1634_A (.DIODE(ch_data_in[81]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1635_A (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1636_A (.DIODE(ch_data_in[80]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1637_A (.DIODE(net1638));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1638_A (.DIODE(ch_data_in[79]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1639_A (.DIODE(net1640));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1640_A (.DIODE(ch_data_in[78]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1641_A (.DIODE(net1642));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1642_A (.DIODE(ch_data_in[77]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1643_A (.DIODE(ch_data_in[43]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1644_A (.DIODE(ch_data_in[42]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1645_A (.DIODE(ch_data_in[41]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1646_A (.DIODE(ch_data_in[40]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1647_A (.DIODE(ch_data_in[39]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1648_A (.DIODE(ch_data_in[38]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1649_A (.DIODE(ch_data_in[37]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1650_A (.DIODE(ch_data_in[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1651_A (.DIODE(ch_data_in[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1652_A (.DIODE(ch_data_in[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1653_A (.DIODE(ch_data_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1654_A (.DIODE(ch_data_in[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1655_A (.DIODE(ch_data_in[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1656_A (.DIODE(ch_data_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1657_A (.DIODE(ch_data_in[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1658_A (.DIODE(ch_data_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1659_A (.DIODE(ch_data_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1660_A (.DIODE(ch_data_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1661_A (.DIODE(ch_data_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1662_A (.DIODE(ch_data_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1663_A (.DIODE(net1664));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1664_A (.DIODE(ch_data_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1665_A (.DIODE(net1666));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1666_A (.DIODE(net1667));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1667_A (.DIODE(ch_data_in[157]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1668_A (.DIODE(net1669));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1669_A (.DIODE(net1670));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1670_A (.DIODE(ch_data_in[156]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1671_A (.DIODE(net1672));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1672_A (.DIODE(net1673));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1673_A (.DIODE(ch_data_in[155]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1674_A (.DIODE(net1675));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1675_A (.DIODE(net1676));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1676_A (.DIODE(ch_data_in[151]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1677_A (.DIODE(net1678));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1678_A (.DIODE(net1679));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1679_A (.DIODE(ch_data_in[150]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1680_A (.DIODE(net1681));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1681_A (.DIODE(ch_data_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1682_A (.DIODE(ch_data_in[143]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1683_A (.DIODE(ch_data_in[142]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1684_A (.DIODE(ch_data_in[141]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1685_A (.DIODE(ch_data_in[140]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1686_A (.DIODE(net1687));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1687_A (.DIODE(ch_data_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1688_A (.DIODE(ch_data_in[139]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1689_A (.DIODE(net1690));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1690_A (.DIODE(ch_data_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1691_A (.DIODE(net1692));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1692_A (.DIODE(ch_data_in[111]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1693_A (.DIODE(net1694));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1694_A (.DIODE(ch_data_in[110]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1695_A (.DIODE(net1696));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1696_A (.DIODE(ch_data_in[109]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1697_A (.DIODE(net1698));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1698_A (.DIODE(ch_data_in[108]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1699_A (.DIODE(net1700));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1700_A (.DIODE(ch_data_in[107]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1701_A (.DIODE(net1702));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1702_A (.DIODE(ch_data_in[106]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1703_A (.DIODE(net1704));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1704_A (.DIODE(ch_data_in[105]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1705_A (.DIODE(net1706));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1706_A (.DIODE(ch_data_in[104]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1707_A (.DIODE(net1708));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1708_A (.DIODE(ch_data_in[103]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1709_A (.DIODE(net1710));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1710_A (.DIODE(ch_data_in[102]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1711_A (.DIODE(net1712));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1712_A (.DIODE(ch_data_in[101]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1713_A (.DIODE(net1714));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1714_A (.DIODE(ch_data_in[100]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1715_A (.DIODE(ch_clk_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1716_A (.DIODE(ch_clk_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1_A (.DIODE(net1734));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire21_A (.DIODE(net1754));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire23_A (.DIODE(net1758));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire24_A (.DIODE(net1757));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire25_A (.DIODE(\clknet_3_5__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire27_A (.DIODE(\clknet_3_7__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire28_A (.DIODE(\clknet_3_7__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire29_A (.DIODE(net1762));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2_A (.DIODE(net1735));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire30_A (.DIODE(net1763));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire31_A (.DIODE(mclk_raw));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire32_A (.DIODE(clknet_0_mclk_raw));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire33_A (.DIODE(clknet_0_mclk_raw));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire34_A (.DIODE(net1767));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire36_A (.DIODE(net1769));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire38_A (.DIODE(clknet_2_2__leaf_mclk_raw));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire39_A (.DIODE(clknet_2_2__leaf_mclk_raw));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire3_A (.DIODE(\u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire40_A (.DIODE(net1773));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire41_A (.DIODE(clknet_2_3__leaf_mclk_raw));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire479_A (.DIODE(_3557_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire480_A (.DIODE(_3553_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire485_A (.DIODE(_3478_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire4_A (.DIODE(\clknet_0_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire510_A (.DIODE(_2783_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire511_A (.DIODE(_2782_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire512_A (.DIODE(_2781_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire515_A (.DIODE(_3586_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire517_A (.DIODE(_3584_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire519_A (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire551_A (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire552_A (.DIODE(_2773_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire553_A (.DIODE(_2752_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire555_A (.DIODE(_2745_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire558_A (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire559_A (.DIODE(_2740_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire560_A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire561_A (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire572_A (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire573_A (.DIODE(\u_dcg_s0.clk_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire585_A (.DIODE(net1885));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire591_A (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire5_A (.DIODE(\clknet_0_u_dsync.out_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire615_A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire628_A (.DIODE(_2024_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire629_A (.DIODE(_1963_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire631_A (.DIODE(_3248_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire632_A (.DIODE(_3245_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire633_A (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire635_A (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire636_A (.DIODE(net1833));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire637_A (.DIODE(net1888));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire638_A (.DIODE(net1919));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire639_A (.DIODE(net1933));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire641_A (.DIODE(_3219_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire642_A (.DIODE(net2014));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire643_A (.DIODE(_3212_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire644_A (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire645_A (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire647_A (.DIODE(net1840));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire649_A (.DIODE(_3200_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire650_A (.DIODE(_3197_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire651_A (.DIODE(_3193_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire652_A (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire654_A (.DIODE(net2020));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire655_A (.DIODE(_3185_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire656_A (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire657_A (.DIODE(net2073));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire661_A (.DIODE(net2069));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire662_A (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire663_A (.DIODE(net1968));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire666_A (.DIODE(_3155_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire667_A (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire669_A (.DIODE(net2053));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire670_A (.DIODE(_3147_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire671_A (.DIODE(_3145_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire672_A (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire673_A (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire674_A (.DIODE(_3140_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire675_A (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire676_A (.DIODE(net1916));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire677_A (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire678_A (.DIODE(net2083));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire679_A (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire680_A (.DIODE(_2871_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire682_A (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire683_A (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire686_A (.DIODE(_2803_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire688_A (.DIODE(net1986));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire690_A (.DIODE(net1896));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire693_A (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire694_A (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire695_A (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire696_A (.DIODE(_2755_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire697_A (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire699_A (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire703_A (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire705_A (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire708_A (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire709_A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire710_A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire719_A (.DIODE(_1970_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire720_A (.DIODE(_1967_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire725_A (.DIODE(_1953_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire726_A (.DIODE(_1944_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire737_A (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire738_A (.DIODE(_1719_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire783_A (.DIODE(_1939_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire784_A (.DIODE(_1938_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire785_A (.DIODE(_1934_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire787_A (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire788_A (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire789_A (.DIODE(_1927_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire790_A (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire791_A (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire792_A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire794_A (.DIODE(_1921_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire795_A (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire8_A (.DIODE(net1741));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire920_A (.DIODE(\u_dcg_peri.reset_n ));
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_5 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_286_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_286_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_286_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_286_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_286_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_286_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_286_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_286_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_287_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_287_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_287_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_287_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_287_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_287_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_287_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_287_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_287_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_288_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_288_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_288_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_288_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_288_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_288_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_288_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_288_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_288_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_288_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_288_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_288_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_288_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_289_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_289_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_289_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_289_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_289_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_289_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_289_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_290_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_290_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_290_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_290_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_290_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_290_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_290_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_290_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_290_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_290_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_290_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_290_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_290_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_290_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_291_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_291_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_291_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_291_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_291_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_291_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_291_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_291_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_291_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_291_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_291_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_291_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_291_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_292_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_292_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_292_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_292_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_292_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_292_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_292_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_292_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_292_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_293_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_293_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_293_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_293_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_293_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_293_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_293_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_293_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_293_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_293_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_293_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_293_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_294_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_294_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_294_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_294_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_294_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_294_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_294_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_294_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_294_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_294_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_294_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_294_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_294_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_294_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_295_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_295_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_295_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_295_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_295_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_295_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_295_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_295_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_295_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_295_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_295_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_295_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_296_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_296_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_296_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_297_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_297_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_297_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_297_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_297_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_297_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_297_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_297_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_297_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_297_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_297_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_297_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_297_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_297_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_297_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_297_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_297_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_298_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_298_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_298_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_298_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_298_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_298_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_298_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_298_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_299_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_299_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_299_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_299_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_299_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_299_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_299_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_299_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_299_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_299_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_299_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_299_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_299_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_300_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_300_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_300_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_300_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_300_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_300_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_300_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_300_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_300_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_300_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_301_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_301_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_301_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_301_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_301_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_301_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_301_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_301_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_301_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_301_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_302_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_302_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_302_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_302_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_302_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_302_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_302_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_302_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_302_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_302_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_302_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_302_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_302_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_302_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_302_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_302_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_302_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_303_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_303_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_303_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_303_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_303_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_303_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_303_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_303_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_303_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_303_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_303_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_304_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_304_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_304_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_304_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_304_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_304_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_304_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_304_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_304_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_304_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_304_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_304_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_304_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_305_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_305_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_305_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_305_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_305_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_305_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_305_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_305_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_305_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_305_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_305_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_305_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_305_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_305_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_305_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_306_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_306_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_306_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_306_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_306_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_306_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_306_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_306_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_306_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_307_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_307_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_307_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_307_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_307_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_307_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_307_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_307_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_307_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_307_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_307_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_307_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_308_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_308_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_308_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_308_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_308_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_308_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_308_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_308_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_308_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_308_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_308_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_308_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_308_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_308_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_308_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_309_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_309_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_309_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_309_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_309_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_309_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_309_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_309_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_309_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_309_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_309_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_309_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_309_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_310_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_310_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_310_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_310_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_310_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_310_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_310_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_310_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_310_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_310_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_310_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_310_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_311_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_311_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_311_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_311_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_311_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_311_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_311_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_311_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_311_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_311_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_311_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_311_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_311_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_311_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_311_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_311_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_312_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_312_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_312_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_312_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_312_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_312_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_312_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_312_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_312_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_312_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_312_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_312_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_312_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_313_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_313_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_313_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_313_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_313_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_313_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_313_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_313_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_313_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_313_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_313_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_313_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_313_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_313_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_314_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_314_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_314_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_315_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_315_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_315_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_315_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_315_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_315_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_315_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_315_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_315_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_315_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_315_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_315_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_315_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_315_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_315_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_315_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_315_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_315_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_315_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_315_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_316_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_316_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_316_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_316_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_316_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_316_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_316_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_316_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_317_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_317_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_317_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_317_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_317_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_317_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_317_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_317_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_317_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_317_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_317_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_317_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_317_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_317_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_318_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_318_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_318_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_318_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_318_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_318_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_318_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_318_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_318_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_318_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_318_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_318_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_318_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_319_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_319_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_319_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_319_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_319_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_319_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_319_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_319_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_319_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_319_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_319_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_319_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_319_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_319_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_320_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_320_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_320_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_320_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_320_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_320_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_320_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_320_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_321_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_321_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_321_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_321_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_321_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_321_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_321_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_321_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_321_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_321_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_321_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_321_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_321_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_321_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_322_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_322_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_322_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_322_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_322_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_322_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_322_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_322_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_322_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_322_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_322_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_322_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_322_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_322_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_323_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_323_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_323_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_323_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_323_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_323_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_323_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_323_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_323_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_323_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_323_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_323_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_323_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_324_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_324_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_324_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_324_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_324_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_324_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_324_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_324_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_324_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_324_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_324_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_324_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_325_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_325_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_325_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_325_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_325_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_325_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_325_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_325_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_326_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_326_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_326_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_326_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_326_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_326_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_326_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_326_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_326_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_326_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_327_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_327_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_327_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_327_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_327_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_327_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_327_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_327_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_327_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_327_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_327_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_327_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_327_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_327_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_327_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_328_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_328_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_328_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_328_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_328_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_328_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_328_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_329_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_329_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_329_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_329_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_329_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_329_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_329_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_329_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_329_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_329_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_329_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_330_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_330_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_330_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_330_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_330_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_330_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_330_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_330_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_330_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_330_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_330_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_330_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_331_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_331_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_331_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_331_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_331_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_331_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_331_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_331_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_331_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_331_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_331_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_331_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_331_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_331_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_331_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_332_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_332_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_332_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_332_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_332_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_332_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_333_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_333_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_333_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_333_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_333_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_333_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_333_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_333_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_334_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_334_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_334_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_334_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_334_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_335_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_335_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_335_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_335_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_335_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_335_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_335_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_335_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_335_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_335_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_335_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_335_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_335_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_335_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_335_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_335_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_336_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_336_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_336_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_336_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_336_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_336_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_336_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_336_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_336_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_336_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_336_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_336_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_336_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_337_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_337_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_337_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_337_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_337_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_337_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_337_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_337_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_337_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_337_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_337_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_337_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_337_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_338_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_338_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_338_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_338_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_338_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_338_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_338_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_338_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_338_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_338_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_338_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_338_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_338_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_339_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_339_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_339_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_339_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_339_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_339_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_339_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_339_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_339_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_339_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_339_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_339_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_340_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_340_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_340_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_340_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_340_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_340_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_340_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_340_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_340_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_340_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_340_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_340_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_340_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_340_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_340_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_340_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_340_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_340_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_341_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_341_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_341_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_341_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_341_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_341_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_341_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_341_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_341_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_341_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_342_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_342_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_342_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_342_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_342_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_342_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_342_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_342_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_342_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_342_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_342_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_342_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_343_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_343_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_343_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_343_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_343_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_343_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_343_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_343_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_343_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_343_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_344_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_344_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_344_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_344_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_344_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_344_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_344_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_344_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_344_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_344_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_345_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_345_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_345_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_345_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_345_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_345_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_345_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_345_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_346_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_346_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_346_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_346_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_346_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_346_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_346_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_346_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_346_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_346_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_346_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_347_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_347_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_347_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_347_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_347_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_347_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_347_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_347_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_347_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_347_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_347_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_347_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_347_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_348_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_348_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_348_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_348_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_348_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_348_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_348_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_348_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_348_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_348_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_348_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_348_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_348_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_348_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_348_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_349_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_349_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_349_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_349_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_349_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_349_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_349_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_349_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_350_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_350_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_350_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_350_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_350_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_350_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_350_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_350_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_350_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_350_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_351_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_351_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_351_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_351_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_351_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_351_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_351_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_351_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_351_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_351_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_351_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_351_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_351_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_351_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_351_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_351_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_352_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_352_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_352_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_352_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_352_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_352_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_352_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_352_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_352_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_352_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_353_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_353_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_353_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_353_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_353_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_353_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_353_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_353_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_353_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_353_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_353_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_353_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_353_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_353_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_353_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_353_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_353_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_354_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_354_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_354_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_354_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_354_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_354_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_354_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_354_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_354_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_354_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_354_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_354_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_354_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_354_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_354_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_354_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_354_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_354_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_355_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_355_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_355_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_355_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_355_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_355_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_355_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_355_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_355_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_355_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_355_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_355_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_355_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_355_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_355_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_355_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_355_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_355_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_355_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_355_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_355_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_355_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_356_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_356_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_356_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_356_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_356_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_356_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_356_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_356_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_356_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_356_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_357_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_357_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_357_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_357_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_357_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_357_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_357_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_357_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_357_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_358_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_358_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_358_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_358_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_358_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_358_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_358_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_358_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_358_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_358_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_358_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_358_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_358_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_358_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_358_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_359_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_359_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_359_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_359_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_359_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_359_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_359_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_359_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_359_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_359_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_359_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_360_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_360_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_360_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_360_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_360_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_360_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_360_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_360_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_360_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_360_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_360_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_360_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_360_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_360_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_361_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_361_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_361_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_361_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_361_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_361_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_361_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_361_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_361_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_361_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_362_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_362_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_362_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_362_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_362_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_362_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_362_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_362_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_363_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_363_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_363_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_363_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_363_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_363_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_363_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_363_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_363_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_363_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_363_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_363_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_363_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_364_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_364_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_364_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_364_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_364_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_364_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_365_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_365_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_365_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_365_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_365_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_365_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_365_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_365_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_365_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_365_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_366_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_366_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_366_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_366_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_366_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_366_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_366_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_366_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_366_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_367_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_367_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_367_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_367_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_367_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_367_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_367_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_367_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_367_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_367_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_367_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_367_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_367_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_367_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_367_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_367_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_367_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_368_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_368_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_368_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_368_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_368_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_368_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_368_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_368_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_368_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_368_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_368_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_368_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_369_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_369_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_369_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_369_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_369_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_369_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_369_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_369_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_369_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_369_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_369_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_369_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_369_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_369_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_369_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_369_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_369_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_370_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_370_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_370_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_370_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_370_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_370_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_370_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_370_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_370_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_370_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_370_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_370_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_370_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_370_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_370_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_371_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_371_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_371_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_371_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_371_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_371_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_371_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_371_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_371_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_371_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_371_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_372_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_372_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_372_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_372_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_372_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_372_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_372_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_372_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_373_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_373_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_373_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_373_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_373_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_373_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_373_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_373_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_373_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_373_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_373_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_373_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_374_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_374_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_374_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_374_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_374_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_374_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_374_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_374_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_374_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_374_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_374_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_374_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_374_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_374_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_374_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_375_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_375_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_375_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_375_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_375_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_375_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_375_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_375_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_375_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_375_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_375_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_375_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_375_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_375_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_375_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_376_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_376_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_376_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_376_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_376_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_376_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_376_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_376_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_376_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_376_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_376_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_377_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_377_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_377_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_377_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_377_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_377_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_377_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_377_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_377_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_377_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_377_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_377_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_377_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_377_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_377_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_378_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_378_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_378_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_378_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_378_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_378_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_378_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_378_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_378_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_378_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_378_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_378_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_378_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_379_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_379_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_379_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_379_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_379_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_379_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_379_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_379_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_379_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_379_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_379_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_380_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_380_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_380_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_380_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_380_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_380_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_381_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_381_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_381_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_381_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_381_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_381_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_381_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_381_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_382_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_382_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_382_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_382_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_382_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_382_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_382_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_382_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_382_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_383_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_383_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_383_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_383_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_383_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_383_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_383_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_383_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_383_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_383_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_383_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_383_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_383_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_383_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_383_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_383_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_383_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_383_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_384_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_384_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_384_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_384_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_384_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_384_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_384_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_384_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_384_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_384_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_385_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_385_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_385_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_385_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_385_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_385_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_385_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_385_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_385_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_386_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_386_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_386_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_386_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_386_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_386_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_386_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_386_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_386_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_386_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_386_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_386_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_386_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_386_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_386_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_386_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_386_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_386_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_386_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_386_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_386_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_386_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_386_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_387_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_387_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_387_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_387_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_387_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_387_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_387_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_387_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_387_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_388_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_388_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_388_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_388_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_388_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_388_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_388_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_388_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_388_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_388_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_388_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_389_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_389_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_389_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_389_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_389_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_389_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_389_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_389_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_389_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_389_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_389_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_389_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_389_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_390_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_390_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_390_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_390_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_390_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_390_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_390_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_390_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_390_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_390_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_390_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_390_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_390_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_390_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_391_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_391_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_391_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_391_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_391_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_391_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_391_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_391_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_391_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_392_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_392_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_392_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_392_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_392_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_392_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_392_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_392_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_392_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_393_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_393_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_393_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_393_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_393_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_393_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_393_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_393_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_393_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_393_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_393_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_394_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_394_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_394_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_394_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_394_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_394_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_394_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_394_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_394_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_394_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_394_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_394_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_394_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_395_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_395_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_395_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_395_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_395_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_395_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_395_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_395_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_395_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_395_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_395_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_395_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_396_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_396_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_396_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_396_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_396_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_396_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_396_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_396_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_396_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_396_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_396_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_396_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_396_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_396_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_396_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_396_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_396_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_396_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_396_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_396_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_396_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_396_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_397_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_397_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_397_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_397_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_397_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_397_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_397_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_397_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_397_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_397_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_397_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_397_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_397_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_397_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_397_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_397_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_397_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_397_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_397_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_397_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_397_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_397_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_397_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_397_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_398_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_398_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_398_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_398_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_398_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_398_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_398_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_398_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_398_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_398_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_398_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_398_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_398_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_398_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_398_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_398_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_398_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_399_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_399_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_399_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_399_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_399_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_399_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_399_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_399_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_399_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_399_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_399_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_399_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_399_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_399_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_399_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_399_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_399_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_399_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_399_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_399_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_399_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_399_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_399_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_399_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_399_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_400_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_400_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_400_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_400_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_400_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_400_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_400_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_400_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_400_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_400_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_400_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_400_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_400_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_400_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_400_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_401_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_401_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_401_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_401_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_401_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_401_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_401_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_401_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_401_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_401_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_401_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_401_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_401_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_401_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_401_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_401_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_401_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_402_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_402_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_402_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_402_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_402_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_402_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_402_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_402_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_402_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_402_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_402_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_402_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_402_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_402_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_402_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_402_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_402_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_402_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_402_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_402_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_402_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_402_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_402_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_403_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_403_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_403_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_403_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_403_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_403_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_403_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_403_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_403_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_403_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_403_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_403_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_403_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_403_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_403_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_403_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_403_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_403_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_403_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_404_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_404_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_404_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_404_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_404_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_404_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_404_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_404_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_404_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_404_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_404_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_404_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_404_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_404_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_405_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_405_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_405_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_405_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_405_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_405_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_405_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_405_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_405_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_405_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_405_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_405_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_405_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_405_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_405_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_405_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_405_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_405_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_406_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_406_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_406_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_406_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_406_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_406_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_406_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_406_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_406_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_406_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_406_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_406_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_406_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_406_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_407_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_407_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_407_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_407_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_407_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_407_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_407_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_407_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_407_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_407_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_407_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_407_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_407_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_407_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_407_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_407_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_407_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_407_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_407_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_407_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_408_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_408_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_408_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_408_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_408_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_408_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_408_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_408_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_408_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_408_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_408_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_408_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_408_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_408_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_408_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_408_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_409_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_409_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_409_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_409_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_409_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_409_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_409_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_409_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_409_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_409_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_409_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_409_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_409_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_409_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_409_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_409_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_409_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_409_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_409_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_409_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_409_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_409_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_409_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_410_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_410_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_410_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_410_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_410_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_410_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_410_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_410_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_410_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_410_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_410_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_410_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_410_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_410_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_410_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_410_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_410_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_410_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_410_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_410_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_410_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_411_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_411_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_411_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_411_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_411_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_411_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_411_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_411_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_411_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_411_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_411_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_411_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_411_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_411_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_411_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_411_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_411_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_411_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_411_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_411_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_411_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_411_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_411_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_411_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_411_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_411_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_411_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_411_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_412_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_412_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_412_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_412_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_412_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_412_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_412_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_412_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_412_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_412_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_412_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_412_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_412_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_412_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_412_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_412_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_412_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_413_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_413_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_413_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_413_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_413_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_413_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_413_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_413_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_413_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_413_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_413_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_413_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_413_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_414_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_414_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_414_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_414_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_414_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_414_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_414_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_414_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_414_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_414_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_414_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_415_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_415_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_415_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_415_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_415_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_415_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_415_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_415_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_415_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_415_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_415_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_415_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_415_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_415_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_416_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_416_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_416_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_416_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_416_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_416_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_416_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_416_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_416_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_417_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_417_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_417_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_417_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_417_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_417_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_417_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_417_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_417_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_417_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_417_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_417_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_417_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_417_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_417_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_417_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_417_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_417_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_417_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_417_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_417_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_418_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_418_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_418_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_418_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_418_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_418_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_418_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_418_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_418_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_418_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_418_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_418_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_418_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_419_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_419_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_419_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_419_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_419_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_419_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_419_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_419_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_419_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_419_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_419_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_419_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_419_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_419_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_419_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_419_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_420_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_420_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_420_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_420_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_420_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_420_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_420_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_420_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_420_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_420_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_420_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_420_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_420_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_420_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_421_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_421_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_421_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_421_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_421_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_421_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_421_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_421_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_421_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_421_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_421_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_421_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_421_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_421_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_421_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_421_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_421_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_421_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_421_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_421_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_421_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_421_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_421_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_421_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_421_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_421_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_421_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_421_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_421_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_422_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_422_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_422_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_422_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_422_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_422_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_422_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_422_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_422_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_422_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_422_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_422_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_422_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_422_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_422_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_422_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_422_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_423_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_423_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_423_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_423_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_423_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_423_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_423_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_423_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_423_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_423_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_423_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_423_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_423_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_423_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_423_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_423_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_423_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_423_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_423_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_423_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_423_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_423_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_423_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_423_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_423_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_423_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_424_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_424_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_424_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_424_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_424_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_424_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_424_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_424_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_424_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_424_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_424_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_424_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_424_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_424_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_424_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_424_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_424_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_424_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_425_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_425_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_425_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_425_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_425_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_425_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_425_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_425_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_425_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_425_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_425_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_425_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_425_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_425_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_425_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_425_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_425_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_425_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_425_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_425_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_425_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_425_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_426_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_426_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_426_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_426_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_426_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_426_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_426_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_426_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_426_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_426_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_426_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_426_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_426_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_426_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_426_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_426_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_426_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_426_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_426_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_426_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_426_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_426_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_427_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_427_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_427_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_427_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_427_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_427_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_427_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_427_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_427_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_427_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_427_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_427_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_427_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_427_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_427_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_427_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_427_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_427_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_427_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_427_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_427_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_427_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_427_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_427_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_428_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_428_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_428_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_428_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_428_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_428_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_428_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_428_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_428_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_428_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_428_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_428_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_428_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_429_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_429_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_429_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_429_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_429_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_429_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_429_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_429_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_429_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_429_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_429_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_429_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_429_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_429_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_429_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_429_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_429_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_429_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_429_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_429_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_429_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_429_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_429_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_429_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_429_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_429_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_429_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_429_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_429_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_430_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_430_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_430_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_430_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_430_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_430_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_430_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_430_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_430_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_430_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_431_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_431_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_431_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_431_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_431_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_431_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_431_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_431_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_431_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_431_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_431_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_431_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_431_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_431_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_432_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_432_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_432_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_432_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_432_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_432_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_432_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_432_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_432_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_432_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_432_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_432_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_432_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_432_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_432_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_433_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_433_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_433_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_433_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_433_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_433_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_433_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_433_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_433_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_433_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_433_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_433_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_433_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_433_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_433_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_433_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_433_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_433_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_433_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_433_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_433_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_433_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_433_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_433_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_433_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_433_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_433_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_434_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_434_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_434_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_434_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_434_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_434_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_434_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_434_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_434_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_434_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_434_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_434_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_434_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_434_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_434_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_434_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_435_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_435_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_435_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_435_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_435_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_435_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_435_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_435_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_435_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_435_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_435_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_435_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_435_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_436_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_436_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_436_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_436_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_436_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_436_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_436_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_436_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_436_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_436_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_436_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_436_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_436_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_436_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_436_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_437_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_437_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_437_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_437_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_437_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_437_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_437_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_437_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_437_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_437_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_437_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_437_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_437_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_437_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_437_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_437_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_437_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_437_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_437_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_437_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_437_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_437_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_437_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_437_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_437_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_437_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_437_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_437_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_438_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_438_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_438_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_438_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_438_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_438_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_438_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_438_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_438_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_438_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_438_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_438_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_438_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_438_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_438_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_438_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_438_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_438_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_439_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_439_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_439_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_439_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_439_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_439_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_439_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_439_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_439_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_439_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_439_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_439_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_439_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_439_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_439_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_439_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_439_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_439_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_439_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_440_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_440_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_440_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_440_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_440_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_440_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_440_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_440_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_440_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_440_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_440_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_440_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_440_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_440_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_440_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_440_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_440_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_440_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_440_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_440_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_441_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_441_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_441_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_441_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_441_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_441_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_441_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_441_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_441_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_441_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_441_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_441_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_441_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_442_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_442_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_442_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_442_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_442_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_442_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_442_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_442_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_442_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_442_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_442_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_442_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_442_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_443_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_443_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_443_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_443_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_443_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_443_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_443_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_443_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_443_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_443_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_443_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_444_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_444_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_444_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_444_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_444_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_444_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_444_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_444_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_444_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_444_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_444_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_444_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_444_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_445_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_445_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_445_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_445_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_445_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_445_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_445_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_445_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_445_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_445_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_445_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_445_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_445_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_445_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_445_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_445_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_445_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_446_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_446_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_446_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_446_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_446_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_446_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_446_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_446_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_446_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_446_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_446_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_446_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_446_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_446_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_446_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_447_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_447_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_447_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_447_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_447_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_447_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_447_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_447_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_447_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_447_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_447_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_447_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_447_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_447_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_447_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_447_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_447_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_447_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_447_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_447_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_447_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_447_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_447_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_447_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_447_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_448_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_448_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_448_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_448_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_448_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_448_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_448_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_448_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_448_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_448_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_448_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_448_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_448_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_448_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_448_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_448_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_448_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_448_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_448_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_448_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_448_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_448_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_448_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_448_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_449_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_449_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_449_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_449_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_449_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_449_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_449_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_449_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_449_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_449_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_449_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_449_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_449_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_449_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_449_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_449_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_449_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_449_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_449_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_449_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_449_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_449_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_449_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_449_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_450_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_450_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_450_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_450_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_450_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_450_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_450_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_450_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_450_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_450_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_450_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_450_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_450_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_450_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_450_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_450_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_450_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_450_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_451_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_451_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_451_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_451_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_451_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_451_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_451_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_451_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_451_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_451_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_451_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_451_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_451_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_451_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_451_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_451_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_451_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_451_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_451_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_451_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_451_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_452_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_452_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_452_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_452_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_452_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_452_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_452_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_452_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_452_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_452_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_452_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_452_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_452_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_452_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_452_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_453_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_453_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_453_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_453_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_453_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_453_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_453_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_453_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_453_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_453_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_453_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_453_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_453_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_453_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_453_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_453_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_453_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_453_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_453_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_453_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_453_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_453_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_453_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_453_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_454_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_454_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_454_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_454_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_454_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_454_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_454_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_454_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_454_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_454_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_454_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_454_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_454_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_455_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_455_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_455_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_455_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_455_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_455_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_455_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_455_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_455_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_455_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_455_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_455_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_455_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_455_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_455_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_455_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_455_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_455_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_455_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_455_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_455_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_455_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_455_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_455_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_455_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_455_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_455_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_455_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_455_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_456_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_456_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_456_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_456_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_456_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_456_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_456_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_456_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_456_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_456_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_456_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_456_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_457_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_457_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_457_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_457_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_457_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_457_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_457_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_457_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_457_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_457_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_457_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_457_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_457_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_457_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_457_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_457_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_457_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_457_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_457_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_457_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_457_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_457_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_457_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_457_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_457_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_457_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_457_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_457_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_457_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_458_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_458_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_458_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_458_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_458_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_458_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_458_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_458_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_458_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_458_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_458_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_458_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_458_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_458_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_458_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_459_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_459_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_459_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_459_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_459_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_459_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_459_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_459_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_459_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_459_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_459_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_459_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_459_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_459_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_459_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_459_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_459_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_459_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_459_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_459_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_459_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_459_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_459_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_459_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_459_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_460_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_460_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_460_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_460_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_460_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_460_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_460_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_460_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_460_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_460_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_460_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_460_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_460_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_460_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_460_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_460_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_460_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_460_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_460_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_460_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_460_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_460_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_460_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_460_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_460_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_461_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_461_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_461_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_461_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_461_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_461_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_461_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_461_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_461_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_461_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_461_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_461_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_461_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_461_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_461_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_461_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_461_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_461_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_461_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_461_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_461_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_461_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_461_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_461_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_461_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_461_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_461_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_461_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_461_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_462_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_462_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_462_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_462_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_462_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_462_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_462_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_462_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_462_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_462_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_462_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_462_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_462_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_462_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_462_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_462_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_462_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_462_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_462_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_463_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_463_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_463_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_463_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_463_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_463_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_463_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_463_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_463_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_463_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_463_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_463_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_463_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_463_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_463_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_463_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_463_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_464_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_464_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_464_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_464_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_464_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_464_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_464_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_464_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_464_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_464_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_464_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_464_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_464_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_464_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_465_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_465_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_465_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_465_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_465_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_465_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_465_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_465_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_465_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_465_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_465_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_465_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_465_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_465_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_465_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_466_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_466_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_466_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_466_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_466_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_466_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_466_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_466_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_466_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_466_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_466_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_466_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_466_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_466_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_466_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_466_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_466_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_466_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_466_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_466_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_466_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_466_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_466_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_466_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_467_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_467_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_467_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_467_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_467_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_467_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_467_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_467_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_467_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_467_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_467_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_467_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_467_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_467_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_467_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_467_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_467_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_467_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_467_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_467_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_467_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_468_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_468_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_468_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_468_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_468_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_468_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_468_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_468_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_468_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_468_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_468_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_468_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_468_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_468_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_468_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_468_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_469_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_469_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_469_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_469_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_469_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_469_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_469_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_469_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_469_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_469_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_469_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_469_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_469_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_469_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_469_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_469_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_469_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_469_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_469_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_469_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_469_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_469_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_469_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_469_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_469_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_469_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_469_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_469_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_469_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_469_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_469_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_470_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_470_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_470_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_470_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_470_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_470_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_470_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_470_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_470_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_470_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_470_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_470_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_470_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_470_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_470_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_470_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_471_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_471_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_472_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_472_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_472_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_472_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_472_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_472_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_472_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_472_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_472_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_472_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_472_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_472_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_472_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_472_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_472_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_473_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_473_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_473_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_473_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_473_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_473_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_473_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_473_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_473_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_473_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_473_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_474_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_474_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_474_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_474_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_474_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_474_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_474_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_474_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_474_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_474_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_474_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_474_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_474_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_474_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_474_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_474_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_474_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_475_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_475_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_475_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_475_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_475_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_475_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_475_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_475_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_475_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_475_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_476_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_476_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_476_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_476_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_476_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_476_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_476_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_476_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_476_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_476_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_477_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_477_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_477_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_477_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_477_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_477_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_477_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_477_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_477_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_477_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_478_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_478_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_478_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_478_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_478_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_478_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_478_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_478_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_478_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_478_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_478_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_478_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_479_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_479_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_479_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_479_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_479_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_479_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_479_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_480_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_480_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_480_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_480_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_480_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_481_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_481_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_481_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_481_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_481_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_481_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_481_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_481_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_481_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_481_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_481_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_481_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_481_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_481_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_482_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_482_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_482_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_482_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_482_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_482_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_482_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_482_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_482_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_482_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_483_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_483_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_483_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_483_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_483_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_483_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_483_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_483_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_483_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_483_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_483_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_483_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_484_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_484_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_484_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_484_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_484_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_484_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_485_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_485_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_485_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_485_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_485_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_485_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_485_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_485_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_485_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_485_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_486_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_486_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_486_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_486_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_486_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_487_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_487_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_487_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_487_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_487_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_487_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_487_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_487_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_487_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_487_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_487_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_487_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_488_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_488_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_488_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_488_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_488_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_488_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_488_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_488_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_488_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_488_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_488_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_488_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_488_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_488_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_488_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_488_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_488_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_489_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_489_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_489_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_489_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_489_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_489_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_489_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_489_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_489_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_489_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_489_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_489_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_489_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_489_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_489_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_489_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_490_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_490_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_490_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_490_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_490_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_490_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_490_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_490_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_490_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_490_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_490_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_490_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_491_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_491_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_491_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_491_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_491_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_491_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_491_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_491_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_491_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_492_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_492_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_492_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_492_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_492_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_492_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_492_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_492_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_492_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_493_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_493_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_493_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_493_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_493_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_493_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_493_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_493_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_493_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_493_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_493_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_493_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_493_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_493_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_493_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_494_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_494_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_494_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_494_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_494_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_494_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_494_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_494_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_494_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_494_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_494_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_494_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_494_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_495_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_495_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_495_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_495_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_495_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_495_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_495_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_495_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_495_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_495_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_495_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_495_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_495_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_495_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_496_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_496_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_496_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_496_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_496_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_496_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_496_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_496_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_496_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_496_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_496_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_497_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_497_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_497_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_497_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_497_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_497_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_497_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_497_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_498_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_499_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_499_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_499_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_499_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_499_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_499_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_499_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_499_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_499_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_500_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_500_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_500_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_500_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_500_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_500_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_500_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_500_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_500_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_500_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_500_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_500_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_500_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_501_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_501_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_501_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_501_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_501_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_501_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_501_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_501_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_501_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_501_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_501_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_501_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_501_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_502_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_502_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_502_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_502_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_502_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_502_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_502_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_502_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_502_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_502_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_502_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_502_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_502_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_502_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_502_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_502_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_502_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_503_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_503_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_503_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_503_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_503_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_503_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_503_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_503_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_503_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_503_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_503_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_503_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_503_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_504_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_504_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_504_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_504_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_504_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_504_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_504_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_504_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_504_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_504_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_504_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_505_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_505_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_505_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_505_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_505_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_505_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_505_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_505_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_505_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_505_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_505_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_505_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_505_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_505_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_506_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_506_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_506_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_506_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_506_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_506_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_506_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_506_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_506_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_506_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_506_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_506_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_506_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_506_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_506_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_506_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_506_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_506_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_506_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_506_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_506_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_506_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_506_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_506_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_506_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_507_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_507_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_507_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_507_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_507_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_507_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_507_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_507_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_507_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_507_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_507_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_507_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_507_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_507_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_507_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_507_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_507_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_507_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_507_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_507_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_507_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_507_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_507_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_507_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_507_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_507_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_507_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_507_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_508_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_508_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_508_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_508_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_508_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_508_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_508_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_508_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_508_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_508_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_508_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_508_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_508_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_508_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_508_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_508_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_508_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_508_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_508_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_508_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_508_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_508_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_509_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_509_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_509_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_509_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_509_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_509_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_509_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_509_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_509_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_509_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_509_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_509_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_509_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_509_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_509_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_509_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_509_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_509_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_509_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_509_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_509_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_509_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_509_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_509_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_509_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_509_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_510_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_510_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_510_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_510_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_510_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_510_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_510_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_510_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_510_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_510_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_510_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_510_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_510_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_510_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_510_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_510_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_510_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_510_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_510_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_510_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_510_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_510_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_510_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_510_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_510_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_510_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_510_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_510_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_510_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_511_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_511_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_511_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_511_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_511_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_511_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_511_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_511_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_511_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_511_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_511_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_511_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_511_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_511_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_511_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_511_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_511_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_511_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_511_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_511_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_511_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_511_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_511_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_511_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_511_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_511_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_512_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_512_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_512_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_512_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_512_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_512_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_512_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_512_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_512_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_512_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_512_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_512_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_512_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_512_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_512_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_512_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_512_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_512_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_512_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_512_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_512_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_512_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_512_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_512_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_512_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_512_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_512_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_512_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_513_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_513_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_513_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_513_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_513_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_513_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_513_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_513_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_513_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_513_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_513_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_513_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_513_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_513_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_513_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_513_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_513_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_513_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_513_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_513_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_513_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_513_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_513_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_513_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_513_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_513_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_514_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_514_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_514_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_514_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_514_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_514_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_514_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_514_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_514_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_514_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_514_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_514_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_514_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_514_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_514_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_514_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_514_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_514_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_514_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_514_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_514_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_514_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_514_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_515_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_515_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_515_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_515_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_515_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_515_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_515_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_515_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_515_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_515_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_515_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_515_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_515_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_515_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_515_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_515_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_515_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_515_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_515_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_515_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_515_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_515_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_515_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_515_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_515_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_515_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_515_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_515_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_516_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_516_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_516_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_516_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_516_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_516_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_516_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_516_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_516_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_516_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_516_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_516_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_516_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_516_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_516_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_516_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_516_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_516_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_516_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_516_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_516_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_516_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_516_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_516_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_516_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_516_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_516_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_516_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_516_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_516_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_517_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_517_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_517_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_517_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_517_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_517_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_517_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_517_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_517_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_517_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_517_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_517_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_517_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_517_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_517_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_517_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_517_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_517_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_517_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_518_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_518_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_518_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_518_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_518_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_518_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_518_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_518_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_518_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_518_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_518_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_518_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_518_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_518_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_518_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_518_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_518_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_518_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_518_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_518_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_518_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_518_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_518_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_518_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_518_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_518_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_518_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_518_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_518_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_519_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_519_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_519_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_519_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_519_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_519_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_519_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_519_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_519_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_519_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_519_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_519_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_519_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_519_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_519_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_519_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_519_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_519_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_519_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_519_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_519_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_519_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_519_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_519_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_519_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_519_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_519_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_519_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_519_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_519_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_520_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_520_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_520_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_520_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_520_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_520_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_520_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_520_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_520_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_520_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_520_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_520_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_520_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_520_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_520_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_520_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_520_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_520_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_520_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_520_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_520_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_520_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_520_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_520_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_520_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_521_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_521_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_521_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_521_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_521_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_521_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_521_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_521_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_521_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_521_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_521_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_521_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_521_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_521_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_521_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_521_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_521_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_521_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_521_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_521_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_521_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_521_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_521_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_521_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_521_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_521_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_521_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_521_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_522_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_522_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_522_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_522_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_522_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_522_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_522_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_522_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_522_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_522_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_522_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_522_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_522_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_522_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_522_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_522_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_522_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_522_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_522_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_522_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_522_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_523_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_523_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_523_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_523_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_523_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_523_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_523_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_523_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_523_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_523_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_523_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_523_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_523_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_523_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_523_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_523_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_523_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_523_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_523_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_523_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_523_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_523_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_523_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_523_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_523_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_523_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_523_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_523_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_523_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_523_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_523_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_524_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_524_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_524_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_524_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_524_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_524_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_524_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_524_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_524_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_524_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_524_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_524_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_524_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_524_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_524_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_524_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_524_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_524_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_524_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_524_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_524_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_524_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_524_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_524_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_524_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_524_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_524_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_524_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_525_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_525_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_525_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_525_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_525_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_525_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_525_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_525_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_525_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_525_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_525_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_525_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_525_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_525_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_525_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_525_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_525_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_525_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_525_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_525_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_525_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_525_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_525_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_525_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_525_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_525_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_525_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_526_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_526_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_526_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_526_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_526_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_526_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_526_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_526_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_526_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_526_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_526_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_526_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_526_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_526_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_526_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_526_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_526_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_526_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_526_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_526_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_526_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_526_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_527_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_527_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_527_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_527_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_527_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_527_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_527_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_527_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_527_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_527_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_527_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_527_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_527_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_527_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_527_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_527_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_527_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_527_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_527_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_527_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_527_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_527_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_527_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_527_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_527_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_527_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_527_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_527_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_527_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_527_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_528_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_528_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_528_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_528_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_528_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_528_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_528_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_528_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_528_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_528_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_528_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_528_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_528_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_528_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_528_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_528_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_528_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_528_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_528_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_528_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_528_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_528_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_528_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_528_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_528_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_528_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_528_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_528_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_528_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_529_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_529_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_529_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_529_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_529_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_529_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_529_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_529_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_529_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_529_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_529_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_529_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_529_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_529_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_529_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_529_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_529_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_529_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_529_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_529_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_529_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_529_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_529_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_529_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_529_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_530_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_530_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_530_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_530_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_530_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_530_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_530_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_530_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_530_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_530_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_530_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_530_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_530_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_530_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_530_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_530_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_530_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_530_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_530_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_530_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_530_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_530_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_530_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_530_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_530_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_530_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_530_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_530_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_531_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_531_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_531_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_531_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_531_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_531_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_531_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_531_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_531_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_531_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_531_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_531_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_531_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_531_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_531_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_531_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_531_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_531_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_531_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_531_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_531_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_531_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_531_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_531_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_531_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_532_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_532_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_532_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_532_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_532_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_532_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_532_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_532_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_532_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_532_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_532_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_532_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_532_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_532_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_532_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_532_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_532_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_532_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_532_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_532_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_532_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_532_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_532_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_532_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_532_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_532_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_532_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_533_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_533_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_533_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_533_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_533_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_533_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_533_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_533_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_533_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_533_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_533_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_533_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_533_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_533_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_533_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_533_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_533_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_533_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_533_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_533_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_533_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_534_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_534_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_534_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_534_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_534_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_534_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_534_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_534_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_534_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_534_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_534_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_534_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_534_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_534_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_534_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_534_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_534_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_534_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_534_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_534_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_534_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_534_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_534_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_534_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_534_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_534_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_534_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_535_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_535_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_535_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_535_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_535_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_535_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_535_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_535_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_535_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_535_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_535_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_535_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_535_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_535_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_535_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_535_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_535_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_535_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_535_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_535_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_535_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_535_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_535_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_535_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_535_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_535_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_535_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_535_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_535_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_536_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_536_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_536_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_536_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_536_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_536_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_536_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_536_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_536_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_536_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_536_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_536_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_536_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_536_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_536_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_536_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_536_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_536_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_536_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_536_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_536_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_536_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_536_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_536_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_536_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_536_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_537_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_537_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_537_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_537_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_537_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_537_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_537_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_537_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_537_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_537_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_537_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_537_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_537_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_537_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_537_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_537_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_537_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_537_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_537_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_537_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_537_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_537_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_537_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_537_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_537_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_538_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_538_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_538_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_538_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_538_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_538_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_538_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_538_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_538_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_538_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_538_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_538_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_538_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_538_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_538_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_538_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_538_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_538_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_538_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_538_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_539_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_539_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_539_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_539_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_539_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_539_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_539_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_539_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_539_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_539_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_539_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_539_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_539_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_539_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_539_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_539_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_539_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_539_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_539_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_539_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_539_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_539_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_539_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_539_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_539_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_539_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_539_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_540_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_540_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_540_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_540_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_540_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_540_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_540_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_540_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_540_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_540_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_540_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_540_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_540_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_540_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_540_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_540_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_540_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_540_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_540_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_540_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_540_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_540_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_541_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_541_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_541_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_541_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_541_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_541_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_541_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_541_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_541_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_541_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_541_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_541_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_541_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_541_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_541_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_541_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_541_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_541_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_541_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_541_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_541_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_541_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_541_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_541_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_541_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_541_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_542_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_542_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_542_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_542_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_542_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_542_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_542_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_542_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_542_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_542_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_542_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_542_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_542_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_542_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_542_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_542_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_542_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_542_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_542_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_542_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_542_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_542_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_542_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_542_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_543_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_543_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_543_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_543_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_543_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_543_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_543_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_543_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_543_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_543_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_543_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_543_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_543_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_543_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_543_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_543_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_543_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_543_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_543_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_543_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_543_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_543_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_543_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_543_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_543_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_543_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_543_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_543_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_543_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_543_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_544_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_544_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_544_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_544_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_544_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_544_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_544_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_544_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_544_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_544_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_544_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_544_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_544_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_544_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_544_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_544_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_544_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_544_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_544_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_544_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_544_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_544_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_544_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_544_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_544_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_545_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_545_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_545_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_545_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_545_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_545_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_545_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_545_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_545_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_545_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_545_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_545_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_545_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_545_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_545_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_545_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_545_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_545_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_546_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_546_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_546_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_546_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_546_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_546_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_546_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_546_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_546_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_546_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_546_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_546_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_546_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_546_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_546_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_546_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_546_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_546_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_546_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_547_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_547_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_547_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_547_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_547_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_547_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_547_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_547_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_547_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_547_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_547_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_547_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_547_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_547_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_547_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_547_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_547_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_547_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_547_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_547_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_547_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_547_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_547_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_547_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_547_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_547_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_547_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_547_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_547_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_547_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_548_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_548_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_548_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_548_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_548_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_548_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_548_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_548_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_548_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_548_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_548_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_548_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_548_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_548_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_548_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_548_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_548_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_548_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_548_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_548_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_548_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_548_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_548_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_548_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_548_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_549_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_549_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_549_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_549_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_549_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_549_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_549_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_549_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_549_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_549_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_549_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_549_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_549_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_549_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_549_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_549_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_549_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_549_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_549_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_549_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_549_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_549_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_549_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_549_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_549_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_549_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_549_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_549_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_549_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_549_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_550_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_550_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_550_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_550_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_550_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_550_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_550_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_550_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_550_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_550_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_550_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_550_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_550_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_550_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_550_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_550_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_550_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_550_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_550_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_550_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_550_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_550_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_550_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_551_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_551_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_551_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_551_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_551_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_551_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_551_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_551_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_551_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_551_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_551_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_551_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_551_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_551_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_551_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_551_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_551_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_551_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_551_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_551_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_551_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_551_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_551_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_551_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_551_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_551_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_552_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_552_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_552_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_552_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_552_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_552_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_552_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_552_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_552_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_552_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_552_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_552_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_552_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_552_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_552_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_552_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_552_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_552_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_552_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_552_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_552_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_552_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_552_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_552_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_552_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_552_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_552_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_552_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_552_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_552_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_553_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_553_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_553_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_553_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_553_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_553_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_553_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_553_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_553_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_553_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_553_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_553_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_553_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_553_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_553_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_553_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_553_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_553_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_553_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_553_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_553_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_553_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_553_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_553_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_553_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_554_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_554_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_554_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_554_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_554_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_554_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_554_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_554_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_554_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_554_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_554_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_554_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_554_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_554_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_554_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_554_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_554_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_554_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_554_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_554_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_554_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_554_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_555_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_555_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_555_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_555_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_555_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_555_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_555_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_555_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_555_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_555_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_555_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_555_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_555_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_555_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_555_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_555_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_555_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_555_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_555_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_555_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_555_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_555_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_555_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_555_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_555_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_555_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_555_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_556_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_556_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_556_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_556_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_556_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_556_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_556_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_556_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_556_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_556_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_556_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_556_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_556_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_556_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_556_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_556_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_556_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_556_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_556_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_556_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_556_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_556_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_557_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_557_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_557_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_557_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_557_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_557_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_557_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_557_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_557_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_557_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_557_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_557_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_557_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_557_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_557_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_557_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_557_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_557_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_557_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_557_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_557_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_557_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_557_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_557_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_557_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_557_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_557_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_557_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_558_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_558_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_558_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_558_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_558_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_558_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_558_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_558_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_558_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_558_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_558_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_558_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_558_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_558_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_558_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_558_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_558_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_558_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_558_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_558_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_558_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_558_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_558_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_558_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_558_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_559_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_559_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_559_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_559_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_559_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_559_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_559_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_559_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_559_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_559_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_559_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_559_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_559_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_559_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_559_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_559_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_559_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_559_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_559_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_559_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_559_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_559_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_559_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_559_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_559_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_559_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_559_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_560_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_560_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_560_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_560_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_560_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_560_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_560_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_560_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_560_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_560_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_560_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_560_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_560_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_560_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_560_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_560_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_560_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_560_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_560_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_560_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_560_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_560_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_560_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_560_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_560_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_560_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_561_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_561_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_561_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_561_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_561_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_561_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_561_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_561_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_561_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_561_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_561_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_561_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_561_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_561_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_561_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_561_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_561_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_561_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_561_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_561_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_561_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_561_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_561_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_561_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_561_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_561_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_561_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_561_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_561_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_562_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_562_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_562_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_562_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_562_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_562_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_562_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_562_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_562_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_562_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_562_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_562_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_562_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_562_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_562_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_562_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_562_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_562_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_562_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_562_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_562_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_562_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_562_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_562_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_562_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_562_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_563_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_563_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_563_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_563_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_563_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_563_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_563_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_563_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_563_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_563_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_563_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_563_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_563_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_563_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_563_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_563_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_563_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_563_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_563_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_563_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_563_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_564_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_564_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_564_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_564_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_564_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_564_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_564_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_564_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_564_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_564_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_564_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_564_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_564_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_564_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_564_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_564_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_564_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_564_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_564_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_564_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_564_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_564_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_564_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_564_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_564_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_564_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_564_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_564_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_565_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_565_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_565_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_565_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_565_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_565_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_565_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_565_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_565_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_565_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_565_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_565_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_565_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_565_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_565_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_565_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_565_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_565_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_565_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_565_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_565_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_565_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_565_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_565_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_565_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_565_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_566_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_566_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_566_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_566_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_566_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_566_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_566_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_566_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_566_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_566_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_566_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_566_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_566_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_566_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_566_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_566_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_566_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_566_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_566_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_566_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_566_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_566_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_566_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_566_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_566_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_566_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_566_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_567_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_567_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_567_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_567_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_567_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_567_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_567_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_567_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_567_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_567_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_567_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_567_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_567_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_567_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_567_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_568_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_568_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_568_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_568_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_568_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_568_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_568_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_568_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_568_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_568_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_568_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_568_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_568_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_568_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_568_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_568_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_568_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_568_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_568_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_568_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_568_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_568_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_568_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_568_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_569_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_569_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_569_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_569_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_569_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_569_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_569_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_569_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_569_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_569_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_569_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_569_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_569_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_569_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_569_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_569_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_569_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_569_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_569_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_569_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_569_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_569_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_569_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_569_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_569_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_569_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_570_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_570_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_570_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_570_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_570_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_570_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_570_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_570_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_570_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_570_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_570_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_570_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_570_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_570_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_570_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_570_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_570_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_570_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_570_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_570_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_570_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_570_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_570_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_570_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_570_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_571_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_571_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_571_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_571_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_571_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_571_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_571_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_571_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_571_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_571_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_571_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_571_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_571_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_571_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_571_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_571_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_571_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_571_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_571_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_571_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_571_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_571_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_571_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_571_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_571_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_571_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_572_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_572_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_572_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_572_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_572_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_572_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_572_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_572_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_572_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_572_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_572_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_572_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_572_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_572_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_572_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_572_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_572_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_572_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_572_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_573_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_573_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_573_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_573_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_573_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_573_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_573_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_573_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_573_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_573_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_573_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_573_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_573_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_573_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_573_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_573_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_573_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_573_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_573_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_573_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_573_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_573_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_573_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_574_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_574_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_574_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_574_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_574_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_574_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_574_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_574_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_574_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_574_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_574_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_574_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_574_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_574_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_574_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_574_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_574_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_574_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_574_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_574_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_574_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_574_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_575_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_575_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_575_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_575_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_575_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_575_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_575_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_575_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_575_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_575_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_575_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_575_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_575_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_575_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_575_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_575_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_575_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_575_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_575_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_575_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_575_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_575_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_575_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_575_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_575_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_575_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_575_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_575_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_575_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_575_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_575_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_576_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_576_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_576_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_576_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_576_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_576_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_576_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_576_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_576_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_576_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_576_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_576_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_576_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_576_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_576_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_576_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_576_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_576_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_576_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_576_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_576_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_576_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_576_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_577_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_577_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_577_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_577_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_577_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_577_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_577_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_577_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_577_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_577_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_577_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_577_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_577_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_577_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_577_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_577_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_577_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_577_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_577_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_577_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_577_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_577_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_577_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_577_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_577_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_577_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_578_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_578_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_578_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_578_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_578_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_578_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_578_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_578_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_578_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_578_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_578_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_578_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_578_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_578_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_578_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_578_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_578_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_578_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_578_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_578_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_578_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_578_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_578_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_578_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_579_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_579_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_579_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_579_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_579_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_579_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_579_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_579_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_579_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_579_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_579_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_579_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_579_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_579_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_579_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_579_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_579_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_579_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_579_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_579_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_579_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_579_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_579_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_579_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_580_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_580_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_580_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_580_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_580_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_580_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_580_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_580_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_580_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_580_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_580_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_580_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_580_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_580_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_580_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_580_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_580_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_580_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_580_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_580_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_580_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_580_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_580_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_580_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_580_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_580_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_580_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_580_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_580_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_580_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_580_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_581_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_581_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_581_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_581_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_581_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_581_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_581_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_581_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_581_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_581_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_581_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_581_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_581_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_581_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_581_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_581_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_581_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_581_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_581_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_581_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_581_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_581_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_581_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_581_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_581_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_582_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_582_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_582_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_582_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_582_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_582_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_582_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_582_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_582_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_582_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_582_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_582_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_582_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_582_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_582_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_582_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_582_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_582_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_582_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_582_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_582_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_582_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_583_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_583_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_583_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_583_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_583_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_583_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_583_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_583_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_583_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_583_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_583_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_583_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_583_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_583_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_583_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_583_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_583_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_583_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_583_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_583_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_583_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_583_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_583_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_583_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_583_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_583_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_583_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_583_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_583_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_583_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_583_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_584_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_584_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_584_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_584_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_584_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_584_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_584_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_584_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_584_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_584_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_584_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_584_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_584_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_584_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_584_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_584_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_584_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_584_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_584_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_584_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_584_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_584_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_584_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_584_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_584_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_585_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_585_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_585_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_585_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_585_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_585_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_585_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_585_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_585_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_585_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_585_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_585_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_585_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_585_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_585_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_585_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_585_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_585_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_585_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_585_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_585_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_585_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_585_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_585_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_586_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_586_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_586_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_586_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_586_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_586_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_586_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_586_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_586_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_586_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_586_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_586_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_586_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_586_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_586_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_586_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_586_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_586_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_586_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_586_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_586_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_586_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_586_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_586_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_586_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_586_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_587_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_587_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_587_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_587_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_587_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_587_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_587_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_587_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_587_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_587_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_587_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_587_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_587_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_587_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_587_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_587_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_587_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_587_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_587_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_587_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_587_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_587_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_587_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_587_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_587_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_587_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_588_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_588_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_588_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_588_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_588_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_588_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_588_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_588_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_588_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_588_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_588_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_588_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_588_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_588_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_588_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_588_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_588_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_588_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_588_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_588_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_588_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_589_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_589_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_589_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_589_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_589_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_589_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_589_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_589_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_589_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_589_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_589_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_589_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_589_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_589_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_589_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_589_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_589_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_589_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_589_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_589_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_589_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_589_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_589_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_589_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_589_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_590_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_590_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_590_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_590_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_590_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_590_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_590_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_590_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_590_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_590_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_590_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_590_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_590_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_590_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_590_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_590_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_590_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_590_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_590_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_590_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_590_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_590_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_590_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_590_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_590_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_590_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_591_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_591_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_591_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_591_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_591_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_591_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_591_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_591_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_591_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_591_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_591_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_591_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_591_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_591_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_591_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_591_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_591_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_591_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_591_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_591_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_591_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_591_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_591_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_591_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_591_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_591_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_591_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_592_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_592_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_592_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_592_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_592_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_592_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_592_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_592_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_592_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_592_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_592_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_592_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_592_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_592_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_592_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_592_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_592_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_592_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_592_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_592_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_592_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_592_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_592_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_592_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_592_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_593_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_593_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_593_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_593_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_593_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_593_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_593_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_593_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_593_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_593_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_593_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_593_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_593_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_593_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_593_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_593_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_593_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_593_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_593_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_593_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_593_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_593_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_593_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_593_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_593_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_593_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_593_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_593_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_593_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_594_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_594_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_594_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_594_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_594_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_594_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_594_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_594_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_594_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_594_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_594_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_594_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_594_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_594_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_594_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_594_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_594_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_594_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_594_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_594_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_594_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_594_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_594_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_594_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_595_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_595_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_595_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_595_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_595_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_595_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_595_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_595_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_595_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_595_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_595_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_595_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_595_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_595_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_595_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_595_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_595_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_595_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_595_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_595_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_595_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_595_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_595_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_595_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_595_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_595_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_595_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_596_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_596_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_596_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_596_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_596_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_596_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_596_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_596_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_596_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_596_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_596_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_596_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_596_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_596_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_596_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_596_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_596_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_596_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_596_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_596_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_596_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_596_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_596_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_597_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_597_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_597_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_597_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_597_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_597_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_597_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_597_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_597_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_597_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_597_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_597_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_597_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_597_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_597_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_597_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_597_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_597_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_597_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_597_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_597_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_597_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_597_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_597_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_597_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_597_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_597_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_597_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_597_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_597_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_598_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_598_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_598_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_598_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_598_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_598_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_598_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_598_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_598_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_598_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_598_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_598_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_598_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_598_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_598_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_598_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_598_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_598_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_598_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_598_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_598_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_599_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_599_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_599_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_599_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_599_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_599_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_599_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_599_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_599_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_599_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_599_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_599_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_599_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_599_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_599_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_599_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_599_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_599_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_599_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_599_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_599_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_599_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_599_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_600_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_600_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_600_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_600_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_600_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_600_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_600_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_600_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_600_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_600_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_600_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_600_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_600_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_600_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_600_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_600_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_600_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_600_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_600_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_600_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_600_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_600_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_600_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_601_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_601_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_601_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_601_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_601_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_601_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_601_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_601_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_601_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_601_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_601_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_601_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_601_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_601_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_601_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_601_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_601_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_601_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_601_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_601_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_601_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_601_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_602_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_602_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_602_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_602_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_602_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_602_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_602_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_602_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_602_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_602_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_602_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_602_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_602_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_602_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_602_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_602_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_602_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_602_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_602_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_602_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_602_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_602_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_602_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_603_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_603_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_603_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_603_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_603_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_603_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_603_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_603_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_603_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_603_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_603_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_603_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_603_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_603_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_603_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_603_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_603_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_603_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_603_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_603_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_603_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_603_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_603_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_603_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_604_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_604_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_604_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_604_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_604_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_604_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_604_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_604_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_604_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_604_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_604_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_604_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_604_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_604_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_604_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_604_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_604_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_604_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_604_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_604_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_604_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_605_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_605_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_605_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_605_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_605_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_605_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_605_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_605_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_605_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_605_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_605_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_605_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_605_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_605_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_605_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_605_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_605_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_605_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_605_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_605_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_605_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_605_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_606_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_606_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_606_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_606_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_606_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_606_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_606_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_606_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_606_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_606_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_606_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_606_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_606_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_606_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_606_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_606_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_606_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_606_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_606_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_606_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_606_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_606_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_606_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_606_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_607_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_607_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_607_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_607_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_607_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_607_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_607_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_607_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_607_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_607_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_607_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_607_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_607_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_607_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_607_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_607_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_607_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_607_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_607_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_607_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_607_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_607_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_607_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_607_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_607_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_607_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_607_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_608_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_608_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_608_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_608_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_608_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_608_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_608_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_608_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_608_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_608_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_608_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_608_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_608_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_608_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_608_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_608_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_608_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_608_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_608_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_608_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_608_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_608_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_608_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_608_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_608_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_608_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_609_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_609_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_609_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_609_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_609_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_609_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_609_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_609_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_609_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_609_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_609_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_609_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_609_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_609_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_609_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_609_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_609_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_609_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_609_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_609_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_609_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_609_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_609_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_609_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_609_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_609_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_609_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_609_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_609_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_609_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_609_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_609_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_609_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_609_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_609_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_609_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_610_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_610_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_610_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_610_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_610_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_610_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_610_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_610_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_610_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_610_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_610_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_610_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_610_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_610_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_610_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_610_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_610_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_610_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_610_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_610_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_610_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_610_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_610_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_610_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_611_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_611_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_611_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_611_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_611_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_611_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_611_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_611_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_611_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_611_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_611_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_611_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_611_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_611_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_611_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_611_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_611_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_611_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_611_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_611_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_611_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_611_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_611_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_611_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_611_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_611_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_611_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_611_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_611_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_612_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_612_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_612_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_612_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_612_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_612_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_612_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_612_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_612_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_612_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_612_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_612_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_612_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_612_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_612_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_612_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_612_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_612_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_612_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_612_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_612_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_612_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_612_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_612_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_613_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_613_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_613_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_613_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_613_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_613_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_613_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_613_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_613_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_613_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_613_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_613_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_613_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_613_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_613_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_613_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_613_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_613_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_613_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_613_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_613_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_613_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_613_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_613_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_613_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_613_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_613_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_613_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_613_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_613_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_613_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_614_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_614_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_614_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_614_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_614_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_614_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_614_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_614_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_614_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_614_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_614_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_614_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_614_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_614_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_614_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_614_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_614_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_614_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_614_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_614_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_615_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_615_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_615_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_615_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_615_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_615_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_615_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_615_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_615_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_615_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_615_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_615_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_615_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_615_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_615_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_615_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_615_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_615_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_615_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_615_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_615_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_615_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_615_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_615_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_615_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_615_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_616_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_616_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_616_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_616_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_616_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_616_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_616_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_616_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_616_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_616_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_616_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_616_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_616_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_616_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_616_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_616_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_616_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_616_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_616_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_616_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_616_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_616_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_616_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_616_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_617_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_617_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_617_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_617_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_617_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_617_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_617_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_617_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_617_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_617_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_617_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_617_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_617_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_617_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_617_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_617_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_617_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_617_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_617_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_617_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_617_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_617_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_617_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_617_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_617_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_617_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_618_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_618_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_618_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_618_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_618_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_618_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_618_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_618_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_618_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_618_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_618_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_618_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_618_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_618_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_618_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_618_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_618_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_618_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_618_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_618_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_618_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_618_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_619_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_619_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_619_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_619_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_619_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_619_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_619_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_619_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_619_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_619_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_619_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_619_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_619_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_619_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_619_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_619_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_619_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_619_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_619_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_619_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_619_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_619_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_619_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_620_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_620_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_620_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_620_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_620_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_620_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_620_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_620_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_620_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_620_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_620_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_620_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_620_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_620_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_620_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_620_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_620_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_620_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_620_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_620_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_620_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_620_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_620_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_621_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_621_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_621_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_621_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_621_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_621_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_621_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_621_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_621_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_621_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_621_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_621_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_621_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_621_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_621_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_621_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_621_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_621_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_621_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_621_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_621_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_621_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_621_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_621_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_621_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_621_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_621_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_622_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_622_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_622_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_622_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_622_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_622_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_622_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_622_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_622_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_622_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_622_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_622_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_622_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_622_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_622_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_622_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_622_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_622_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_622_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_622_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_622_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_622_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_622_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_622_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_623_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_623_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_623_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_623_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_623_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_623_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_623_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_623_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_623_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_623_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_623_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_623_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_623_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_623_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_623_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_623_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_623_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_623_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_623_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_623_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_623_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_623_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_623_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_623_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_623_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_623_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_623_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_623_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_623_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_624_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_624_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_624_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_624_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_624_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_624_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_624_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_624_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_624_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_624_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_624_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_624_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_624_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_624_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_624_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_624_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_624_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_624_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_624_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_624_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_624_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_624_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_624_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_624_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_624_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_625_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_625_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_625_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_625_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_625_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_625_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_625_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_625_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_625_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_625_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_625_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_625_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_625_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_625_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_625_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_625_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_625_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_625_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_625_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_625_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_625_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_625_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_625_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_625_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_626_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_626_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_626_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_626_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_626_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_626_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_626_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_626_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_626_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_626_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_626_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_626_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_626_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_626_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_626_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_626_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_626_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_626_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_626_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_626_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_626_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_626_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_626_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_626_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_626_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_627_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_627_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_627_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_627_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_627_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_627_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_627_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_627_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_627_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_627_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_627_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_627_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_627_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_627_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_627_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_627_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_627_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_627_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_627_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_627_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_627_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_627_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_627_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_627_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_628_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_628_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_628_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_628_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_628_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_628_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_628_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_628_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_628_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_628_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_628_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_628_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_628_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_628_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_628_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_628_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_628_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_628_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_628_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_628_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_628_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_628_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_628_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_628_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_628_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_628_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_629_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_629_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_629_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_629_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_629_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_629_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_629_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_629_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_629_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_629_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_629_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_629_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_629_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_629_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_629_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_629_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_629_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_629_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_629_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_629_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_629_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_629_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_629_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_629_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_629_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_629_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_629_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_630_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_630_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_630_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_630_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_630_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_630_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_630_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_630_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_630_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_630_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_630_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_630_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_630_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_630_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_630_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_630_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_630_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_630_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_630_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_630_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_630_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_630_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_630_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_631_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_631_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_631_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_631_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_631_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_631_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_631_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_631_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_631_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_631_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_631_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_631_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_631_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_631_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_631_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_631_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_631_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_631_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_631_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_631_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_631_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_631_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_631_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_631_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_631_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_631_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_631_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_631_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_631_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_631_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_632_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_632_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_632_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_632_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_632_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_632_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_632_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_632_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_632_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_632_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_632_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_632_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_632_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_632_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_632_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_632_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_632_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_632_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_632_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_632_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_632_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_632_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_632_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_632_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_633_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_633_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_633_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_633_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_633_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_633_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_633_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_633_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_633_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_633_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_633_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_633_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_633_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_633_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_633_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_633_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_633_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_633_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_633_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_633_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_633_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_633_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_634_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_634_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_634_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_634_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_634_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_634_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_634_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_634_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_634_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_634_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_634_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_634_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_634_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_634_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_634_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_634_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_634_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_634_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_634_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_634_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_634_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_634_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_634_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_635_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_635_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_635_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_635_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_635_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_635_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_635_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_635_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_635_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_635_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_635_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_635_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_635_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_635_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_635_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_635_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_635_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_635_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_635_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_635_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_635_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_635_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_635_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_635_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_635_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_636_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_636_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_636_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_636_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_636_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_636_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_636_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_636_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_636_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_636_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_636_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_636_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_636_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_636_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_636_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_636_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_636_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_636_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_636_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_636_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_636_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_636_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_636_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_637_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_637_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_637_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_637_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_637_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_637_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_637_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_637_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_637_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_637_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_637_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_637_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_637_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_637_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_637_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_637_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_637_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_637_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_637_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_637_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_637_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_637_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_637_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_638_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_638_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_638_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_638_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_638_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_638_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_638_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_638_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_638_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_638_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_638_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_638_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_638_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_638_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_638_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_638_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_638_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_638_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_638_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_638_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_638_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_638_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_638_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_638_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_638_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_638_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_638_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_639_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_639_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_639_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_639_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_639_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_639_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_639_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_639_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_639_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_639_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_639_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_639_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_639_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_639_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_639_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_639_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_639_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_639_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_639_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_639_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_639_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_639_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_639_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_639_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_639_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_639_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_640_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_640_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_640_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_640_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_640_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_640_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_640_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_640_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_640_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_640_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_640_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_640_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_640_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_640_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_640_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_640_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_640_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_640_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_640_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_640_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_640_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_640_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_640_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_640_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_641_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_641_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_641_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_641_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_641_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_641_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_641_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_641_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_641_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_641_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_641_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_641_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_641_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_641_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_641_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_641_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_641_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_641_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_641_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_641_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_641_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_641_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_641_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_642_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_642_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_642_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_642_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_642_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_642_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_642_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_642_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_642_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_642_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_642_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_642_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_642_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_642_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_642_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_642_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_642_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_642_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_642_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_642_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_642_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_642_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_642_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_642_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_642_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_642_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_643_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_643_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_643_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_643_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_643_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_643_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_643_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_643_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_643_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_643_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_643_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_643_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_643_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_643_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_643_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_643_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_643_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_643_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_643_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_643_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_643_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_643_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_643_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_643_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_643_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_643_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_643_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_644_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_644_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_644_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_644_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_644_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_644_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_644_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_644_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_644_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_644_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_644_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_644_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_644_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_644_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_644_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_644_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_644_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_644_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_644_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_644_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_644_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_645_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_645_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_645_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_645_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_645_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_645_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_645_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_645_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_645_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_645_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_645_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_645_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_645_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_645_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_645_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_645_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_645_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_645_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_645_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_645_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_645_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_645_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_646_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_646_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_646_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_646_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_646_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_646_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_646_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_646_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_646_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_646_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_646_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_646_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_646_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_646_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_646_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_646_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_646_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_646_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_646_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_646_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_646_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_647_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_647_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_647_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_647_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_647_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_647_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_647_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_647_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_647_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_647_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_647_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_647_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_647_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_647_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_647_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_647_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_647_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_647_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_647_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_647_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_647_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_647_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_647_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_648_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_648_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_648_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_648_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_648_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_648_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_648_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_648_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_648_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_648_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_648_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_648_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_648_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_648_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_648_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_648_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_648_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_648_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_648_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_648_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_648_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_649_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_649_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_649_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_649_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_649_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_649_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_649_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_649_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_649_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_649_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_649_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_649_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_649_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_649_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_649_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_649_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_649_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_649_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_649_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_649_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_649_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_649_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_649_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_650_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_650_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_650_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_650_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_650_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_650_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_650_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_650_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_650_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_650_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_650_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_650_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_650_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_650_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_650_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_650_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_650_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_650_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_650_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_650_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_650_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_651_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_651_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_651_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_651_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_651_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_651_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_651_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_651_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_651_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_651_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_651_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_651_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_651_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_651_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_651_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_651_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_651_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_651_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_651_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_651_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_651_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_651_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_651_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_652_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_652_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_652_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_5 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_1000 ();
 sky130_fd_sc_hd__decap_3 PHY_1001 ();
 sky130_fd_sc_hd__decap_3 PHY_1002 ();
 sky130_fd_sc_hd__decap_3 PHY_1003 ();
 sky130_fd_sc_hd__decap_3 PHY_1004 ();
 sky130_fd_sc_hd__decap_3 PHY_1005 ();
 sky130_fd_sc_hd__decap_3 PHY_1006 ();
 sky130_fd_sc_hd__decap_3 PHY_1007 ();
 sky130_fd_sc_hd__decap_3 PHY_1008 ();
 sky130_fd_sc_hd__decap_3 PHY_1009 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_1010 ();
 sky130_fd_sc_hd__decap_3 PHY_1011 ();
 sky130_fd_sc_hd__decap_3 PHY_1012 ();
 sky130_fd_sc_hd__decap_3 PHY_1013 ();
 sky130_fd_sc_hd__decap_3 PHY_1014 ();
 sky130_fd_sc_hd__decap_3 PHY_1015 ();
 sky130_fd_sc_hd__decap_3 PHY_1016 ();
 sky130_fd_sc_hd__decap_3 PHY_1017 ();
 sky130_fd_sc_hd__decap_3 PHY_1018 ();
 sky130_fd_sc_hd__decap_3 PHY_1019 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_1020 ();
 sky130_fd_sc_hd__decap_3 PHY_1021 ();
 sky130_fd_sc_hd__decap_3 PHY_1022 ();
 sky130_fd_sc_hd__decap_3 PHY_1023 ();
 sky130_fd_sc_hd__decap_3 PHY_1024 ();
 sky130_fd_sc_hd__decap_3 PHY_1025 ();
 sky130_fd_sc_hd__decap_3 PHY_1026 ();
 sky130_fd_sc_hd__decap_3 PHY_1027 ();
 sky130_fd_sc_hd__decap_3 PHY_1028 ();
 sky130_fd_sc_hd__decap_3 PHY_1029 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_1030 ();
 sky130_fd_sc_hd__decap_3 PHY_1031 ();
 sky130_fd_sc_hd__decap_3 PHY_1032 ();
 sky130_fd_sc_hd__decap_3 PHY_1033 ();
 sky130_fd_sc_hd__decap_3 PHY_1034 ();
 sky130_fd_sc_hd__decap_3 PHY_1035 ();
 sky130_fd_sc_hd__decap_3 PHY_1036 ();
 sky130_fd_sc_hd__decap_3 PHY_1037 ();
 sky130_fd_sc_hd__decap_3 PHY_1038 ();
 sky130_fd_sc_hd__decap_3 PHY_1039 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_1040 ();
 sky130_fd_sc_hd__decap_3 PHY_1041 ();
 sky130_fd_sc_hd__decap_3 PHY_1042 ();
 sky130_fd_sc_hd__decap_3 PHY_1043 ();
 sky130_fd_sc_hd__decap_3 PHY_1044 ();
 sky130_fd_sc_hd__decap_3 PHY_1045 ();
 sky130_fd_sc_hd__decap_3 PHY_1046 ();
 sky130_fd_sc_hd__decap_3 PHY_1047 ();
 sky130_fd_sc_hd__decap_3 PHY_1048 ();
 sky130_fd_sc_hd__decap_3 PHY_1049 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_1050 ();
 sky130_fd_sc_hd__decap_3 PHY_1051 ();
 sky130_fd_sc_hd__decap_3 PHY_1052 ();
 sky130_fd_sc_hd__decap_3 PHY_1053 ();
 sky130_fd_sc_hd__decap_3 PHY_1054 ();
 sky130_fd_sc_hd__decap_3 PHY_1055 ();
 sky130_fd_sc_hd__decap_3 PHY_1056 ();
 sky130_fd_sc_hd__decap_3 PHY_1057 ();
 sky130_fd_sc_hd__decap_3 PHY_1058 ();
 sky130_fd_sc_hd__decap_3 PHY_1059 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_1060 ();
 sky130_fd_sc_hd__decap_3 PHY_1061 ();
 sky130_fd_sc_hd__decap_3 PHY_1062 ();
 sky130_fd_sc_hd__decap_3 PHY_1063 ();
 sky130_fd_sc_hd__decap_3 PHY_1064 ();
 sky130_fd_sc_hd__decap_3 PHY_1065 ();
 sky130_fd_sc_hd__decap_3 PHY_1066 ();
 sky130_fd_sc_hd__decap_3 PHY_1067 ();
 sky130_fd_sc_hd__decap_3 PHY_1068 ();
 sky130_fd_sc_hd__decap_3 PHY_1069 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_1070 ();
 sky130_fd_sc_hd__decap_3 PHY_1071 ();
 sky130_fd_sc_hd__decap_3 PHY_1072 ();
 sky130_fd_sc_hd__decap_3 PHY_1073 ();
 sky130_fd_sc_hd__decap_3 PHY_1074 ();
 sky130_fd_sc_hd__decap_3 PHY_1075 ();
 sky130_fd_sc_hd__decap_3 PHY_1076 ();
 sky130_fd_sc_hd__decap_3 PHY_1077 ();
 sky130_fd_sc_hd__decap_3 PHY_1078 ();
 sky130_fd_sc_hd__decap_3 PHY_1079 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_1080 ();
 sky130_fd_sc_hd__decap_3 PHY_1081 ();
 sky130_fd_sc_hd__decap_3 PHY_1082 ();
 sky130_fd_sc_hd__decap_3 PHY_1083 ();
 sky130_fd_sc_hd__decap_3 PHY_1084 ();
 sky130_fd_sc_hd__decap_3 PHY_1085 ();
 sky130_fd_sc_hd__decap_3 PHY_1086 ();
 sky130_fd_sc_hd__decap_3 PHY_1087 ();
 sky130_fd_sc_hd__decap_3 PHY_1088 ();
 sky130_fd_sc_hd__decap_3 PHY_1089 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_1090 ();
 sky130_fd_sc_hd__decap_3 PHY_1091 ();
 sky130_fd_sc_hd__decap_3 PHY_1092 ();
 sky130_fd_sc_hd__decap_3 PHY_1093 ();
 sky130_fd_sc_hd__decap_3 PHY_1094 ();
 sky130_fd_sc_hd__decap_3 PHY_1095 ();
 sky130_fd_sc_hd__decap_3 PHY_1096 ();
 sky130_fd_sc_hd__decap_3 PHY_1097 ();
 sky130_fd_sc_hd__decap_3 PHY_1098 ();
 sky130_fd_sc_hd__decap_3 PHY_1099 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_1100 ();
 sky130_fd_sc_hd__decap_3 PHY_1101 ();
 sky130_fd_sc_hd__decap_3 PHY_1102 ();
 sky130_fd_sc_hd__decap_3 PHY_1103 ();
 sky130_fd_sc_hd__decap_3 PHY_1104 ();
 sky130_fd_sc_hd__decap_3 PHY_1105 ();
 sky130_fd_sc_hd__decap_3 PHY_1106 ();
 sky130_fd_sc_hd__decap_3 PHY_1107 ();
 sky130_fd_sc_hd__decap_3 PHY_1108 ();
 sky130_fd_sc_hd__decap_3 PHY_1109 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_1110 ();
 sky130_fd_sc_hd__decap_3 PHY_1111 ();
 sky130_fd_sc_hd__decap_3 PHY_1112 ();
 sky130_fd_sc_hd__decap_3 PHY_1113 ();
 sky130_fd_sc_hd__decap_3 PHY_1114 ();
 sky130_fd_sc_hd__decap_3 PHY_1115 ();
 sky130_fd_sc_hd__decap_3 PHY_1116 ();
 sky130_fd_sc_hd__decap_3 PHY_1117 ();
 sky130_fd_sc_hd__decap_3 PHY_1118 ();
 sky130_fd_sc_hd__decap_3 PHY_1119 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_1120 ();
 sky130_fd_sc_hd__decap_3 PHY_1121 ();
 sky130_fd_sc_hd__decap_3 PHY_1122 ();
 sky130_fd_sc_hd__decap_3 PHY_1123 ();
 sky130_fd_sc_hd__decap_3 PHY_1124 ();
 sky130_fd_sc_hd__decap_3 PHY_1125 ();
 sky130_fd_sc_hd__decap_3 PHY_1126 ();
 sky130_fd_sc_hd__decap_3 PHY_1127 ();
 sky130_fd_sc_hd__decap_3 PHY_1128 ();
 sky130_fd_sc_hd__decap_3 PHY_1129 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_1130 ();
 sky130_fd_sc_hd__decap_3 PHY_1131 ();
 sky130_fd_sc_hd__decap_3 PHY_1132 ();
 sky130_fd_sc_hd__decap_3 PHY_1133 ();
 sky130_fd_sc_hd__decap_3 PHY_1134 ();
 sky130_fd_sc_hd__decap_3 PHY_1135 ();
 sky130_fd_sc_hd__decap_3 PHY_1136 ();
 sky130_fd_sc_hd__decap_3 PHY_1137 ();
 sky130_fd_sc_hd__decap_3 PHY_1138 ();
 sky130_fd_sc_hd__decap_3 PHY_1139 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_1140 ();
 sky130_fd_sc_hd__decap_3 PHY_1141 ();
 sky130_fd_sc_hd__decap_3 PHY_1142 ();
 sky130_fd_sc_hd__decap_3 PHY_1143 ();
 sky130_fd_sc_hd__decap_3 PHY_1144 ();
 sky130_fd_sc_hd__decap_3 PHY_1145 ();
 sky130_fd_sc_hd__decap_3 PHY_1146 ();
 sky130_fd_sc_hd__decap_3 PHY_1147 ();
 sky130_fd_sc_hd__decap_3 PHY_1148 ();
 sky130_fd_sc_hd__decap_3 PHY_1149 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_1150 ();
 sky130_fd_sc_hd__decap_3 PHY_1151 ();
 sky130_fd_sc_hd__decap_3 PHY_1152 ();
 sky130_fd_sc_hd__decap_3 PHY_1153 ();
 sky130_fd_sc_hd__decap_3 PHY_1154 ();
 sky130_fd_sc_hd__decap_3 PHY_1155 ();
 sky130_fd_sc_hd__decap_3 PHY_1156 ();
 sky130_fd_sc_hd__decap_3 PHY_1157 ();
 sky130_fd_sc_hd__decap_3 PHY_1158 ();
 sky130_fd_sc_hd__decap_3 PHY_1159 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_1160 ();
 sky130_fd_sc_hd__decap_3 PHY_1161 ();
 sky130_fd_sc_hd__decap_3 PHY_1162 ();
 sky130_fd_sc_hd__decap_3 PHY_1163 ();
 sky130_fd_sc_hd__decap_3 PHY_1164 ();
 sky130_fd_sc_hd__decap_3 PHY_1165 ();
 sky130_fd_sc_hd__decap_3 PHY_1166 ();
 sky130_fd_sc_hd__decap_3 PHY_1167 ();
 sky130_fd_sc_hd__decap_3 PHY_1168 ();
 sky130_fd_sc_hd__decap_3 PHY_1169 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_1170 ();
 sky130_fd_sc_hd__decap_3 PHY_1171 ();
 sky130_fd_sc_hd__decap_3 PHY_1172 ();
 sky130_fd_sc_hd__decap_3 PHY_1173 ();
 sky130_fd_sc_hd__decap_3 PHY_1174 ();
 sky130_fd_sc_hd__decap_3 PHY_1175 ();
 sky130_fd_sc_hd__decap_3 PHY_1176 ();
 sky130_fd_sc_hd__decap_3 PHY_1177 ();
 sky130_fd_sc_hd__decap_3 PHY_1178 ();
 sky130_fd_sc_hd__decap_3 PHY_1179 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_1180 ();
 sky130_fd_sc_hd__decap_3 PHY_1181 ();
 sky130_fd_sc_hd__decap_3 PHY_1182 ();
 sky130_fd_sc_hd__decap_3 PHY_1183 ();
 sky130_fd_sc_hd__decap_3 PHY_1184 ();
 sky130_fd_sc_hd__decap_3 PHY_1185 ();
 sky130_fd_sc_hd__decap_3 PHY_1186 ();
 sky130_fd_sc_hd__decap_3 PHY_1187 ();
 sky130_fd_sc_hd__decap_3 PHY_1188 ();
 sky130_fd_sc_hd__decap_3 PHY_1189 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_1190 ();
 sky130_fd_sc_hd__decap_3 PHY_1191 ();
 sky130_fd_sc_hd__decap_3 PHY_1192 ();
 sky130_fd_sc_hd__decap_3 PHY_1193 ();
 sky130_fd_sc_hd__decap_3 PHY_1194 ();
 sky130_fd_sc_hd__decap_3 PHY_1195 ();
 sky130_fd_sc_hd__decap_3 PHY_1196 ();
 sky130_fd_sc_hd__decap_3 PHY_1197 ();
 sky130_fd_sc_hd__decap_3 PHY_1198 ();
 sky130_fd_sc_hd__decap_3 PHY_1199 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_1200 ();
 sky130_fd_sc_hd__decap_3 PHY_1201 ();
 sky130_fd_sc_hd__decap_3 PHY_1202 ();
 sky130_fd_sc_hd__decap_3 PHY_1203 ();
 sky130_fd_sc_hd__decap_3 PHY_1204 ();
 sky130_fd_sc_hd__decap_3 PHY_1205 ();
 sky130_fd_sc_hd__decap_3 PHY_1206 ();
 sky130_fd_sc_hd__decap_3 PHY_1207 ();
 sky130_fd_sc_hd__decap_3 PHY_1208 ();
 sky130_fd_sc_hd__decap_3 PHY_1209 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_1210 ();
 sky130_fd_sc_hd__decap_3 PHY_1211 ();
 sky130_fd_sc_hd__decap_3 PHY_1212 ();
 sky130_fd_sc_hd__decap_3 PHY_1213 ();
 sky130_fd_sc_hd__decap_3 PHY_1214 ();
 sky130_fd_sc_hd__decap_3 PHY_1215 ();
 sky130_fd_sc_hd__decap_3 PHY_1216 ();
 sky130_fd_sc_hd__decap_3 PHY_1217 ();
 sky130_fd_sc_hd__decap_3 PHY_1218 ();
 sky130_fd_sc_hd__decap_3 PHY_1219 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_1220 ();
 sky130_fd_sc_hd__decap_3 PHY_1221 ();
 sky130_fd_sc_hd__decap_3 PHY_1222 ();
 sky130_fd_sc_hd__decap_3 PHY_1223 ();
 sky130_fd_sc_hd__decap_3 PHY_1224 ();
 sky130_fd_sc_hd__decap_3 PHY_1225 ();
 sky130_fd_sc_hd__decap_3 PHY_1226 ();
 sky130_fd_sc_hd__decap_3 PHY_1227 ();
 sky130_fd_sc_hd__decap_3 PHY_1228 ();
 sky130_fd_sc_hd__decap_3 PHY_1229 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_1230 ();
 sky130_fd_sc_hd__decap_3 PHY_1231 ();
 sky130_fd_sc_hd__decap_3 PHY_1232 ();
 sky130_fd_sc_hd__decap_3 PHY_1233 ();
 sky130_fd_sc_hd__decap_3 PHY_1234 ();
 sky130_fd_sc_hd__decap_3 PHY_1235 ();
 sky130_fd_sc_hd__decap_3 PHY_1236 ();
 sky130_fd_sc_hd__decap_3 PHY_1237 ();
 sky130_fd_sc_hd__decap_3 PHY_1238 ();
 sky130_fd_sc_hd__decap_3 PHY_1239 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_1240 ();
 sky130_fd_sc_hd__decap_3 PHY_1241 ();
 sky130_fd_sc_hd__decap_3 PHY_1242 ();
 sky130_fd_sc_hd__decap_3 PHY_1243 ();
 sky130_fd_sc_hd__decap_3 PHY_1244 ();
 sky130_fd_sc_hd__decap_3 PHY_1245 ();
 sky130_fd_sc_hd__decap_3 PHY_1246 ();
 sky130_fd_sc_hd__decap_3 PHY_1247 ();
 sky130_fd_sc_hd__decap_3 PHY_1248 ();
 sky130_fd_sc_hd__decap_3 PHY_1249 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_1250 ();
 sky130_fd_sc_hd__decap_3 PHY_1251 ();
 sky130_fd_sc_hd__decap_3 PHY_1252 ();
 sky130_fd_sc_hd__decap_3 PHY_1253 ();
 sky130_fd_sc_hd__decap_3 PHY_1254 ();
 sky130_fd_sc_hd__decap_3 PHY_1255 ();
 sky130_fd_sc_hd__decap_3 PHY_1256 ();
 sky130_fd_sc_hd__decap_3 PHY_1257 ();
 sky130_fd_sc_hd__decap_3 PHY_1258 ();
 sky130_fd_sc_hd__decap_3 PHY_1259 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_1260 ();
 sky130_fd_sc_hd__decap_3 PHY_1261 ();
 sky130_fd_sc_hd__decap_3 PHY_1262 ();
 sky130_fd_sc_hd__decap_3 PHY_1263 ();
 sky130_fd_sc_hd__decap_3 PHY_1264 ();
 sky130_fd_sc_hd__decap_3 PHY_1265 ();
 sky130_fd_sc_hd__decap_3 PHY_1266 ();
 sky130_fd_sc_hd__decap_3 PHY_1267 ();
 sky130_fd_sc_hd__decap_3 PHY_1268 ();
 sky130_fd_sc_hd__decap_3 PHY_1269 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_1270 ();
 sky130_fd_sc_hd__decap_3 PHY_1271 ();
 sky130_fd_sc_hd__decap_3 PHY_1272 ();
 sky130_fd_sc_hd__decap_3 PHY_1273 ();
 sky130_fd_sc_hd__decap_3 PHY_1274 ();
 sky130_fd_sc_hd__decap_3 PHY_1275 ();
 sky130_fd_sc_hd__decap_3 PHY_1276 ();
 sky130_fd_sc_hd__decap_3 PHY_1277 ();
 sky130_fd_sc_hd__decap_3 PHY_1278 ();
 sky130_fd_sc_hd__decap_3 PHY_1279 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_1280 ();
 sky130_fd_sc_hd__decap_3 PHY_1281 ();
 sky130_fd_sc_hd__decap_3 PHY_1282 ();
 sky130_fd_sc_hd__decap_3 PHY_1283 ();
 sky130_fd_sc_hd__decap_3 PHY_1284 ();
 sky130_fd_sc_hd__decap_3 PHY_1285 ();
 sky130_fd_sc_hd__decap_3 PHY_1286 ();
 sky130_fd_sc_hd__decap_3 PHY_1287 ();
 sky130_fd_sc_hd__decap_3 PHY_1288 ();
 sky130_fd_sc_hd__decap_3 PHY_1289 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_1290 ();
 sky130_fd_sc_hd__decap_3 PHY_1291 ();
 sky130_fd_sc_hd__decap_3 PHY_1292 ();
 sky130_fd_sc_hd__decap_3 PHY_1293 ();
 sky130_fd_sc_hd__decap_3 PHY_1294 ();
 sky130_fd_sc_hd__decap_3 PHY_1295 ();
 sky130_fd_sc_hd__decap_3 PHY_1296 ();
 sky130_fd_sc_hd__decap_3 PHY_1297 ();
 sky130_fd_sc_hd__decap_3 PHY_1298 ();
 sky130_fd_sc_hd__decap_3 PHY_1299 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_1300 ();
 sky130_fd_sc_hd__decap_3 PHY_1301 ();
 sky130_fd_sc_hd__decap_3 PHY_1302 ();
 sky130_fd_sc_hd__decap_3 PHY_1303 ();
 sky130_fd_sc_hd__decap_3 PHY_1304 ();
 sky130_fd_sc_hd__decap_3 PHY_1305 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__decap_3 PHY_572 ();
 sky130_fd_sc_hd__decap_3 PHY_573 ();
 sky130_fd_sc_hd__decap_3 PHY_574 ();
 sky130_fd_sc_hd__decap_3 PHY_575 ();
 sky130_fd_sc_hd__decap_3 PHY_576 ();
 sky130_fd_sc_hd__decap_3 PHY_577 ();
 sky130_fd_sc_hd__decap_3 PHY_578 ();
 sky130_fd_sc_hd__decap_3 PHY_579 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_580 ();
 sky130_fd_sc_hd__decap_3 PHY_581 ();
 sky130_fd_sc_hd__decap_3 PHY_582 ();
 sky130_fd_sc_hd__decap_3 PHY_583 ();
 sky130_fd_sc_hd__decap_3 PHY_584 ();
 sky130_fd_sc_hd__decap_3 PHY_585 ();
 sky130_fd_sc_hd__decap_3 PHY_586 ();
 sky130_fd_sc_hd__decap_3 PHY_587 ();
 sky130_fd_sc_hd__decap_3 PHY_588 ();
 sky130_fd_sc_hd__decap_3 PHY_589 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_590 ();
 sky130_fd_sc_hd__decap_3 PHY_591 ();
 sky130_fd_sc_hd__decap_3 PHY_592 ();
 sky130_fd_sc_hd__decap_3 PHY_593 ();
 sky130_fd_sc_hd__decap_3 PHY_594 ();
 sky130_fd_sc_hd__decap_3 PHY_595 ();
 sky130_fd_sc_hd__decap_3 PHY_596 ();
 sky130_fd_sc_hd__decap_3 PHY_597 ();
 sky130_fd_sc_hd__decap_3 PHY_598 ();
 sky130_fd_sc_hd__decap_3 PHY_599 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_600 ();
 sky130_fd_sc_hd__decap_3 PHY_601 ();
 sky130_fd_sc_hd__decap_3 PHY_602 ();
 sky130_fd_sc_hd__decap_3 PHY_603 ();
 sky130_fd_sc_hd__decap_3 PHY_604 ();
 sky130_fd_sc_hd__decap_3 PHY_605 ();
 sky130_fd_sc_hd__decap_3 PHY_606 ();
 sky130_fd_sc_hd__decap_3 PHY_607 ();
 sky130_fd_sc_hd__decap_3 PHY_608 ();
 sky130_fd_sc_hd__decap_3 PHY_609 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_610 ();
 sky130_fd_sc_hd__decap_3 PHY_611 ();
 sky130_fd_sc_hd__decap_3 PHY_612 ();
 sky130_fd_sc_hd__decap_3 PHY_613 ();
 sky130_fd_sc_hd__decap_3 PHY_614 ();
 sky130_fd_sc_hd__decap_3 PHY_615 ();
 sky130_fd_sc_hd__decap_3 PHY_616 ();
 sky130_fd_sc_hd__decap_3 PHY_617 ();
 sky130_fd_sc_hd__decap_3 PHY_618 ();
 sky130_fd_sc_hd__decap_3 PHY_619 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_620 ();
 sky130_fd_sc_hd__decap_3 PHY_621 ();
 sky130_fd_sc_hd__decap_3 PHY_622 ();
 sky130_fd_sc_hd__decap_3 PHY_623 ();
 sky130_fd_sc_hd__decap_3 PHY_624 ();
 sky130_fd_sc_hd__decap_3 PHY_625 ();
 sky130_fd_sc_hd__decap_3 PHY_626 ();
 sky130_fd_sc_hd__decap_3 PHY_627 ();
 sky130_fd_sc_hd__decap_3 PHY_628 ();
 sky130_fd_sc_hd__decap_3 PHY_629 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_630 ();
 sky130_fd_sc_hd__decap_3 PHY_631 ();
 sky130_fd_sc_hd__decap_3 PHY_632 ();
 sky130_fd_sc_hd__decap_3 PHY_633 ();
 sky130_fd_sc_hd__decap_3 PHY_634 ();
 sky130_fd_sc_hd__decap_3 PHY_635 ();
 sky130_fd_sc_hd__decap_3 PHY_636 ();
 sky130_fd_sc_hd__decap_3 PHY_637 ();
 sky130_fd_sc_hd__decap_3 PHY_638 ();
 sky130_fd_sc_hd__decap_3 PHY_639 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_640 ();
 sky130_fd_sc_hd__decap_3 PHY_641 ();
 sky130_fd_sc_hd__decap_3 PHY_642 ();
 sky130_fd_sc_hd__decap_3 PHY_643 ();
 sky130_fd_sc_hd__decap_3 PHY_644 ();
 sky130_fd_sc_hd__decap_3 PHY_645 ();
 sky130_fd_sc_hd__decap_3 PHY_646 ();
 sky130_fd_sc_hd__decap_3 PHY_647 ();
 sky130_fd_sc_hd__decap_3 PHY_648 ();
 sky130_fd_sc_hd__decap_3 PHY_649 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_650 ();
 sky130_fd_sc_hd__decap_3 PHY_651 ();
 sky130_fd_sc_hd__decap_3 PHY_652 ();
 sky130_fd_sc_hd__decap_3 PHY_653 ();
 sky130_fd_sc_hd__decap_3 PHY_654 ();
 sky130_fd_sc_hd__decap_3 PHY_655 ();
 sky130_fd_sc_hd__decap_3 PHY_656 ();
 sky130_fd_sc_hd__decap_3 PHY_657 ();
 sky130_fd_sc_hd__decap_3 PHY_658 ();
 sky130_fd_sc_hd__decap_3 PHY_659 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_660 ();
 sky130_fd_sc_hd__decap_3 PHY_661 ();
 sky130_fd_sc_hd__decap_3 PHY_662 ();
 sky130_fd_sc_hd__decap_3 PHY_663 ();
 sky130_fd_sc_hd__decap_3 PHY_664 ();
 sky130_fd_sc_hd__decap_3 PHY_665 ();
 sky130_fd_sc_hd__decap_3 PHY_666 ();
 sky130_fd_sc_hd__decap_3 PHY_667 ();
 sky130_fd_sc_hd__decap_3 PHY_668 ();
 sky130_fd_sc_hd__decap_3 PHY_669 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_670 ();
 sky130_fd_sc_hd__decap_3 PHY_671 ();
 sky130_fd_sc_hd__decap_3 PHY_672 ();
 sky130_fd_sc_hd__decap_3 PHY_673 ();
 sky130_fd_sc_hd__decap_3 PHY_674 ();
 sky130_fd_sc_hd__decap_3 PHY_675 ();
 sky130_fd_sc_hd__decap_3 PHY_676 ();
 sky130_fd_sc_hd__decap_3 PHY_677 ();
 sky130_fd_sc_hd__decap_3 PHY_678 ();
 sky130_fd_sc_hd__decap_3 PHY_679 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_680 ();
 sky130_fd_sc_hd__decap_3 PHY_681 ();
 sky130_fd_sc_hd__decap_3 PHY_682 ();
 sky130_fd_sc_hd__decap_3 PHY_683 ();
 sky130_fd_sc_hd__decap_3 PHY_684 ();
 sky130_fd_sc_hd__decap_3 PHY_685 ();
 sky130_fd_sc_hd__decap_3 PHY_686 ();
 sky130_fd_sc_hd__decap_3 PHY_687 ();
 sky130_fd_sc_hd__decap_3 PHY_688 ();
 sky130_fd_sc_hd__decap_3 PHY_689 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_690 ();
 sky130_fd_sc_hd__decap_3 PHY_691 ();
 sky130_fd_sc_hd__decap_3 PHY_692 ();
 sky130_fd_sc_hd__decap_3 PHY_693 ();
 sky130_fd_sc_hd__decap_3 PHY_694 ();
 sky130_fd_sc_hd__decap_3 PHY_695 ();
 sky130_fd_sc_hd__decap_3 PHY_696 ();
 sky130_fd_sc_hd__decap_3 PHY_697 ();
 sky130_fd_sc_hd__decap_3 PHY_698 ();
 sky130_fd_sc_hd__decap_3 PHY_699 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_700 ();
 sky130_fd_sc_hd__decap_3 PHY_701 ();
 sky130_fd_sc_hd__decap_3 PHY_702 ();
 sky130_fd_sc_hd__decap_3 PHY_703 ();
 sky130_fd_sc_hd__decap_3 PHY_704 ();
 sky130_fd_sc_hd__decap_3 PHY_705 ();
 sky130_fd_sc_hd__decap_3 PHY_706 ();
 sky130_fd_sc_hd__decap_3 PHY_707 ();
 sky130_fd_sc_hd__decap_3 PHY_708 ();
 sky130_fd_sc_hd__decap_3 PHY_709 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_710 ();
 sky130_fd_sc_hd__decap_3 PHY_711 ();
 sky130_fd_sc_hd__decap_3 PHY_712 ();
 sky130_fd_sc_hd__decap_3 PHY_713 ();
 sky130_fd_sc_hd__decap_3 PHY_714 ();
 sky130_fd_sc_hd__decap_3 PHY_715 ();
 sky130_fd_sc_hd__decap_3 PHY_716 ();
 sky130_fd_sc_hd__decap_3 PHY_717 ();
 sky130_fd_sc_hd__decap_3 PHY_718 ();
 sky130_fd_sc_hd__decap_3 PHY_719 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_720 ();
 sky130_fd_sc_hd__decap_3 PHY_721 ();
 sky130_fd_sc_hd__decap_3 PHY_722 ();
 sky130_fd_sc_hd__decap_3 PHY_723 ();
 sky130_fd_sc_hd__decap_3 PHY_724 ();
 sky130_fd_sc_hd__decap_3 PHY_725 ();
 sky130_fd_sc_hd__decap_3 PHY_726 ();
 sky130_fd_sc_hd__decap_3 PHY_727 ();
 sky130_fd_sc_hd__decap_3 PHY_728 ();
 sky130_fd_sc_hd__decap_3 PHY_729 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_730 ();
 sky130_fd_sc_hd__decap_3 PHY_731 ();
 sky130_fd_sc_hd__decap_3 PHY_732 ();
 sky130_fd_sc_hd__decap_3 PHY_733 ();
 sky130_fd_sc_hd__decap_3 PHY_734 ();
 sky130_fd_sc_hd__decap_3 PHY_735 ();
 sky130_fd_sc_hd__decap_3 PHY_736 ();
 sky130_fd_sc_hd__decap_3 PHY_737 ();
 sky130_fd_sc_hd__decap_3 PHY_738 ();
 sky130_fd_sc_hd__decap_3 PHY_739 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_740 ();
 sky130_fd_sc_hd__decap_3 PHY_741 ();
 sky130_fd_sc_hd__decap_3 PHY_742 ();
 sky130_fd_sc_hd__decap_3 PHY_743 ();
 sky130_fd_sc_hd__decap_3 PHY_744 ();
 sky130_fd_sc_hd__decap_3 PHY_745 ();
 sky130_fd_sc_hd__decap_3 PHY_746 ();
 sky130_fd_sc_hd__decap_3 PHY_747 ();
 sky130_fd_sc_hd__decap_3 PHY_748 ();
 sky130_fd_sc_hd__decap_3 PHY_749 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_750 ();
 sky130_fd_sc_hd__decap_3 PHY_751 ();
 sky130_fd_sc_hd__decap_3 PHY_752 ();
 sky130_fd_sc_hd__decap_3 PHY_753 ();
 sky130_fd_sc_hd__decap_3 PHY_754 ();
 sky130_fd_sc_hd__decap_3 PHY_755 ();
 sky130_fd_sc_hd__decap_3 PHY_756 ();
 sky130_fd_sc_hd__decap_3 PHY_757 ();
 sky130_fd_sc_hd__decap_3 PHY_758 ();
 sky130_fd_sc_hd__decap_3 PHY_759 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_760 ();
 sky130_fd_sc_hd__decap_3 PHY_761 ();
 sky130_fd_sc_hd__decap_3 PHY_762 ();
 sky130_fd_sc_hd__decap_3 PHY_763 ();
 sky130_fd_sc_hd__decap_3 PHY_764 ();
 sky130_fd_sc_hd__decap_3 PHY_765 ();
 sky130_fd_sc_hd__decap_3 PHY_766 ();
 sky130_fd_sc_hd__decap_3 PHY_767 ();
 sky130_fd_sc_hd__decap_3 PHY_768 ();
 sky130_fd_sc_hd__decap_3 PHY_769 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_770 ();
 sky130_fd_sc_hd__decap_3 PHY_771 ();
 sky130_fd_sc_hd__decap_3 PHY_772 ();
 sky130_fd_sc_hd__decap_3 PHY_773 ();
 sky130_fd_sc_hd__decap_3 PHY_774 ();
 sky130_fd_sc_hd__decap_3 PHY_775 ();
 sky130_fd_sc_hd__decap_3 PHY_776 ();
 sky130_fd_sc_hd__decap_3 PHY_777 ();
 sky130_fd_sc_hd__decap_3 PHY_778 ();
 sky130_fd_sc_hd__decap_3 PHY_779 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_780 ();
 sky130_fd_sc_hd__decap_3 PHY_781 ();
 sky130_fd_sc_hd__decap_3 PHY_782 ();
 sky130_fd_sc_hd__decap_3 PHY_783 ();
 sky130_fd_sc_hd__decap_3 PHY_784 ();
 sky130_fd_sc_hd__decap_3 PHY_785 ();
 sky130_fd_sc_hd__decap_3 PHY_786 ();
 sky130_fd_sc_hd__decap_3 PHY_787 ();
 sky130_fd_sc_hd__decap_3 PHY_788 ();
 sky130_fd_sc_hd__decap_3 PHY_789 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_790 ();
 sky130_fd_sc_hd__decap_3 PHY_791 ();
 sky130_fd_sc_hd__decap_3 PHY_792 ();
 sky130_fd_sc_hd__decap_3 PHY_793 ();
 sky130_fd_sc_hd__decap_3 PHY_794 ();
 sky130_fd_sc_hd__decap_3 PHY_795 ();
 sky130_fd_sc_hd__decap_3 PHY_796 ();
 sky130_fd_sc_hd__decap_3 PHY_797 ();
 sky130_fd_sc_hd__decap_3 PHY_798 ();
 sky130_fd_sc_hd__decap_3 PHY_799 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_800 ();
 sky130_fd_sc_hd__decap_3 PHY_801 ();
 sky130_fd_sc_hd__decap_3 PHY_802 ();
 sky130_fd_sc_hd__decap_3 PHY_803 ();
 sky130_fd_sc_hd__decap_3 PHY_804 ();
 sky130_fd_sc_hd__decap_3 PHY_805 ();
 sky130_fd_sc_hd__decap_3 PHY_806 ();
 sky130_fd_sc_hd__decap_3 PHY_807 ();
 sky130_fd_sc_hd__decap_3 PHY_808 ();
 sky130_fd_sc_hd__decap_3 PHY_809 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_810 ();
 sky130_fd_sc_hd__decap_3 PHY_811 ();
 sky130_fd_sc_hd__decap_3 PHY_812 ();
 sky130_fd_sc_hd__decap_3 PHY_813 ();
 sky130_fd_sc_hd__decap_3 PHY_814 ();
 sky130_fd_sc_hd__decap_3 PHY_815 ();
 sky130_fd_sc_hd__decap_3 PHY_816 ();
 sky130_fd_sc_hd__decap_3 PHY_817 ();
 sky130_fd_sc_hd__decap_3 PHY_818 ();
 sky130_fd_sc_hd__decap_3 PHY_819 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_820 ();
 sky130_fd_sc_hd__decap_3 PHY_821 ();
 sky130_fd_sc_hd__decap_3 PHY_822 ();
 sky130_fd_sc_hd__decap_3 PHY_823 ();
 sky130_fd_sc_hd__decap_3 PHY_824 ();
 sky130_fd_sc_hd__decap_3 PHY_825 ();
 sky130_fd_sc_hd__decap_3 PHY_826 ();
 sky130_fd_sc_hd__decap_3 PHY_827 ();
 sky130_fd_sc_hd__decap_3 PHY_828 ();
 sky130_fd_sc_hd__decap_3 PHY_829 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_830 ();
 sky130_fd_sc_hd__decap_3 PHY_831 ();
 sky130_fd_sc_hd__decap_3 PHY_832 ();
 sky130_fd_sc_hd__decap_3 PHY_833 ();
 sky130_fd_sc_hd__decap_3 PHY_834 ();
 sky130_fd_sc_hd__decap_3 PHY_835 ();
 sky130_fd_sc_hd__decap_3 PHY_836 ();
 sky130_fd_sc_hd__decap_3 PHY_837 ();
 sky130_fd_sc_hd__decap_3 PHY_838 ();
 sky130_fd_sc_hd__decap_3 PHY_839 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_840 ();
 sky130_fd_sc_hd__decap_3 PHY_841 ();
 sky130_fd_sc_hd__decap_3 PHY_842 ();
 sky130_fd_sc_hd__decap_3 PHY_843 ();
 sky130_fd_sc_hd__decap_3 PHY_844 ();
 sky130_fd_sc_hd__decap_3 PHY_845 ();
 sky130_fd_sc_hd__decap_3 PHY_846 ();
 sky130_fd_sc_hd__decap_3 PHY_847 ();
 sky130_fd_sc_hd__decap_3 PHY_848 ();
 sky130_fd_sc_hd__decap_3 PHY_849 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_850 ();
 sky130_fd_sc_hd__decap_3 PHY_851 ();
 sky130_fd_sc_hd__decap_3 PHY_852 ();
 sky130_fd_sc_hd__decap_3 PHY_853 ();
 sky130_fd_sc_hd__decap_3 PHY_854 ();
 sky130_fd_sc_hd__decap_3 PHY_855 ();
 sky130_fd_sc_hd__decap_3 PHY_856 ();
 sky130_fd_sc_hd__decap_3 PHY_857 ();
 sky130_fd_sc_hd__decap_3 PHY_858 ();
 sky130_fd_sc_hd__decap_3 PHY_859 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_860 ();
 sky130_fd_sc_hd__decap_3 PHY_861 ();
 sky130_fd_sc_hd__decap_3 PHY_862 ();
 sky130_fd_sc_hd__decap_3 PHY_863 ();
 sky130_fd_sc_hd__decap_3 PHY_864 ();
 sky130_fd_sc_hd__decap_3 PHY_865 ();
 sky130_fd_sc_hd__decap_3 PHY_866 ();
 sky130_fd_sc_hd__decap_3 PHY_867 ();
 sky130_fd_sc_hd__decap_3 PHY_868 ();
 sky130_fd_sc_hd__decap_3 PHY_869 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_870 ();
 sky130_fd_sc_hd__decap_3 PHY_871 ();
 sky130_fd_sc_hd__decap_3 PHY_872 ();
 sky130_fd_sc_hd__decap_3 PHY_873 ();
 sky130_fd_sc_hd__decap_3 PHY_874 ();
 sky130_fd_sc_hd__decap_3 PHY_875 ();
 sky130_fd_sc_hd__decap_3 PHY_876 ();
 sky130_fd_sc_hd__decap_3 PHY_877 ();
 sky130_fd_sc_hd__decap_3 PHY_878 ();
 sky130_fd_sc_hd__decap_3 PHY_879 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_880 ();
 sky130_fd_sc_hd__decap_3 PHY_881 ();
 sky130_fd_sc_hd__decap_3 PHY_882 ();
 sky130_fd_sc_hd__decap_3 PHY_883 ();
 sky130_fd_sc_hd__decap_3 PHY_884 ();
 sky130_fd_sc_hd__decap_3 PHY_885 ();
 sky130_fd_sc_hd__decap_3 PHY_886 ();
 sky130_fd_sc_hd__decap_3 PHY_887 ();
 sky130_fd_sc_hd__decap_3 PHY_888 ();
 sky130_fd_sc_hd__decap_3 PHY_889 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_890 ();
 sky130_fd_sc_hd__decap_3 PHY_891 ();
 sky130_fd_sc_hd__decap_3 PHY_892 ();
 sky130_fd_sc_hd__decap_3 PHY_893 ();
 sky130_fd_sc_hd__decap_3 PHY_894 ();
 sky130_fd_sc_hd__decap_3 PHY_895 ();
 sky130_fd_sc_hd__decap_3 PHY_896 ();
 sky130_fd_sc_hd__decap_3 PHY_897 ();
 sky130_fd_sc_hd__decap_3 PHY_898 ();
 sky130_fd_sc_hd__decap_3 PHY_899 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_900 ();
 sky130_fd_sc_hd__decap_3 PHY_901 ();
 sky130_fd_sc_hd__decap_3 PHY_902 ();
 sky130_fd_sc_hd__decap_3 PHY_903 ();
 sky130_fd_sc_hd__decap_3 PHY_904 ();
 sky130_fd_sc_hd__decap_3 PHY_905 ();
 sky130_fd_sc_hd__decap_3 PHY_906 ();
 sky130_fd_sc_hd__decap_3 PHY_907 ();
 sky130_fd_sc_hd__decap_3 PHY_908 ();
 sky130_fd_sc_hd__decap_3 PHY_909 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_910 ();
 sky130_fd_sc_hd__decap_3 PHY_911 ();
 sky130_fd_sc_hd__decap_3 PHY_912 ();
 sky130_fd_sc_hd__decap_3 PHY_913 ();
 sky130_fd_sc_hd__decap_3 PHY_914 ();
 sky130_fd_sc_hd__decap_3 PHY_915 ();
 sky130_fd_sc_hd__decap_3 PHY_916 ();
 sky130_fd_sc_hd__decap_3 PHY_917 ();
 sky130_fd_sc_hd__decap_3 PHY_918 ();
 sky130_fd_sc_hd__decap_3 PHY_919 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_920 ();
 sky130_fd_sc_hd__decap_3 PHY_921 ();
 sky130_fd_sc_hd__decap_3 PHY_922 ();
 sky130_fd_sc_hd__decap_3 PHY_923 ();
 sky130_fd_sc_hd__decap_3 PHY_924 ();
 sky130_fd_sc_hd__decap_3 PHY_925 ();
 sky130_fd_sc_hd__decap_3 PHY_926 ();
 sky130_fd_sc_hd__decap_3 PHY_927 ();
 sky130_fd_sc_hd__decap_3 PHY_928 ();
 sky130_fd_sc_hd__decap_3 PHY_929 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_930 ();
 sky130_fd_sc_hd__decap_3 PHY_931 ();
 sky130_fd_sc_hd__decap_3 PHY_932 ();
 sky130_fd_sc_hd__decap_3 PHY_933 ();
 sky130_fd_sc_hd__decap_3 PHY_934 ();
 sky130_fd_sc_hd__decap_3 PHY_935 ();
 sky130_fd_sc_hd__decap_3 PHY_936 ();
 sky130_fd_sc_hd__decap_3 PHY_937 ();
 sky130_fd_sc_hd__decap_3 PHY_938 ();
 sky130_fd_sc_hd__decap_3 PHY_939 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_940 ();
 sky130_fd_sc_hd__decap_3 PHY_941 ();
 sky130_fd_sc_hd__decap_3 PHY_942 ();
 sky130_fd_sc_hd__decap_3 PHY_943 ();
 sky130_fd_sc_hd__decap_3 PHY_944 ();
 sky130_fd_sc_hd__decap_3 PHY_945 ();
 sky130_fd_sc_hd__decap_3 PHY_946 ();
 sky130_fd_sc_hd__decap_3 PHY_947 ();
 sky130_fd_sc_hd__decap_3 PHY_948 ();
 sky130_fd_sc_hd__decap_3 PHY_949 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_950 ();
 sky130_fd_sc_hd__decap_3 PHY_951 ();
 sky130_fd_sc_hd__decap_3 PHY_952 ();
 sky130_fd_sc_hd__decap_3 PHY_953 ();
 sky130_fd_sc_hd__decap_3 PHY_954 ();
 sky130_fd_sc_hd__decap_3 PHY_955 ();
 sky130_fd_sc_hd__decap_3 PHY_956 ();
 sky130_fd_sc_hd__decap_3 PHY_957 ();
 sky130_fd_sc_hd__decap_3 PHY_958 ();
 sky130_fd_sc_hd__decap_3 PHY_959 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_960 ();
 sky130_fd_sc_hd__decap_3 PHY_961 ();
 sky130_fd_sc_hd__decap_3 PHY_962 ();
 sky130_fd_sc_hd__decap_3 PHY_963 ();
 sky130_fd_sc_hd__decap_3 PHY_964 ();
 sky130_fd_sc_hd__decap_3 PHY_965 ();
 sky130_fd_sc_hd__decap_3 PHY_966 ();
 sky130_fd_sc_hd__decap_3 PHY_967 ();
 sky130_fd_sc_hd__decap_3 PHY_968 ();
 sky130_fd_sc_hd__decap_3 PHY_969 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_970 ();
 sky130_fd_sc_hd__decap_3 PHY_971 ();
 sky130_fd_sc_hd__decap_3 PHY_972 ();
 sky130_fd_sc_hd__decap_3 PHY_973 ();
 sky130_fd_sc_hd__decap_3 PHY_974 ();
 sky130_fd_sc_hd__decap_3 PHY_975 ();
 sky130_fd_sc_hd__decap_3 PHY_976 ();
 sky130_fd_sc_hd__decap_3 PHY_977 ();
 sky130_fd_sc_hd__decap_3 PHY_978 ();
 sky130_fd_sc_hd__decap_3 PHY_979 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_980 ();
 sky130_fd_sc_hd__decap_3 PHY_981 ();
 sky130_fd_sc_hd__decap_3 PHY_982 ();
 sky130_fd_sc_hd__decap_3 PHY_983 ();
 sky130_fd_sc_hd__decap_3 PHY_984 ();
 sky130_fd_sc_hd__decap_3 PHY_985 ();
 sky130_fd_sc_hd__decap_3 PHY_986 ();
 sky130_fd_sc_hd__decap_3 PHY_987 ();
 sky130_fd_sc_hd__decap_3 PHY_988 ();
 sky130_fd_sc_hd__decap_3 PHY_989 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_990 ();
 sky130_fd_sc_hd__decap_3 PHY_991 ();
 sky130_fd_sc_hd__decap_3 PHY_992 ();
 sky130_fd_sc_hd__decap_3 PHY_993 ();
 sky130_fd_sc_hd__decap_3 PHY_994 ();
 sky130_fd_sc_hd__decap_3 PHY_995 ();
 sky130_fd_sc_hd__decap_3 PHY_996 ();
 sky130_fd_sc_hd__decap_3 PHY_997 ();
 sky130_fd_sc_hd__decap_3 PHY_998 ();
 sky130_fd_sc_hd__decap_3 PHY_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8510 ();
 sky130_fd_sc_hd__inv_2 _3612_ (.A(net1369),
    .Y(_1669_));
 sky130_fd_sc_hd__inv_2 _3613_ (.A(net1372),
    .Y(_1670_));
 sky130_fd_sc_hd__inv_2 _3614_ (.A(m2_wbd_bl_i[0]),
    .Y(_1671_));
 sky130_fd_sc_hd__inv_2 _3615_ (.A(net1404),
    .Y(_1672_));
 sky130_fd_sc_hd__clkinv_4 _3616_ (.A(net1405),
    .Y(_1673_));
 sky130_fd_sc_hd__clkinv_2 _3617_ (.A(net1874),
    .Y(_1674_));
 sky130_fd_sc_hd__inv_2 _3618_ (.A(\u_s1.u_sync_wbb.u_resp_if.wr_ptr[0] ),
    .Y(_1675_));
 sky130_fd_sc_hd__inv_2 _3619_ (.A(net1409),
    .Y(_1676_));
 sky130_fd_sc_hd__inv_2 _3620_ (.A(net1408),
    .Y(_1677_));
 sky130_fd_sc_hd__inv_2 _3621_ (.A(m2_wbd_bry_i),
    .Y(_1678_));
 sky130_fd_sc_hd__inv_2 _3622_ (.A(\u_s2.u_sync_wbb.m_bl_cnt[0] ),
    .Y(_1679_));
 sky130_fd_sc_hd__inv_2 _3623_ (.A(net1817),
    .Y(_1680_));
 sky130_fd_sc_hd__inv_2 _3624_ (.A(net1798),
    .Y(_1681_));
 sky130_fd_sc_hd__inv_2 _3625_ (.A(net1396),
    .Y(_1682_));
 sky130_fd_sc_hd__inv_2 _3626_ (.A(net1900),
    .Y(_1683_));
 sky130_fd_sc_hd__clkinv_2 _3627_ (.A(m0_wbd_adr_i[17]),
    .Y(_1684_));
 sky130_fd_sc_hd__clkinv_2 _3628_ (.A(m0_wbd_adr_i[16]),
    .Y(_1685_));
 sky130_fd_sc_hd__inv_2 _3629_ (.A(m0_wbd_stb_i),
    .Y(_1686_));
 sky130_fd_sc_hd__inv_2 _3630_ (.A(m3_wbd_stb_i),
    .Y(_1687_));
 sky130_fd_sc_hd__inv_2 _3631_ (.A(m2_wbd_stb_i),
    .Y(_1688_));
 sky130_fd_sc_hd__inv_2 _3632_ (.A(m1_wbd_adr_i[17]),
    .Y(_1689_));
 sky130_fd_sc_hd__clkinv_4 _3633_ (.A(m1_wbd_stb_i),
    .Y(_1690_));
 sky130_fd_sc_hd__inv_2 _3634_ (.A(net1826),
    .Y(_1691_));
 sky130_fd_sc_hd__inv_2 _3635_ (.A(\u_s1.u_sync_wbb.m_state[1] ),
    .Y(_1692_));
 sky130_fd_sc_hd__inv_2 _3636_ (.A(\u_s1.u_sync_wbb.m_cmd_wr_en ),
    .Y(_1693_));
 sky130_fd_sc_hd__clkinv_4 _3637_ (.A(\u_s1.u_sync_wbb.wbm_lack_o ),
    .Y(_1694_));
 sky130_fd_sc_hd__inv_2 _3638_ (.A(net1925),
    .Y(_1695_));
 sky130_fd_sc_hd__inv_2 _3639_ (.A(\u_s0.u_sync_wbb.wbs_ack_f ),
    .Y(_1696_));
 sky130_fd_sc_hd__inv_2 _3640_ (.A(\u_dcg_s0.hcnt[0] ),
    .Y(_1697_));
 sky130_fd_sc_hd__inv_2 _3641_ (.A(\u_dcg_s0.hcnt[3] ),
    .Y(_1698_));
 sky130_fd_sc_hd__inv_2 _3642_ (.A(\u_s0.u_sync_wbb.m_bl_cnt[0] ),
    .Y(_1699_));
 sky130_fd_sc_hd__clkinv_2 _3643_ (.A(\u_s0.u_sync_wbb.m_state[0] ),
    .Y(_1700_));
 sky130_fd_sc_hd__inv_2 _3644_ (.A(\u_s0.u_sync_wbb.m_state[2] ),
    .Y(_1701_));
 sky130_fd_sc_hd__inv_2 _3645_ (.A(\u_s1.u_sync_wbb.wbs_ack_f ),
    .Y(_1702_));
 sky130_fd_sc_hd__inv_2 _3646_ (.A(\u_s1.u_sync_wbb.wbs_stb_l ),
    .Y(_1703_));
 sky130_fd_sc_hd__inv_2 _3647_ (.A(net1508),
    .Y(_1704_));
 sky130_fd_sc_hd__inv_2 _3648_ (.A(\u_s0.u_sync_wbb.wbs_stb_l ),
    .Y(_1705_));
 sky130_fd_sc_hd__inv_2 _3649_ (.A(s0_wbd_lack_i),
    .Y(_1706_));
 sky130_fd_sc_hd__inv_2 _3650_ (.A(net1276),
    .Y(_1707_));
 sky130_fd_sc_hd__inv_2 _3651_ (.A(net1274),
    .Y(_1708_));
 sky130_fd_sc_hd__inv_2 _3652_ (.A(\u_s2.u_sync_wbb.wbs_ack_f ),
    .Y(_1709_));
 sky130_fd_sc_hd__inv_2 _3653_ (.A(\u_s2.u_sync_wbb.wbs_stb_l ),
    .Y(_1710_));
 sky130_fd_sc_hd__inv_2 _3654_ (.A(net1499),
    .Y(_1711_));
 sky130_fd_sc_hd__nand2b_1 _3655_ (.A_N(net1328),
    .B(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .Y(_1712_));
 sky130_fd_sc_hd__xor2_2 _3656_ (.A(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .B(net1328),
    .X(_1713_));
 sky130_fd_sc_hd__and2b_1 _3657_ (.A_N(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .B(net1338),
    .X(_1714_));
 sky130_fd_sc_hd__xor2_1 _3658_ (.A(net1338),
    .B(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .X(_1715_));
 sky130_fd_sc_hd__nor2_1 _3659_ (.A(_1713_),
    .B(_1715_),
    .Y(_1716_));
 sky130_fd_sc_hd__xor2_2 _3660_ (.A(\u_s0.u_sync_wbb.u_cmd_if.rd_ptr[2] ),
    .B(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[2] ),
    .X(_1717_));
 sky130_fd_sc_hd__or3_1 _3661_ (.A(_1713_),
    .B(_1715_),
    .C(_1717_),
    .X(_1718_));
 sky130_fd_sc_hd__a21oi_2 _3662_ (.A1(_1696_),
    .A2(net827),
    .B1(\u_s0.u_sync_wbb.wbs_burst ),
    .Y(_1719_));
 sky130_fd_sc_hd__clkinv_2 _3663_ (.A(_1719_),
    .Y(net342));
 sky130_fd_sc_hd__o21a_1 _3664_ (.A1(_1713_),
    .A2(_1714_),
    .B1(_1712_),
    .X(_1720_));
 sky130_fd_sc_hd__xnor2_1 _3665_ (.A(_1717_),
    .B(_1720_),
    .Y(_1721_));
 sky130_fd_sc_hd__xor2_1 _3666_ (.A(_1713_),
    .B(_1714_),
    .X(_1722_));
 sky130_fd_sc_hd__and3_1 _3667_ (.A(\u_s0.u_sync_wbb.m_cmd_wr_en ),
    .B(_1715_),
    .C(_1722_),
    .X(_1723_));
 sky130_fd_sc_hd__nor2_2 _3668_ (.A(net1368),
    .B(net1254),
    .Y(_1724_));
 sky130_fd_sc_hd__nand2_1 _3669_ (.A(net1264),
    .B(net1372),
    .Y(_1725_));
 sky130_fd_sc_hd__and3b_1 _3670_ (.A_N(net1371),
    .B(net1375),
    .C(net1563),
    .X(_1726_));
 sky130_fd_sc_hd__and2_1 _3671_ (.A(net1369),
    .B(net1373),
    .X(_1727_));
 sky130_fd_sc_hd__and3_1 _3672_ (.A(net1371),
    .B(net1375),
    .C(m3_wbd_bry_i),
    .X(_1728_));
 sky130_fd_sc_hd__nor2_4 _3673_ (.A(net1368),
    .B(net1372),
    .Y(_1729_));
 sky130_fd_sc_hd__or2_2 _3674_ (.A(net1371),
    .B(net1375),
    .X(_1730_));
 sky130_fd_sc_hd__and2b_1 _3675_ (.A_N(\u_s0.gnt[0] ),
    .B(net1371),
    .X(_1731_));
 sky130_fd_sc_hd__inv_2 _3676_ (.A(net1193),
    .Y(_1732_));
 sky130_fd_sc_hd__a2111o_2 _3677_ (.A1(net1259),
    .A2(m2_wbd_bry_i),
    .B1(_1726_),
    .C1(_1728_),
    .D1(net1205),
    .X(_1733_));
 sky130_fd_sc_hd__a21bo_1 _3678_ (.A1(_1716_),
    .A2(_1717_),
    .B1_N(_1733_),
    .X(_1734_));
 sky130_fd_sc_hd__a21o_2 _3679_ (.A1(_1721_),
    .A2(_1723_),
    .B1(_1734_),
    .X(_1735_));
 sky130_fd_sc_hd__or4_1 _3680_ (.A(m3_wbd_adr_i[21]),
    .B(m3_wbd_adr_i[20]),
    .C(m3_wbd_adr_i[23]),
    .D(m3_wbd_adr_i[22]),
    .X(_1736_));
 sky130_fd_sc_hd__or4b_2 _3681_ (.A(m3_wbd_adr_i[29]),
    .B(m3_wbd_adr_i[31]),
    .C(m3_wbd_adr_i[30]),
    .D_N(m3_wbd_adr_i[28]),
    .X(_1737_));
 sky130_fd_sc_hd__or4_1 _3682_ (.A(m3_wbd_adr_i[25]),
    .B(m3_wbd_adr_i[24]),
    .C(m3_wbd_adr_i[27]),
    .D(m3_wbd_adr_i[26]),
    .X(_1738_));
 sky130_fd_sc_hd__or2_1 _3683_ (.A(m3_wbd_adr_i[19]),
    .B(m3_wbd_adr_i[18]),
    .X(_1739_));
 sky130_fd_sc_hd__or3b_1 _3684_ (.A(m3_wbd_adr_i[19]),
    .B(m3_wbd_adr_i[18]),
    .C_N(m3_wbd_adr_i[16]),
    .X(_1740_));
 sky130_fd_sc_hd__or4_4 _3685_ (.A(_1736_),
    .B(_1737_),
    .C(_1738_),
    .D(_1740_),
    .X(_1741_));
 sky130_fd_sc_hd__or3b_1 _3686_ (.A(m3_wbd_adr_i[19]),
    .B(m3_wbd_adr_i[18]),
    .C_N(m3_wbd_adr_i[17]),
    .X(_1742_));
 sky130_fd_sc_hd__or4_4 _3687_ (.A(_1736_),
    .B(_1737_),
    .C(_1738_),
    .D(_1742_),
    .X(_1743_));
 sky130_fd_sc_hd__or4_1 _3688_ (.A(_1736_),
    .B(_1737_),
    .C(_1738_),
    .D(_1740_),
    .X(_1744_));
 sky130_fd_sc_hd__or4_1 _3689_ (.A(_1736_),
    .B(_1737_),
    .C(_1738_),
    .D(_1742_),
    .X(_1745_));
 sky130_fd_sc_hd__or4_1 _3690_ (.A(_1736_),
    .B(_1737_),
    .C(_1738_),
    .D(_1739_),
    .X(_1746_));
 sky130_fd_sc_hd__and3_4 _3691_ (.A(net1208),
    .B(_1741_),
    .C(_1743_),
    .X(_1747_));
 sky130_fd_sc_hd__or2_1 _3692_ (.A(m0_wbd_adr_i[25]),
    .B(m0_wbd_adr_i[24]),
    .X(_1748_));
 sky130_fd_sc_hd__or4b_4 _3693_ (.A(m0_wbd_adr_i[27]),
    .B(m0_wbd_adr_i[26]),
    .C(m0_wbd_adr_i[29]),
    .D_N(m0_wbd_adr_i[28]),
    .X(_1749_));
 sky130_fd_sc_hd__or4_4 _3694_ (.A(m0_wbd_adr_i[31]),
    .B(m0_wbd_adr_i[30]),
    .C(m0_wbd_adr_i[21]),
    .D(m0_wbd_adr_i[20]),
    .X(_1750_));
 sky130_fd_sc_hd__or4_4 _3695_ (.A(m0_wbd_adr_i[23]),
    .B(m0_wbd_adr_i[22]),
    .C(m0_wbd_adr_i[19]),
    .D(m0_wbd_adr_i[18]),
    .X(_1751_));
 sky130_fd_sc_hd__or4_4 _3696_ (.A(_1748_),
    .B(_1749_),
    .C(_1750_),
    .D(_1751_),
    .X(_1752_));
 sky130_fd_sc_hd__nor3_1 _3697_ (.A(_1748_),
    .B(_1749_),
    .C(_1750_),
    .Y(_1753_));
 sky130_fd_sc_hd__or4_4 _3698_ (.A(_1748_),
    .B(_1749_),
    .C(_1750_),
    .D(_1751_),
    .X(_1754_));
 sky130_fd_sc_hd__nor2_1 _3699_ (.A(_1684_),
    .B(_1751_),
    .Y(_1755_));
 sky130_fd_sc_hd__a2bb2oi_4 _3700_ (.A1_N(_1685_),
    .A2_N(_1754_),
    .B1(_1755_),
    .B2(_1753_),
    .Y(_1756_));
 sky130_fd_sc_hd__and2_4 _3701_ (.A(net1203),
    .B(_1756_),
    .X(_1757_));
 sky130_fd_sc_hd__and2_1 _3702_ (.A(m0_wbd_stb_i),
    .B(_1756_),
    .X(_1758_));
 sky130_fd_sc_hd__a32oi_4 _3703_ (.A1(m0_wbd_stb_i),
    .A2(net1203),
    .A3(_1756_),
    .B1(_1747_),
    .B2(m3_wbd_stb_i),
    .Y(_1759_));
 sky130_fd_sc_hd__or3b_1 _3704_ (.A(m1_wbd_adr_i[21]),
    .B(m1_wbd_adr_i[20]),
    .C_N(m1_wbd_adr_i[16]),
    .X(_1760_));
 sky130_fd_sc_hd__or4b_4 _3705_ (.A(m1_wbd_adr_i[29]),
    .B(m1_wbd_adr_i[31]),
    .C(m1_wbd_adr_i[30]),
    .D_N(m1_wbd_adr_i[28]),
    .X(_1761_));
 sky130_fd_sc_hd__or4_1 _3706_ (.A(m1_wbd_adr_i[25]),
    .B(m1_wbd_adr_i[24]),
    .C(m1_wbd_adr_i[27]),
    .D(m1_wbd_adr_i[26]),
    .X(_1762_));
 sky130_fd_sc_hd__or4_1 _3707_ (.A(m1_wbd_adr_i[23]),
    .B(m1_wbd_adr_i[22]),
    .C(m1_wbd_adr_i[19]),
    .D(m1_wbd_adr_i[18]),
    .X(_1763_));
 sky130_fd_sc_hd__or4_4 _3708_ (.A(_1760_),
    .B(_1761_),
    .C(_1762_),
    .D(_1763_),
    .X(_1764_));
 sky130_fd_sc_hd__or3b_1 _3709_ (.A(m1_wbd_adr_i[21]),
    .B(m1_wbd_adr_i[20]),
    .C_N(m1_wbd_adr_i[17]),
    .X(_1765_));
 sky130_fd_sc_hd__or4_4 _3710_ (.A(_1761_),
    .B(_1762_),
    .C(_1763_),
    .D(_1765_),
    .X(_1766_));
 sky130_fd_sc_hd__or4_4 _3711_ (.A(_1760_),
    .B(_1761_),
    .C(_1762_),
    .D(_1763_),
    .X(_1767_));
 sky130_fd_sc_hd__or4_4 _3712_ (.A(_1761_),
    .B(_1762_),
    .C(_1763_),
    .D(_1765_),
    .X(_1768_));
 sky130_fd_sc_hd__and3_4 _3713_ (.A(net821),
    .B(_1767_),
    .C(_1768_),
    .X(_1769_));
 sky130_fd_sc_hd__or4_4 _3714_ (.A(m2_wbd_adr_i[21]),
    .B(m2_wbd_adr_i[20]),
    .C(m2_wbd_adr_i[23]),
    .D(m2_wbd_adr_i[22]),
    .X(_1770_));
 sky130_fd_sc_hd__or4b_4 _3715_ (.A(m2_wbd_adr_i[29]),
    .B(m2_wbd_adr_i[31]),
    .C(m2_wbd_adr_i[30]),
    .D_N(m2_wbd_adr_i[28]),
    .X(_1771_));
 sky130_fd_sc_hd__or4_1 _3716_ (.A(m2_wbd_adr_i[25]),
    .B(m2_wbd_adr_i[24]),
    .C(m2_wbd_adr_i[27]),
    .D(m2_wbd_adr_i[26]),
    .X(_1772_));
 sky130_fd_sc_hd__or2_1 _3717_ (.A(m2_wbd_adr_i[19]),
    .B(m2_wbd_adr_i[18]),
    .X(_1773_));
 sky130_fd_sc_hd__or3b_1 _3718_ (.A(m2_wbd_adr_i[19]),
    .B(m2_wbd_adr_i[18]),
    .C_N(m2_wbd_adr_i[16]),
    .X(_1774_));
 sky130_fd_sc_hd__or4_4 _3719_ (.A(_1770_),
    .B(_1771_),
    .C(_1772_),
    .D(_1774_),
    .X(_1775_));
 sky130_fd_sc_hd__or3b_1 _3720_ (.A(m2_wbd_adr_i[19]),
    .B(m2_wbd_adr_i[18]),
    .C_N(m2_wbd_adr_i[17]),
    .X(_1776_));
 sky130_fd_sc_hd__or4_4 _3721_ (.A(_1770_),
    .B(_1771_),
    .C(_1772_),
    .D(_1776_),
    .X(_1777_));
 sky130_fd_sc_hd__or4_1 _3722_ (.A(_1770_),
    .B(_1771_),
    .C(_1772_),
    .D(_1774_),
    .X(_1778_));
 sky130_fd_sc_hd__or4_1 _3723_ (.A(_1770_),
    .B(_1771_),
    .C(_1772_),
    .D(_1773_),
    .X(_1779_));
 sky130_fd_sc_hd__and3_4 _3724_ (.A(net1193),
    .B(_1775_),
    .C(_1777_),
    .X(_1780_));
 sky130_fd_sc_hd__and3_1 _3725_ (.A(m2_wbd_stb_i),
    .B(_1775_),
    .C(_1777_),
    .X(_1781_));
 sky130_fd_sc_hd__a22oi_4 _3726_ (.A1(m1_wbd_stb_i),
    .A2(net736),
    .B1(net810),
    .B2(m2_wbd_stb_i),
    .Y(_1782_));
 sky130_fd_sc_hd__a21o_1 _3727_ (.A1(_1759_),
    .A2(_1782_),
    .B1(\u_s0.u_sync_wbb.wbm_lack_o ),
    .X(_1783_));
 sky130_fd_sc_hd__a211o_2 _3728_ (.A1(_1759_),
    .A2(_1782_),
    .B1(\u_s0.u_sync_wbb.wbm_lack_o ),
    .C1(_1735_),
    .X(_1784_));
 sky130_fd_sc_hd__a221o_1 _3729_ (.A1(net1262),
    .A2(m2_wbd_bl_i[0]),
    .B1(net1207),
    .B2(m3_wbd_bl_i[0]),
    .C1(_1729_),
    .X(_1785_));
 sky130_fd_sc_hd__a21o_2 _3730_ (.A1(net1564),
    .A2(net823),
    .B1(_1785_),
    .X(_1786_));
 sky130_fd_sc_hd__a22o_4 _3731_ (.A1(m3_wbd_bl_i[9]),
    .A2(net1207),
    .B1(net1193),
    .B2(m2_wbd_bl_i[9]),
    .X(_1787_));
 sky130_fd_sc_hd__a22o_1 _3732_ (.A1(m3_wbd_bl_i[1]),
    .A2(net1207),
    .B1(net1193),
    .B2(m2_wbd_bl_i[1]),
    .X(_1788_));
 sky130_fd_sc_hd__a21o_4 _3733_ (.A1(m1_wbd_bl_i[1]),
    .A2(net823),
    .B1(_1788_),
    .X(_1789_));
 sky130_fd_sc_hd__or3b_1 _3734_ (.A(_1787_),
    .B(_1789_),
    .C_N(_1786_),
    .X(_1790_));
 sky130_fd_sc_hd__a22o_1 _3735_ (.A1(m3_wbd_bl_i[2]),
    .A2(net1207),
    .B1(net1193),
    .B2(m2_wbd_bl_i[2]),
    .X(_1791_));
 sky130_fd_sc_hd__a21o_2 _3736_ (.A1(m1_wbd_bl_i[2]),
    .A2(net823),
    .B1(_1791_),
    .X(_1792_));
 sky130_fd_sc_hd__a22o_2 _3737_ (.A1(m3_wbd_bl_i[4]),
    .A2(net1207),
    .B1(net1193),
    .B2(m2_wbd_bl_i[4]),
    .X(_1793_));
 sky130_fd_sc_hd__a22o_2 _3738_ (.A1(m3_wbd_bl_i[3]),
    .A2(net1207),
    .B1(net1193),
    .B2(m2_wbd_bl_i[3]),
    .X(_1794_));
 sky130_fd_sc_hd__or2_1 _3739_ (.A(_1792_),
    .B(_1794_),
    .X(_1795_));
 sky130_fd_sc_hd__a22o_2 _3740_ (.A1(m3_wbd_bl_i[7]),
    .A2(net1207),
    .B1(net1193),
    .B2(m2_wbd_bl_i[7]),
    .X(_1796_));
 sky130_fd_sc_hd__a22o_2 _3741_ (.A1(m3_wbd_bl_i[6]),
    .A2(net1207),
    .B1(net1193),
    .B2(m2_wbd_bl_i[6]),
    .X(_1797_));
 sky130_fd_sc_hd__or2_1 _3742_ (.A(_1796_),
    .B(_1797_),
    .X(_1798_));
 sky130_fd_sc_hd__a22o_2 _3743_ (.A1(m3_wbd_bl_i[8]),
    .A2(net1207),
    .B1(net1193),
    .B2(m2_wbd_bl_i[8]),
    .X(_1799_));
 sky130_fd_sc_hd__a22o_1 _3744_ (.A1(m3_wbd_bl_i[5]),
    .A2(net1209),
    .B1(_1731_),
    .B2(m2_wbd_bl_i[5]),
    .X(_1800_));
 sky130_fd_sc_hd__nor3_1 _3745_ (.A(_1798_),
    .B(_1799_),
    .C(net808),
    .Y(_1801_));
 sky130_fd_sc_hd__inv_2 _3746_ (.A(_1801_),
    .Y(_1802_));
 sky130_fd_sc_hd__nor4_2 _3747_ (.A(_1790_),
    .B(_1793_),
    .C(_1795_),
    .D(_1802_),
    .Y(_1803_));
 sky130_fd_sc_hd__and3_1 _3748_ (.A(net1271),
    .B(net1375),
    .C(m1_wbd_we_i),
    .X(_1804_));
 sky130_fd_sc_hd__a221o_1 _3749_ (.A1(net1259),
    .A2(m2_wbd_we_i),
    .B1(net1208),
    .B2(m3_wbd_we_i),
    .C1(net1204),
    .X(_1805_));
 sky130_fd_sc_hd__o22a_4 _3750_ (.A1(m0_wbd_we_i),
    .A2(net1199),
    .B1(_1804_),
    .B2(_1805_),
    .X(_1806_));
 sky130_fd_sc_hd__inv_2 _3751_ (.A(_1806_),
    .Y(_1807_));
 sky130_fd_sc_hd__and3b_1 _3752_ (.A_N(\u_s0.u_sync_wbb.wbm_lack_o ),
    .B(\u_s0.u_sync_wbb.m_state[0] ),
    .C(_1733_),
    .X(_1808_));
 sky130_fd_sc_hd__and3_1 _3753_ (.A(_1803_),
    .B(_1806_),
    .C(_1808_),
    .X(_1809_));
 sky130_fd_sc_hd__and2b_1 _3754_ (.A_N(net1315),
    .B(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .X(_1810_));
 sky130_fd_sc_hd__nand2b_1 _3755_ (.A_N(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[0] ),
    .B(net1320),
    .Y(_1811_));
 sky130_fd_sc_hd__xnor2_2 _3756_ (.A(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .B(net1315),
    .Y(_1812_));
 sky130_fd_sc_hd__a21o_1 _3757_ (.A1(_1811_),
    .A2(_1812_),
    .B1(_1810_),
    .X(_1813_));
 sky130_fd_sc_hd__xor2_4 _3758_ (.A(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[2] ),
    .B(\u_s0.u_sync_wbb.u_resp_if.rd_ptr[2] ),
    .X(_1814_));
 sky130_fd_sc_hd__xnor2_4 _3759_ (.A(_1813_),
    .B(_1814_),
    .Y(_1815_));
 sky130_fd_sc_hd__xnor2_1 _3760_ (.A(_1811_),
    .B(_1812_),
    .Y(_1816_));
 sky130_fd_sc_hd__xnor2_1 _3761_ (.A(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[0] ),
    .B(net1321),
    .Y(_1817_));
 sky130_fd_sc_hd__xor2_1 _3762_ (.A(\u_s0.u_sync_wbb.wbm_ack_o ),
    .B(_1817_),
    .X(_1818_));
 sky130_fd_sc_hd__nand2_1 _3763_ (.A(_1816_),
    .B(_1818_),
    .Y(_1819_));
 sky130_fd_sc_hd__o21ai_1 _3764_ (.A1(_1815_),
    .A2(_1819_),
    .B1(_1733_),
    .Y(_1820_));
 sky130_fd_sc_hd__o211a_1 _3765_ (.A1(_1815_),
    .A2(_1819_),
    .B1(\u_s0.u_sync_wbb.m_state[1] ),
    .C1(_1733_),
    .X(_1821_));
 sky130_fd_sc_hd__nor2_1 _3766_ (.A(_1701_),
    .B(_1735_),
    .Y(_1822_));
 sky130_fd_sc_hd__or2_1 _3767_ (.A(_1821_),
    .B(_1822_),
    .X(_1823_));
 sky130_fd_sc_hd__or4_4 _3768_ (.A(\u_s0.u_sync_wbb.m_bl_cnt[7] ),
    .B(\u_s0.u_sync_wbb.m_bl_cnt[6] ),
    .C(\u_s0.u_sync_wbb.m_bl_cnt[9] ),
    .D(\u_s0.u_sync_wbb.m_bl_cnt[8] ),
    .X(_1824_));
 sky130_fd_sc_hd__or4_1 _3769_ (.A(_1699_),
    .B(\u_s0.u_sync_wbb.m_bl_cnt[1] ),
    .C(\u_s0.u_sync_wbb.m_bl_cnt[5] ),
    .D(\u_s0.u_sync_wbb.m_bl_cnt[4] ),
    .X(_1825_));
 sky130_fd_sc_hd__nor4_1 _3770_ (.A(\u_s0.u_sync_wbb.m_bl_cnt[3] ),
    .B(\u_s0.u_sync_wbb.m_bl_cnt[2] ),
    .C(_1824_),
    .D(_1825_),
    .Y(_1826_));
 sky130_fd_sc_hd__or4_1 _3771_ (.A(\u_s0.u_sync_wbb.m_bl_cnt[3] ),
    .B(\u_s0.u_sync_wbb.m_bl_cnt[2] ),
    .C(_1824_),
    .D(_1825_),
    .X(_1827_));
 sky130_fd_sc_hd__or4_1 _3772_ (.A(_1699_),
    .B(\u_s0.u_sync_wbb.m_bl_cnt[1] ),
    .C(\u_s0.u_sync_wbb.m_bl_cnt[3] ),
    .D(\u_s0.u_sync_wbb.m_bl_cnt[4] ),
    .X(_1828_));
 sky130_fd_sc_hd__nor4_1 _3773_ (.A(\u_s0.u_sync_wbb.m_bl_cnt[2] ),
    .B(\u_s0.u_sync_wbb.m_bl_cnt[5] ),
    .C(_1824_),
    .D(_1828_),
    .Y(_1829_));
 sky130_fd_sc_hd__a221o_1 _3774_ (.A1(\u_s0.u_sync_wbb.m_state[0] ),
    .A2(_1784_),
    .B1(_1823_),
    .B2(_1826_),
    .C1(_1809_),
    .X(_0000_));
 sky130_fd_sc_hd__nor2_4 _3775_ (.A(net1404),
    .B(net1405),
    .Y(_1830_));
 sky130_fd_sc_hd__or2_4 _3776_ (.A(net1404),
    .B(net1405),
    .X(_1831_));
 sky130_fd_sc_hd__and2_2 _3777_ (.A(net1404),
    .B(net1405),
    .X(_1832_));
 sky130_fd_sc_hd__and2b_4 _3778_ (.A_N(\u_s1.gnt[1] ),
    .B(net1406),
    .X(_1833_));
 sky130_fd_sc_hd__nand2_2 _3779_ (.A(net1245),
    .B(net1405),
    .Y(_1834_));
 sky130_fd_sc_hd__and2_1 _3780_ (.A(m1_wbd_we_i),
    .B(net1183),
    .X(_1835_));
 sky130_fd_sc_hd__a221o_1 _3781_ (.A1(net1240),
    .A2(m2_wbd_we_i),
    .B1(net1185),
    .B2(m3_wbd_we_i),
    .C1(net1192),
    .X(_1836_));
 sky130_fd_sc_hd__o22a_1 _3782_ (.A1(m0_wbd_we_i),
    .A2(net1187),
    .B1(_1835_),
    .B2(_1836_),
    .X(_1837_));
 sky130_fd_sc_hd__and2b_1 _3783_ (.A_N(net1358),
    .B(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .X(_1838_));
 sky130_fd_sc_hd__xor2_1 _3784_ (.A(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[2] ),
    .B(\u_s1.u_sync_wbb.u_cmd_if.rd_ptr[2] ),
    .X(_1839_));
 sky130_fd_sc_hd__xnor2_1 _3785_ (.A(_1838_),
    .B(_1839_),
    .Y(_1840_));
 sky130_fd_sc_hd__and2b_1 _3786_ (.A_N(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .B(net1365),
    .X(_1841_));
 sky130_fd_sc_hd__xnor2_1 _3787_ (.A(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .B(net1357),
    .Y(_1842_));
 sky130_fd_sc_hd__and2b_1 _3788_ (.A_N(_1841_),
    .B(_1842_),
    .X(_1843_));
 sky130_fd_sc_hd__and2b_1 _3789_ (.A_N(net1365),
    .B(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .X(_1844_));
 sky130_fd_sc_hd__nor2_1 _3790_ (.A(_1842_),
    .B(_1844_),
    .Y(_1845_));
 sky130_fd_sc_hd__a21oi_1 _3791_ (.A1(net1404),
    .A2(_1678_),
    .B1(net1406),
    .Y(_1846_));
 sky130_fd_sc_hd__a221o_1 _3792_ (.A1(net1252),
    .A2(net1563),
    .B1(net1186),
    .B2(m3_wbd_bry_i),
    .C1(_1846_),
    .X(_1847_));
 sky130_fd_sc_hd__or4bb_1 _3793_ (.A(_1841_),
    .B(_1844_),
    .C_N(_1842_),
    .D_N(_1839_),
    .X(_1848_));
 sky130_fd_sc_hd__o41a_2 _3794_ (.A1(_1693_),
    .A2(_1840_),
    .A3(_1843_),
    .A4(_1845_),
    .B1(_1848_),
    .X(_1849_));
 sky130_fd_sc_hd__nand2_1 _3795_ (.A(net807),
    .B(_1849_),
    .Y(_1850_));
 sky130_fd_sc_hd__and2b_4 _3796_ (.A_N(net1405),
    .B(net1404),
    .X(_1851_));
 sky130_fd_sc_hd__nor3b_2 _3797_ (.A(m2_wbd_adr_i[17]),
    .B(_1775_),
    .C_N(net1182),
    .Y(_1852_));
 sky130_fd_sc_hd__nor2_2 _3798_ (.A(m3_wbd_adr_i[17]),
    .B(_1741_),
    .Y(_1853_));
 sky130_fd_sc_hd__or4b_1 _3799_ (.A(m3_wbd_adr_i[17]),
    .B(_1687_),
    .C(_1741_),
    .D_N(net1185),
    .X(_1854_));
 sky130_fd_sc_hd__and4b_2 _3800_ (.A_N(_1752_),
    .B(_1684_),
    .C(m0_wbd_adr_i[16]),
    .D(_1830_),
    .X(_1855_));
 sky130_fd_sc_hd__a22o_4 _3801_ (.A1(m3_wbd_bl_i[4]),
    .A2(net1186),
    .B1(net1182),
    .B2(m2_wbd_bl_i[4]),
    .X(_1856_));
 sky130_fd_sc_hd__and3_1 _3802_ (.A(net1404),
    .B(net1406),
    .C(m3_wbd_bl_i[2]),
    .X(_1857_));
 sky130_fd_sc_hd__a221o_1 _3803_ (.A1(m1_wbd_bl_i[2]),
    .A2(net1183),
    .B1(net1182),
    .B2(m2_wbd_bl_i[2]),
    .C1(_1857_),
    .X(_1858_));
 sky130_fd_sc_hd__inv_2 _3804_ (.A(net798),
    .Y(_1859_));
 sky130_fd_sc_hd__a22o_4 _3805_ (.A1(m3_wbd_bl_i[3]),
    .A2(net1186),
    .B1(net1182),
    .B2(m2_wbd_bl_i[3]),
    .X(_1860_));
 sky130_fd_sc_hd__inv_2 _3806_ (.A(_1860_),
    .Y(_1861_));
 sky130_fd_sc_hd__and3_1 _3807_ (.A(net1404),
    .B(net1405),
    .C(m3_wbd_bl_i[1]),
    .X(_1862_));
 sky130_fd_sc_hd__a221o_1 _3808_ (.A1(m1_wbd_bl_i[1]),
    .A2(net1184),
    .B1(net1182),
    .B2(m2_wbd_bl_i[1]),
    .C1(_1862_),
    .X(_1863_));
 sky130_fd_sc_hd__inv_2 _3809_ (.A(net797),
    .Y(_1864_));
 sky130_fd_sc_hd__or4_1 _3810_ (.A(_1856_),
    .B(net798),
    .C(_1860_),
    .D(net797),
    .X(_1865_));
 sky130_fd_sc_hd__a22o_4 _3811_ (.A1(m3_wbd_bl_i[8]),
    .A2(net1186),
    .B1(net1182),
    .B2(m2_wbd_bl_i[8]),
    .X(_1866_));
 sky130_fd_sc_hd__a22o_2 _3812_ (.A1(m3_wbd_bl_i[7]),
    .A2(net1186),
    .B1(net1182),
    .B2(m2_wbd_bl_i[7]),
    .X(_1867_));
 sky130_fd_sc_hd__a22o_4 _3813_ (.A1(m3_wbd_bl_i[6]),
    .A2(net1186),
    .B1(net1182),
    .B2(m2_wbd_bl_i[6]),
    .X(_1868_));
 sky130_fd_sc_hd__a22o_4 _3814_ (.A1(m3_wbd_bl_i[5]),
    .A2(net1186),
    .B1(_1851_),
    .B2(m2_wbd_bl_i[5]),
    .X(_1869_));
 sky130_fd_sc_hd__or3_1 _3815_ (.A(_1867_),
    .B(_1868_),
    .C(_1869_),
    .X(_1870_));
 sky130_fd_sc_hd__nor2_1 _3816_ (.A(_1866_),
    .B(_1870_),
    .Y(_1871_));
 sky130_fd_sc_hd__or2_1 _3817_ (.A(_1866_),
    .B(_1870_),
    .X(_1872_));
 sky130_fd_sc_hd__a22o_4 _3818_ (.A1(m3_wbd_bl_i[9]),
    .A2(_1832_),
    .B1(_1851_),
    .B2(m2_wbd_bl_i[9]),
    .X(_1873_));
 sky130_fd_sc_hd__a21oi_1 _3819_ (.A1(_1671_),
    .A2(\u_s1.gnt[1] ),
    .B1(net1406),
    .Y(_1874_));
 sky130_fd_sc_hd__a221o_4 _3820_ (.A1(net1564),
    .A2(net1252),
    .B1(_1832_),
    .B2(m3_wbd_bl_i[0]),
    .C1(_1874_),
    .X(_1875_));
 sky130_fd_sc_hd__or4b_1 _3821_ (.A(_1865_),
    .B(_1872_),
    .C(_1873_),
    .D_N(_1875_),
    .X(_1876_));
 sky130_fd_sc_hd__and3_1 _3822_ (.A(_1694_),
    .B(net807),
    .C(_1849_),
    .X(_1877_));
 sky130_fd_sc_hd__or4_4 _3823_ (.A(m0_wbd_adr_i[17]),
    .B(_1685_),
    .C(_1686_),
    .D(_1754_),
    .X(_1878_));
 sky130_fd_sc_hd__and2b_2 _3824_ (.A_N(_1767_),
    .B(_1765_),
    .X(_1879_));
 sky130_fd_sc_hd__or4b_4 _3825_ (.A(_1690_),
    .B(_1767_),
    .C(_1834_),
    .D_N(_1765_),
    .X(_1880_));
 sky130_fd_sc_hd__or4b_1 _3826_ (.A(m2_wbd_adr_i[17]),
    .B(_1688_),
    .C(_1775_),
    .D_N(net1182),
    .X(_1881_));
 sky130_fd_sc_hd__o2111ai_2 _3827_ (.A1(net1187),
    .A2(_1878_),
    .B1(_1880_),
    .C1(_1881_),
    .D1(_1854_),
    .Y(_1882_));
 sky130_fd_sc_hd__and2_1 _3828_ (.A(_1877_),
    .B(net630),
    .X(_1883_));
 sky130_fd_sc_hd__and2b_1 _3829_ (.A_N(\u_s1.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .B(net1345),
    .X(_1884_));
 sky130_fd_sc_hd__xnor2_2 _3830_ (.A(\u_s1.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .B(net1344),
    .Y(_1885_));
 sky130_fd_sc_hd__a22oi_4 _3831_ (.A1(_1675_),
    .A2(net1348),
    .B1(\u_s1.u_sync_wbb.wbm_ack_o ),
    .B2(_1885_),
    .Y(_1886_));
 sky130_fd_sc_hd__o21ai_2 _3832_ (.A1(_1675_),
    .A2(net1348),
    .B1(_1885_),
    .Y(_1887_));
 sky130_fd_sc_hd__a21oi_4 _3833_ (.A1(\u_s1.u_sync_wbb.wbm_ack_o ),
    .A2(_1887_),
    .B1(_1886_),
    .Y(_1888_));
 sky130_fd_sc_hd__xnor2_1 _3834_ (.A(\u_s1.u_sync_wbb.u_resp_if.wr_ptr[2] ),
    .B(\u_s1.u_sync_wbb.u_resp_if.rd_ptr[2] ),
    .Y(_1889_));
 sky130_fd_sc_hd__xnor2_1 _3835_ (.A(_1884_),
    .B(_1889_),
    .Y(_1890_));
 sky130_fd_sc_hd__a21o_1 _3836_ (.A1(_1886_),
    .A2(_1887_),
    .B1(_1890_),
    .X(_1891_));
 sky130_fd_sc_hd__o21ai_4 _3837_ (.A1(_1888_),
    .A2(_1891_),
    .B1(net807),
    .Y(_1892_));
 sky130_fd_sc_hd__nor2_1 _3838_ (.A(_1692_),
    .B(_1892_),
    .Y(_1893_));
 sky130_fd_sc_hd__and3_1 _3839_ (.A(\u_s1.u_sync_wbb.m_state[2] ),
    .B(net807),
    .C(_1849_),
    .X(_1894_));
 sky130_fd_sc_hd__or2_2 _3840_ (.A(_1893_),
    .B(_1894_),
    .X(_1895_));
 sky130_fd_sc_hd__or4_4 _3841_ (.A(\u_s1.u_sync_wbb.m_bl_cnt[7] ),
    .B(\u_s1.u_sync_wbb.m_bl_cnt[6] ),
    .C(\u_s1.u_sync_wbb.m_bl_cnt[9] ),
    .D(\u_s1.u_sync_wbb.m_bl_cnt[8] ),
    .X(_1896_));
 sky130_fd_sc_hd__or4b_1 _3842_ (.A(\u_s1.u_sync_wbb.m_bl_cnt[1] ),
    .B(\u_s1.u_sync_wbb.m_bl_cnt[5] ),
    .C(\u_s1.u_sync_wbb.m_bl_cnt[4] ),
    .D_N(\u_s1.u_sync_wbb.m_bl_cnt[0] ),
    .X(_1897_));
 sky130_fd_sc_hd__or4_2 _3843_ (.A(net1962),
    .B(\u_s1.u_sync_wbb.m_bl_cnt[2] ),
    .C(_1896_),
    .D(_1897_),
    .X(_1898_));
 sky130_fd_sc_hd__nand2_1 _3844_ (.A(\u_s1.u_sync_wbb.m_state[0] ),
    .B(net732),
    .Y(_1899_));
 sky130_fd_sc_hd__nor2_1 _3845_ (.A(_1876_),
    .B(_1899_),
    .Y(_1900_));
 sky130_fd_sc_hd__or4b_1 _3846_ (.A(\u_s1.u_sync_wbb.m_bl_cnt[1] ),
    .B(\u_s1.u_sync_wbb.m_bl_cnt[3] ),
    .C(\u_s1.u_sync_wbb.m_bl_cnt[4] ),
    .D_N(\u_s1.u_sync_wbb.m_bl_cnt[0] ),
    .X(_1901_));
 sky130_fd_sc_hd__nor4_2 _3847_ (.A(\u_s1.u_sync_wbb.m_bl_cnt[2] ),
    .B(\u_s1.u_sync_wbb.m_bl_cnt[5] ),
    .C(_1896_),
    .D(_1901_),
    .Y(_1902_));
 sky130_fd_sc_hd__a21oi_2 _3848_ (.A1(_1877_),
    .A2(net630),
    .B1(_1695_),
    .Y(_1903_));
 sky130_fd_sc_hd__a211o_1 _3849_ (.A1(_1895_),
    .A2(_1902_),
    .B1(_1903_),
    .C1(_1900_),
    .X(_0003_));
 sky130_fd_sc_hd__mux4_2 _3850_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][9] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][9] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][9] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][9] ),
    .S0(net1339),
    .S1(net1329),
    .X(_1904_));
 sky130_fd_sc_hd__mux2_4 _3851_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[9] ),
    .A1(_1904_),
    .S(net832),
    .X(net340));
 sky130_fd_sc_hd__mux4_2 _3852_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][8] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][8] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][8] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][8] ),
    .S0(net1341),
    .S1(net1331),
    .X(_1905_));
 sky130_fd_sc_hd__mux2_1 _3853_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[8] ),
    .A1(_1905_),
    .S(net831),
    .X(net339));
 sky130_fd_sc_hd__mux4_2 _3854_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][7] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][7] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][7] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][7] ),
    .S0(net1341),
    .S1(net1331),
    .X(_1906_));
 sky130_fd_sc_hd__mux2_1 _3855_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[7] ),
    .A1(_1906_),
    .S(net831),
    .X(net338));
 sky130_fd_sc_hd__mux4_2 _3856_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][6] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][6] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][6] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][6] ),
    .S0(net1340),
    .S1(net1330),
    .X(_1907_));
 sky130_fd_sc_hd__mux2_1 _3857_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[6] ),
    .A1(_1907_),
    .S(net831),
    .X(net337));
 sky130_fd_sc_hd__mux4_2 _3858_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][5] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][5] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][5] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][5] ),
    .S0(net1340),
    .S1(net1330),
    .X(_1908_));
 sky130_fd_sc_hd__mux2_1 _3859_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[5] ),
    .A1(_1908_),
    .S(net832),
    .X(net336));
 sky130_fd_sc_hd__mux4_2 _3860_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][4] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][4] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][4] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][4] ),
    .S0(net1340),
    .S1(net1330),
    .X(_1909_));
 sky130_fd_sc_hd__mux2_2 _3861_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[4] ),
    .A1(_1909_),
    .S(net830),
    .X(net335));
 sky130_fd_sc_hd__mux4_2 _3862_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][3] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][3] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][3] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][3] ),
    .S0(net1341),
    .S1(net1331),
    .X(_1910_));
 sky130_fd_sc_hd__mux2_1 _3863_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[3] ),
    .A1(_1910_),
    .S(net831),
    .X(net334));
 sky130_fd_sc_hd__mux4_1 _3864_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][2] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][2] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][2] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][2] ),
    .S0(net1340),
    .S1(net1330),
    .X(_1911_));
 sky130_fd_sc_hd__mux2_1 _3865_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[2] ),
    .A1(net1181),
    .S(net827),
    .X(net333));
 sky130_fd_sc_hd__mux4_2 _3866_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][1] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][1] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][1] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][1] ),
    .S0(net1334),
    .S1(net1324),
    .X(_1912_));
 sky130_fd_sc_hd__mux2_1 _3867_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[1] ),
    .A1(_1912_),
    .S(net827),
    .X(net332));
 sky130_fd_sc_hd__or2_1 _3868_ (.A(_1700_),
    .B(_1784_),
    .X(_1913_));
 sky130_fd_sc_hd__o21ai_1 _3869_ (.A1(_1735_),
    .A2(_1827_),
    .B1(\u_s0.u_sync_wbb.m_state[2] ),
    .Y(_1914_));
 sky130_fd_sc_hd__o31ai_1 _3870_ (.A1(_1803_),
    .A2(_1807_),
    .A3(_1913_),
    .B1(_1914_),
    .Y(_0002_));
 sky130_fd_sc_hd__and2b_1 _3871_ (.A_N(net1410),
    .B(net1408),
    .X(_1915_));
 sky130_fd_sc_hd__nand2_2 _3872_ (.A(net1232),
    .B(net1407),
    .Y(_1916_));
 sky130_fd_sc_hd__and2_1 _3873_ (.A(net1410),
    .B(\u_s2.gnt[1] ),
    .X(_1917_));
 sky130_fd_sc_hd__a22o_1 _3874_ (.A1(m2_wbd_bl_i[4]),
    .A2(net1180),
    .B1(net1177),
    .B2(m3_wbd_bl_i[4]),
    .X(_1918_));
 sky130_fd_sc_hd__and3_1 _3875_ (.A(m3_wbd_bl_i[2]),
    .B(net1410),
    .C(net1408),
    .X(_1919_));
 sky130_fd_sc_hd__and2b_1 _3876_ (.A_N(net1407),
    .B(net1409),
    .X(_1920_));
 sky130_fd_sc_hd__a221o_2 _3877_ (.A1(m2_wbd_bl_i[2]),
    .A2(net1180),
    .B1(net1174),
    .B2(m1_wbd_bl_i[2]),
    .C1(_1919_),
    .X(_1921_));
 sky130_fd_sc_hd__a22o_1 _3878_ (.A1(m2_wbd_bl_i[3]),
    .A2(net1180),
    .B1(net1177),
    .B2(m3_wbd_bl_i[3]),
    .X(_1922_));
 sky130_fd_sc_hd__and3_1 _3879_ (.A(m3_wbd_bl_i[1]),
    .B(net1410),
    .C(net1408),
    .X(_1923_));
 sky130_fd_sc_hd__a221o_2 _3880_ (.A1(m2_wbd_bl_i[1]),
    .A2(net1180),
    .B1(net1174),
    .B2(m1_wbd_bl_i[1]),
    .C1(_1923_),
    .X(_1924_));
 sky130_fd_sc_hd__or4_2 _3881_ (.A(net796),
    .B(net794),
    .C(net793),
    .D(net791),
    .X(_1925_));
 sky130_fd_sc_hd__a22o_1 _3882_ (.A1(m2_wbd_bl_i[8]),
    .A2(net1180),
    .B1(net1177),
    .B2(m3_wbd_bl_i[8]),
    .X(_1926_));
 sky130_fd_sc_hd__a22o_2 _3883_ (.A1(m2_wbd_bl_i[7]),
    .A2(net1180),
    .B1(net1177),
    .B2(m3_wbd_bl_i[7]),
    .X(_1927_));
 sky130_fd_sc_hd__inv_2 _3884_ (.A(net789),
    .Y(_1928_));
 sky130_fd_sc_hd__a22o_2 _3885_ (.A1(m2_wbd_bl_i[6]),
    .A2(net1180),
    .B1(net1177),
    .B2(m3_wbd_bl_i[6]),
    .X(_1929_));
 sky130_fd_sc_hd__inv_2 _3886_ (.A(net788),
    .Y(_1930_));
 sky130_fd_sc_hd__a22oi_4 _3887_ (.A1(m2_wbd_bl_i[5]),
    .A2(net1180),
    .B1(net1177),
    .B2(m3_wbd_bl_i[5]),
    .Y(_1931_));
 sky130_fd_sc_hd__a22o_1 _3888_ (.A1(m2_wbd_bl_i[5]),
    .A2(net1180),
    .B1(net1178),
    .B2(m3_wbd_bl_i[5]),
    .X(_1932_));
 sky130_fd_sc_hd__or3_1 _3889_ (.A(net789),
    .B(net788),
    .C(net786),
    .X(_1933_));
 sky130_fd_sc_hd__a22o_2 _3890_ (.A1(m2_wbd_bl_i[9]),
    .A2(_1915_),
    .B1(net1177),
    .B2(m3_wbd_bl_i[9]),
    .X(_1934_));
 sky130_fd_sc_hd__nor2_1 _3891_ (.A(net1409),
    .B(net1407),
    .Y(_1935_));
 sky130_fd_sc_hd__or2_1 _3892_ (.A(net1409),
    .B(net1407),
    .X(_1936_));
 sky130_fd_sc_hd__a21oi_2 _3893_ (.A1(_1671_),
    .A2(\u_s2.gnt[1] ),
    .B1(\u_s2.gnt[0] ),
    .Y(_1937_));
 sky130_fd_sc_hd__a221oi_4 _3894_ (.A1(net1564),
    .A2(net1225),
    .B1(net1177),
    .B2(m3_wbd_bl_i[0]),
    .C1(_1937_),
    .Y(_1938_));
 sky130_fd_sc_hd__a221o_2 _3895_ (.A1(net1564),
    .A2(net1225),
    .B1(net1177),
    .B2(m3_wbd_bl_i[0]),
    .C1(_1937_),
    .X(_1939_));
 sky130_fd_sc_hd__or3_1 _3896_ (.A(_1925_),
    .B(net790),
    .C(_1933_),
    .X(_1940_));
 sky130_fd_sc_hd__or3_1 _3897_ (.A(net785),
    .B(net784),
    .C(_1940_),
    .X(_1941_));
 sky130_fd_sc_hd__and3_1 _3898_ (.A(net1410),
    .B(net1408),
    .C(m3_wbd_we_i),
    .X(_1942_));
 sky130_fd_sc_hd__a221o_1 _3899_ (.A1(net1233),
    .A2(m2_wbd_we_i),
    .B1(m1_wbd_we_i),
    .B2(net1174),
    .C1(net1172),
    .X(_1943_));
 sky130_fd_sc_hd__o22a_4 _3900_ (.A1(m0_wbd_we_i),
    .A2(net1166),
    .B1(_1942_),
    .B2(_1943_),
    .X(_1944_));
 sky130_fd_sc_hd__nand2b_1 _3901_ (.A_N(net1389),
    .B(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .Y(_1945_));
 sky130_fd_sc_hd__xor2_4 _3902_ (.A(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[2] ),
    .B(\u_s2.u_sync_wbb.u_cmd_if.rd_ptr[2] ),
    .X(_1946_));
 sky130_fd_sc_hd__xnor2_1 _3903_ (.A(_1945_),
    .B(_1946_),
    .Y(_1947_));
 sky130_fd_sc_hd__xnor2_1 _3904_ (.A(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .B(net1389),
    .Y(_1948_));
 sky130_fd_sc_hd__o21ai_1 _3905_ (.A1(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .A2(_1682_),
    .B1(_1948_),
    .Y(_1949_));
 sky130_fd_sc_hd__and2_1 _3906_ (.A(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .B(_1682_),
    .X(_1950_));
 sky130_fd_sc_hd__o2111a_1 _3907_ (.A1(_1948_),
    .A2(_1950_),
    .B1(_1949_),
    .C1(\u_s2.u_sync_wbb.m_cmd_wr_en ),
    .D1(_1947_),
    .X(_1951_));
 sky130_fd_sc_hd__a22oi_1 _3908_ (.A1(m3_wbd_bry_i),
    .A2(net1177),
    .B1(net1174),
    .B2(net1563),
    .Y(_1952_));
 sky130_fd_sc_hd__o211a_4 _3909_ (.A1(\u_s2.gnt[0] ),
    .A2(_1678_),
    .B1(net1167),
    .C1(_1952_),
    .X(_1953_));
 sky130_fd_sc_hd__nor2_1 _3910_ (.A(_1949_),
    .B(_1950_),
    .Y(_1954_));
 sky130_fd_sc_hd__a211o_4 _3911_ (.A1(_1946_),
    .A2(_1954_),
    .B1(net725),
    .C1(_1951_),
    .X(_1955_));
 sky130_fd_sc_hd__nor3b_4 _3912_ (.A(m1_wbd_adr_i[16]),
    .B(_1766_),
    .C_N(net1176),
    .Y(_1956_));
 sky130_fd_sc_hd__or4b_4 _3913_ (.A(m1_wbd_adr_i[16]),
    .B(_1690_),
    .C(_1766_),
    .D_N(net1176),
    .X(_1957_));
 sky130_fd_sc_hd__nor2_1 _3914_ (.A(m3_wbd_adr_i[16]),
    .B(_1743_),
    .Y(_1958_));
 sky130_fd_sc_hd__or4b_1 _3915_ (.A(m3_wbd_adr_i[16]),
    .B(_1687_),
    .C(_1743_),
    .D_N(net1179),
    .X(_1959_));
 sky130_fd_sc_hd__nor3_4 _3916_ (.A(m2_wbd_adr_i[16]),
    .B(_1777_),
    .C(_1916_),
    .Y(_1960_));
 sky130_fd_sc_hd__or4_1 _3917_ (.A(m2_wbd_adr_i[16]),
    .B(_1688_),
    .C(_1777_),
    .D(_1916_),
    .X(_1961_));
 sky130_fd_sc_hd__or4_4 _3918_ (.A(_1684_),
    .B(m0_wbd_adr_i[16]),
    .C(_1686_),
    .D(_1752_),
    .X(_1962_));
 sky130_fd_sc_hd__o2111a_4 _3919_ (.A1(net1166),
    .A2(_1962_),
    .B1(_1961_),
    .C1(_1959_),
    .D1(_1957_),
    .X(_1963_));
 sky130_fd_sc_hd__nor3_1 _3920_ (.A(m3_wbd_adr_i[16]),
    .B(_1687_),
    .C(_1745_),
    .Y(_1964_));
 sky130_fd_sc_hd__or4b_2 _3921_ (.A(m2_wbd_adr_i[16]),
    .B(_1688_),
    .C(_1779_),
    .D_N(m2_wbd_adr_i[17]),
    .X(_1965_));
 sky130_fd_sc_hd__or4bb_1 _3922_ (.A(m3_wbd_adr_i[16]),
    .B(_1746_),
    .C_N(net1179),
    .D_N(m3_wbd_adr_i[17]),
    .X(_1966_));
 sky130_fd_sc_hd__o22a_4 _3923_ (.A1(_1916_),
    .A2(_1965_),
    .B1(_1966_),
    .B2(_1687_),
    .X(_1967_));
 sky130_fd_sc_hd__and4_2 _3924_ (.A(_1685_),
    .B(m0_wbd_stb_i),
    .C(_1753_),
    .D(_1755_),
    .X(_1968_));
 sky130_fd_sc_hd__and4bb_2 _3925_ (.A_N(_1690_),
    .B_N(_1768_),
    .C(net1176),
    .D(_1760_),
    .X(_1969_));
 sky130_fd_sc_hd__a21oi_4 _3926_ (.A1(net1173),
    .A2(_1968_),
    .B1(_1969_),
    .Y(_1970_));
 sky130_fd_sc_hd__a211oi_4 _3927_ (.A1(net720),
    .A2(net719),
    .B1(net1400),
    .C1(_1955_),
    .Y(_1971_));
 sky130_fd_sc_hd__o31ai_4 _3928_ (.A1(net1400),
    .A2(_1955_),
    .A3(net629),
    .B1(net1826),
    .Y(_1972_));
 sky130_fd_sc_hd__nand2b_2 _3929_ (.A_N(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .B(net1378),
    .Y(_1973_));
 sky130_fd_sc_hd__xnor2_2 _3930_ (.A(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .B(net1379),
    .Y(_1974_));
 sky130_fd_sc_hd__a22oi_1 _3931_ (.A1(_1674_),
    .A2(net1383),
    .B1(\u_s2.u_sync_wbb.wbm_ack_o ),
    .B2(_1974_),
    .Y(_1975_));
 sky130_fd_sc_hd__o21ai_1 _3932_ (.A1(_1674_),
    .A2(net1383),
    .B1(_1974_),
    .Y(_1976_));
 sky130_fd_sc_hd__nand2_1 _3933_ (.A(_1975_),
    .B(_1976_),
    .Y(_1977_));
 sky130_fd_sc_hd__a21o_1 _3934_ (.A1(\u_s2.u_sync_wbb.wbm_ack_o ),
    .A2(_1976_),
    .B1(_1975_),
    .X(_1978_));
 sky130_fd_sc_hd__xnor2_4 _3935_ (.A(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[2] ),
    .B(\u_s2.u_sync_wbb.u_resp_if.rd_ptr[2] ),
    .Y(_1979_));
 sky130_fd_sc_hd__xnor2_4 _3936_ (.A(_1973_),
    .B(_1979_),
    .Y(_1980_));
 sky130_fd_sc_hd__a31o_4 _3937_ (.A1(_1977_),
    .A2(_1978_),
    .A3(_1980_),
    .B1(net725),
    .X(_1981_));
 sky130_fd_sc_hd__nor2_2 _3938_ (.A(_1680_),
    .B(_1981_),
    .Y(_1982_));
 sky130_fd_sc_hd__nor2_2 _3939_ (.A(_1681_),
    .B(_1955_),
    .Y(_1983_));
 sky130_fd_sc_hd__nor2_1 _3940_ (.A(_1982_),
    .B(_1983_),
    .Y(_1984_));
 sky130_fd_sc_hd__or4_2 _3941_ (.A(\u_s2.u_sync_wbb.m_bl_cnt[7] ),
    .B(\u_s2.u_sync_wbb.m_bl_cnt[6] ),
    .C(\u_s2.u_sync_wbb.m_bl_cnt[9] ),
    .D(\u_s2.u_sync_wbb.m_bl_cnt[8] ),
    .X(_1985_));
 sky130_fd_sc_hd__or4_1 _3942_ (.A(_1679_),
    .B(\u_s2.u_sync_wbb.m_bl_cnt[1] ),
    .C(\u_s2.u_sync_wbb.m_bl_cnt[3] ),
    .D(\u_s2.u_sync_wbb.m_bl_cnt[4] ),
    .X(_1986_));
 sky130_fd_sc_hd__or4_4 _3943_ (.A(\u_s2.u_sync_wbb.m_bl_cnt[2] ),
    .B(\u_s2.u_sync_wbb.m_bl_cnt[5] ),
    .C(_1985_),
    .D(_1986_),
    .X(_1987_));
 sky130_fd_sc_hd__inv_2 _3944_ (.A(_1987_),
    .Y(_1988_));
 sky130_fd_sc_hd__nand2_1 _3945_ (.A(net726),
    .B(_1971_),
    .Y(_1989_));
 sky130_fd_sc_hd__o32a_1 _3946_ (.A1(_1691_),
    .A2(_1941_),
    .A3(_1989_),
    .B1(_1987_),
    .B2(_1984_),
    .X(_1990_));
 sky130_fd_sc_hd__nand2_1 _3947_ (.A(_1972_),
    .B(_1990_),
    .Y(_0006_));
 sky130_fd_sc_hd__o21ai_1 _3948_ (.A1(_1981_),
    .A2(_1987_),
    .B1(\u_s2.u_sync_wbb.m_state[1] ),
    .Y(_1991_));
 sky130_fd_sc_hd__a2111o_1 _3949_ (.A1(net720),
    .A2(net719),
    .B1(net1400),
    .C1(net726),
    .D1(_1955_),
    .X(_1992_));
 sky130_fd_sc_hd__o21ai_1 _3950_ (.A1(_1691_),
    .A2(net583),
    .B1(_1991_),
    .Y(_0007_));
 sky130_fd_sc_hd__o21a_1 _3951_ (.A1(_1955_),
    .A2(_1987_),
    .B1(\u_s2.u_sync_wbb.m_state[2] ),
    .X(_1993_));
 sky130_fd_sc_hd__and4_1 _3952_ (.A(\u_s2.u_sync_wbb.m_state[0] ),
    .B(_1941_),
    .C(net726),
    .D(_1971_),
    .X(_1994_));
 sky130_fd_sc_hd__or2_1 _3953_ (.A(_1993_),
    .B(_1994_),
    .X(_0008_));
 sky130_fd_sc_hd__and4_1 _3954_ (.A(\u_s1.u_sync_wbb.m_state[0] ),
    .B(net732),
    .C(_1876_),
    .D(_1883_),
    .X(_1995_));
 sky130_fd_sc_hd__o21a_1 _3955_ (.A1(_1850_),
    .A2(_1898_),
    .B1(\u_s1.u_sync_wbb.m_state[2] ),
    .X(_1996_));
 sky130_fd_sc_hd__or2_1 _3956_ (.A(_1995_),
    .B(_1996_),
    .X(_0005_));
 sky130_fd_sc_hd__a2111o_2 _3957_ (.A1(_1721_),
    .A2(_1723_),
    .B1(_1734_),
    .C1(_1806_),
    .D1(\u_s0.u_sync_wbb.wbm_lack_o ),
    .X(_1997_));
 sky130_fd_sc_hd__a21oi_4 _3958_ (.A1(_1759_),
    .A2(_1782_),
    .B1(_1997_),
    .Y(_1998_));
 sky130_fd_sc_hd__or2_1 _3959_ (.A(_1820_),
    .B(_1827_),
    .X(_1999_));
 sky130_fd_sc_hd__a22o_1 _3960_ (.A1(\u_s0.u_sync_wbb.m_state[0] ),
    .A2(net580),
    .B1(_1999_),
    .B2(\u_s0.u_sync_wbb.m_state[1] ),
    .X(_0001_));
 sky130_fd_sc_hd__nand2b_1 _3961_ (.A_N(\u_dcg_s2.cfg_mode_ss[0] ),
    .B(\u_dcg_s2.cfg_mode_ss[1] ),
    .Y(\u_dcg_s2.clk_enb ));
 sky130_fd_sc_hd__o21ai_1 _3962_ (.A1(_1892_),
    .A2(_1898_),
    .B1(\u_s1.u_sync_wbb.m_state[1] ),
    .Y(_2000_));
 sky130_fd_sc_hd__and4b_4 _3963_ (.A_N(net732),
    .B(_1849_),
    .C(net807),
    .D(_1694_),
    .X(_2001_));
 sky130_fd_sc_hd__nand2_1 _3964_ (.A(net630),
    .B(_2001_),
    .Y(_2002_));
 sky130_fd_sc_hd__o21ai_1 _3965_ (.A1(_1695_),
    .A2(_2002_),
    .B1(_2000_),
    .Y(_0004_));
 sky130_fd_sc_hd__nand2b_2 _3966_ (.A_N(\u_dcg_s1.cfg_mode_ss[0] ),
    .B(\u_dcg_s1.cfg_mode_ss[1] ),
    .Y(\u_dcg_s1.clk_enb ));
 sky130_fd_sc_hd__nand2b_1 _3967_ (.A_N(\u_dcg_riscv.cfg_mode_ss[0] ),
    .B(net1492),
    .Y(\u_dcg_riscv.clk_enb ));
 sky130_fd_sc_hd__nand2b_1 _3968_ (.A_N(\u_dcg_peri.cfg_mode_ss[0] ),
    .B(\u_dcg_peri.cfg_mode_ss[1] ),
    .Y(\u_dcg_peri.clk_enb ));
 sky130_fd_sc_hd__or3_1 _3969_ (.A(_1946_),
    .B(_1949_),
    .C(_1950_),
    .X(_2003_));
 sky130_fd_sc_hd__mux4_1 _3970_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][50] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][50] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][50] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][50] ),
    .S0(net1396),
    .S1(net1389),
    .X(_2004_));
 sky130_fd_sc_hd__mux2_2 _3971_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[50] ),
    .A1(_2004_),
    .S(net716),
    .X(net476));
 sky130_fd_sc_hd__or4b_1 _3972_ (.A(_1839_),
    .B(_1841_),
    .C(_1844_),
    .D_N(_1842_),
    .X(_2005_));
 sky130_fd_sc_hd__mux4_2 _3973_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][50] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][50] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][50] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][50] ),
    .S0(net1362),
    .S1(net1355),
    .X(_2006_));
 sky130_fd_sc_hd__mux2_2 _3974_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[50] ),
    .A1(_2006_),
    .S(net774),
    .X(net427));
 sky130_fd_sc_hd__mux4_2 _3975_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][50] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][50] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][50] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][50] ),
    .S0(net1339),
    .S1(net1329),
    .X(_2007_));
 sky130_fd_sc_hd__mux2_1 _3976_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[50] ),
    .A1(_2007_),
    .S(net831),
    .X(net380));
 sky130_fd_sc_hd__a21o_4 _3977_ (.A1(_1709_),
    .A2(net717),
    .B1(\u_s2.u_sync_wbb.wbs_burst ),
    .X(net438));
 sky130_fd_sc_hd__a21o_4 _3978_ (.A1(_1702_),
    .A2(net775),
    .B1(\u_s1.u_sync_wbb.wbs_burst ),
    .X(net389));
 sky130_fd_sc_hd__nor2_4 _3979_ (.A(_1689_),
    .B(_1764_),
    .Y(_2008_));
 sky130_fd_sc_hd__o31a_1 _3980_ (.A1(_1689_),
    .A2(_1690_),
    .A3(_1764_),
    .B1(net1278),
    .X(_2009_));
 sky130_fd_sc_hd__or2_1 _3981_ (.A(net1275),
    .B(_2009_),
    .X(_2010_));
 sky130_fd_sc_hd__nor2_1 _3982_ (.A(_1775_),
    .B(_1776_),
    .Y(_2011_));
 sky130_fd_sc_hd__nand2_1 _3983_ (.A(m2_wbd_stb_i),
    .B(net1161),
    .Y(_2012_));
 sky130_fd_sc_hd__and2_1 _3984_ (.A(net1277),
    .B(net1274),
    .X(_2013_));
 sky130_fd_sc_hd__nor2_1 _3985_ (.A(_1741_),
    .B(_1742_),
    .Y(_2014_));
 sky130_fd_sc_hd__or4_1 _3986_ (.A(_1688_),
    .B(net1277),
    .C(_1776_),
    .D(_1778_),
    .X(_2015_));
 sky130_fd_sc_hd__or3_1 _3987_ (.A(_1687_),
    .B(_1742_),
    .C(_1744_),
    .X(_2016_));
 sky130_fd_sc_hd__o31a_1 _3988_ (.A1(net1219),
    .A2(net1210),
    .A3(_2016_),
    .B1(_2015_),
    .X(_2017_));
 sky130_fd_sc_hd__nand2_1 _3989_ (.A(_2010_),
    .B(_2017_),
    .Y(_2018_));
 sky130_fd_sc_hd__nor2_4 _3990_ (.A(net1278),
    .B(net1275),
    .Y(_2019_));
 sky130_fd_sc_hd__or2_1 _3991_ (.A(net1276),
    .B(net1274),
    .X(_2020_));
 sky130_fd_sc_hd__nor3_4 _3992_ (.A(_1684_),
    .B(_1685_),
    .C(_1752_),
    .Y(_2021_));
 sky130_fd_sc_hd__nand2_1 _3993_ (.A(m0_wbd_stb_i),
    .B(net1147),
    .Y(_2022_));
 sky130_fd_sc_hd__a22o_1 _3994_ (.A1(_2010_),
    .A2(_2017_),
    .B1(_2019_),
    .B2(_2022_),
    .X(_2023_));
 sky130_fd_sc_hd__or2_4 _3995_ (.A(\u_reg.reg_ack ),
    .B(net711),
    .X(_2024_));
 sky130_fd_sc_hd__inv_2 _3996_ (.A(net627),
    .Y(_0009_));
 sky130_fd_sc_hd__a22o_1 _3997_ (.A1(net1366),
    .A2(net804),
    .B1(net1158),
    .B2(\u_reg.reg_ack ),
    .X(_2025_));
 sky130_fd_sc_hd__a22o_1 _3998_ (.A1(\u_s0.u_sync_wbb.wbm_lack_o ),
    .A2(net812),
    .B1(net722),
    .B2(net1401),
    .X(_2026_));
 sky130_fd_sc_hd__or2_1 _3999_ (.A(_2025_),
    .B(_2026_),
    .X(net263));
 sky130_fd_sc_hd__a22o_1 _4000_ (.A1(net1367),
    .A2(net806),
    .B1(net1159),
    .B2(\u_reg.reg_ack ),
    .X(_2027_));
 sky130_fd_sc_hd__a22o_1 _4001_ (.A1(\u_s0.u_sync_wbb.wbm_ack_o ),
    .A2(net811),
    .B1(net724),
    .B2(net1402),
    .X(_2028_));
 sky130_fd_sc_hd__or2_1 _4002_ (.A(_2027_),
    .B(_2028_),
    .X(net230));
 sky130_fd_sc_hd__mux4_1 _4003_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][0] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][0] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][0] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][0] ),
    .S0(net1319),
    .S1(net1314),
    .X(_2029_));
 sky130_fd_sc_hd__a22o_1 _4004_ (.A1(net1312),
    .A2(net1159),
    .B1(net1142),
    .B2(net811),
    .X(_2030_));
 sky130_fd_sc_hd__mux4_2 _4005_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][0] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][0] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][0] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][0] ),
    .S0(net1383),
    .S1(net1379),
    .X(_2031_));
 sky130_fd_sc_hd__mux4_2 _4006_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][0] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][0] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][0] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][0] ),
    .S0(net1349),
    .S1(net1345),
    .X(_2032_));
 sky130_fd_sc_hd__a22o_1 _4007_ (.A1(net723),
    .A2(net1140),
    .B1(net1138),
    .B2(net805),
    .X(_2033_));
 sky130_fd_sc_hd__or2_1 _4008_ (.A(_2030_),
    .B(_2033_),
    .X(net231));
 sky130_fd_sc_hd__mux4_2 _4009_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][1] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][1] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][1] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][1] ),
    .S0(net1350),
    .S1(net1346),
    .X(_2034_));
 sky130_fd_sc_hd__a22o_1 _4010_ (.A1(\u_reg.reg_rdata[1] ),
    .A2(net1159),
    .B1(net1137),
    .B2(net806),
    .X(_2035_));
 sky130_fd_sc_hd__mux4_2 _4011_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][1] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][1] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][1] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][1] ),
    .S0(net1321),
    .S1(net1316),
    .X(_2036_));
 sky130_fd_sc_hd__mux4_2 _4012_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][1] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][1] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][1] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][1] ),
    .S0(net1382),
    .S1(net1378),
    .X(_2037_));
 sky130_fd_sc_hd__a22o_1 _4013_ (.A1(net811),
    .A2(_2036_),
    .B1(net1135),
    .B2(net724),
    .X(_2038_));
 sky130_fd_sc_hd__or2_1 _4014_ (.A(_2035_),
    .B(_2038_),
    .X(net242));
 sky130_fd_sc_hd__mux4_1 _4015_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][2] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][2] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][2] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][2] ),
    .S0(net1322),
    .S1(net1315),
    .X(_2039_));
 sky130_fd_sc_hd__a22o_1 _4016_ (.A1(\u_reg.reg_rdata[2] ),
    .A2(net1159),
    .B1(net1134),
    .B2(net811),
    .X(_2040_));
 sky130_fd_sc_hd__mux4_2 _4017_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][2] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][2] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][2] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][2] ),
    .S0(net1382),
    .S1(net1378),
    .X(_2041_));
 sky130_fd_sc_hd__mux4_2 _4018_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][2] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][2] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][2] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][2] ),
    .S0(net1350),
    .S1(net1346),
    .X(_2042_));
 sky130_fd_sc_hd__a22o_1 _4019_ (.A1(net724),
    .A2(net1131),
    .B1(net1129),
    .B2(net806),
    .X(_2043_));
 sky130_fd_sc_hd__or2_1 _4020_ (.A(_2040_),
    .B(_2043_),
    .X(net253));
 sky130_fd_sc_hd__mux4_2 _4021_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][3] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][3] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][3] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][3] ),
    .S0(net1348),
    .S1(net1344),
    .X(_2044_));
 sky130_fd_sc_hd__a22o_1 _4022_ (.A1(\u_reg.reg_rdata[3] ),
    .A2(net1159),
    .B1(net1128),
    .B2(net805),
    .X(_2045_));
 sky130_fd_sc_hd__mux4_2 _4023_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][3] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][3] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][3] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][3] ),
    .S0(net1321),
    .S1(net1316),
    .X(_2046_));
 sky130_fd_sc_hd__mux4_2 _4024_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][3] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][3] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][3] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][3] ),
    .S0(net1382),
    .S1(net1378),
    .X(_2047_));
 sky130_fd_sc_hd__a22o_1 _4025_ (.A1(net811),
    .A2(_2046_),
    .B1(net1126),
    .B2(net723),
    .X(_2048_));
 sky130_fd_sc_hd__or2_1 _4026_ (.A(_2045_),
    .B(_2048_),
    .X(net256));
 sky130_fd_sc_hd__mux4_1 _4027_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][4] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][4] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][4] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][4] ),
    .S0(net1320),
    .S1(net1317),
    .X(_2049_));
 sky130_fd_sc_hd__a22o_1 _4028_ (.A1(net1311),
    .A2(net1159),
    .B1(net1125),
    .B2(net811),
    .X(_2050_));
 sky130_fd_sc_hd__mux4_2 _4029_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][4] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][4] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][4] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][4] ),
    .S0(net1382),
    .S1(net1378),
    .X(_2051_));
 sky130_fd_sc_hd__mux4_2 _4030_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][4] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][4] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][4] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][4] ),
    .S0(net1349),
    .S1(net1345),
    .X(_2052_));
 sky130_fd_sc_hd__a22o_1 _4031_ (.A1(net724),
    .A2(net1123),
    .B1(net1122),
    .B2(net806),
    .X(_2053_));
 sky130_fd_sc_hd__or2_1 _4032_ (.A(_2050_),
    .B(_2053_),
    .X(net257));
 sky130_fd_sc_hd__mux4_2 _4033_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][5] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][5] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][5] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][5] ),
    .S0(net1350),
    .S1(net1346),
    .X(_2054_));
 sky130_fd_sc_hd__a22o_1 _4034_ (.A1(net1310),
    .A2(net1159),
    .B1(net1120),
    .B2(net805),
    .X(_2055_));
 sky130_fd_sc_hd__mux4_2 _4035_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][5] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][5] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][5] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][5] ),
    .S0(net1320),
    .S1(net1317),
    .X(_2056_));
 sky130_fd_sc_hd__mux4_2 _4036_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][5] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][5] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][5] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][5] ),
    .S0(net1382),
    .S1(net1378),
    .X(_2057_));
 sky130_fd_sc_hd__a22o_1 _4037_ (.A1(net811),
    .A2(net1119),
    .B1(net1116),
    .B2(net723),
    .X(_2058_));
 sky130_fd_sc_hd__or2_1 _4038_ (.A(_2055_),
    .B(_2058_),
    .X(net258));
 sky130_fd_sc_hd__mux4_2 _4039_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][6] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][6] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][6] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][6] ),
    .S0(net1350),
    .S1(net1346),
    .X(_2059_));
 sky130_fd_sc_hd__a22o_1 _4040_ (.A1(\u_reg.reg_rdata[6] ),
    .A2(net1158),
    .B1(net1115),
    .B2(net805),
    .X(_2060_));
 sky130_fd_sc_hd__mux4_1 _4041_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][6] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][6] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][6] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][6] ),
    .S0(net1320),
    .S1(net1315),
    .X(_2061_));
 sky130_fd_sc_hd__mux4_2 _4042_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][6] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][6] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][6] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][6] ),
    .S0(net1382),
    .S1(net1378),
    .X(_2062_));
 sky130_fd_sc_hd__a22o_1 _4043_ (.A1(net812),
    .A2(net1114),
    .B1(net1112),
    .B2(net723),
    .X(_2063_));
 sky130_fd_sc_hd__or2_1 _4044_ (.A(_2060_),
    .B(_2063_),
    .X(net259));
 sky130_fd_sc_hd__mux4_2 _4045_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][7] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][7] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][7] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][7] ),
    .S0(net1322),
    .S1(net1315),
    .X(_2064_));
 sky130_fd_sc_hd__a22o_1 _4046_ (.A1(net1309),
    .A2(net1159),
    .B1(net1111),
    .B2(net811),
    .X(_2065_));
 sky130_fd_sc_hd__mux4_1 _4047_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][7] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][7] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][7] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][7] ),
    .S0(net1380),
    .S1(net1376),
    .X(_2066_));
 sky130_fd_sc_hd__mux4_2 _4048_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][7] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][7] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][7] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][7] ),
    .S0(net1349),
    .S1(net1345),
    .X(_2067_));
 sky130_fd_sc_hd__a22o_1 _4049_ (.A1(net723),
    .A2(net1109),
    .B1(net1108),
    .B2(net805),
    .X(_2068_));
 sky130_fd_sc_hd__or2_1 _4050_ (.A(_2065_),
    .B(_2068_),
    .X(net260));
 sky130_fd_sc_hd__mux4_2 _4051_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][8] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][8] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][8] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][8] ),
    .S0(net1349),
    .S1(net1346),
    .X(_2069_));
 sky130_fd_sc_hd__a22o_1 _4052_ (.A1(net1308),
    .A2(net1160),
    .B1(net1106),
    .B2(net806),
    .X(_2070_));
 sky130_fd_sc_hd__mux4_2 _4053_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][8] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][8] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][8] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][8] ),
    .S0(net1321),
    .S1(net1316),
    .X(_2071_));
 sky130_fd_sc_hd__mux4_1 _4054_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][8] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][8] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][8] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][8] ),
    .S0(net1383),
    .S1(net1379),
    .X(_2072_));
 sky130_fd_sc_hd__a22o_1 _4055_ (.A1(net811),
    .A2(_2071_),
    .B1(net1103),
    .B2(net724),
    .X(_2073_));
 sky130_fd_sc_hd__or2_1 _4056_ (.A(_2070_),
    .B(_2073_),
    .X(net261));
 sky130_fd_sc_hd__mux4_2 _4057_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][9] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][9] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][9] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][9] ),
    .S0(net1349),
    .S1(net1345),
    .X(_2074_));
 sky130_fd_sc_hd__a22o_1 _4058_ (.A1(net1307),
    .A2(net1159),
    .B1(net1102),
    .B2(net806),
    .X(_2075_));
 sky130_fd_sc_hd__mux4_2 _4059_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][9] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][9] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][9] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][9] ),
    .S0(net1321),
    .S1(net1316),
    .X(_2076_));
 sky130_fd_sc_hd__mux4_2 _4060_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][9] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][9] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][9] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][9] ),
    .S0(net1383),
    .S1(net1379),
    .X(_2077_));
 sky130_fd_sc_hd__a22o_1 _4061_ (.A1(_1780_),
    .A2(net1101),
    .B1(net1099),
    .B2(net724),
    .X(_2078_));
 sky130_fd_sc_hd__or2_1 _4062_ (.A(_2075_),
    .B(_2078_),
    .X(net262));
 sky130_fd_sc_hd__mux4_2 _4063_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][10] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][10] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][10] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][10] ),
    .S0(net1347),
    .S1(net1343),
    .X(_2079_));
 sky130_fd_sc_hd__a22o_1 _4064_ (.A1(net1306),
    .A2(net1160),
    .B1(net1098),
    .B2(net806),
    .X(_2080_));
 sky130_fd_sc_hd__mux4_2 _4065_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][10] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][10] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][10] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][10] ),
    .S0(net1321),
    .S1(net1316),
    .X(_2081_));
 sky130_fd_sc_hd__mux4_2 _4066_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][10] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][10] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][10] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][10] ),
    .S0(net1382),
    .S1(net1378),
    .X(_2082_));
 sky130_fd_sc_hd__a22o_1 _4067_ (.A1(net812),
    .A2(net1097),
    .B1(net1094),
    .B2(net724),
    .X(_2083_));
 sky130_fd_sc_hd__or2_1 _4068_ (.A(_2080_),
    .B(_2083_),
    .X(net232));
 sky130_fd_sc_hd__mux4_1 _4069_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][11] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][11] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][11] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][11] ),
    .S0(net1319),
    .S1(net1314),
    .X(_2084_));
 sky130_fd_sc_hd__a22o_1 _4070_ (.A1(net1305),
    .A2(net1158),
    .B1(net1093),
    .B2(net809),
    .X(_2085_));
 sky130_fd_sc_hd__mux4_2 _4071_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][11] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][11] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][11] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][11] ),
    .S0(net1381),
    .S1(net1377),
    .X(_2086_));
 sky130_fd_sc_hd__mux4_1 _4072_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][11] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][11] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][11] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][11] ),
    .S0(net1347),
    .S1(net1344),
    .X(_2087_));
 sky130_fd_sc_hd__a22o_1 _4073_ (.A1(net721),
    .A2(net1092),
    .B1(net1091),
    .B2(net803),
    .X(_2088_));
 sky130_fd_sc_hd__or2_1 _4074_ (.A(_2085_),
    .B(_2088_),
    .X(net233));
 sky130_fd_sc_hd__mux4_2 _4075_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][12] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][12] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][12] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][12] ),
    .S0(net1348),
    .S1(net1344),
    .X(_2089_));
 sky130_fd_sc_hd__a22o_1 _4076_ (.A1(net1304),
    .A2(net1160),
    .B1(net1090),
    .B2(net805),
    .X(_2090_));
 sky130_fd_sc_hd__mux4_2 _4077_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][12] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][12] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][12] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][12] ),
    .S0(net1318),
    .S1(net1313),
    .X(_2091_));
 sky130_fd_sc_hd__mux4_1 _4078_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][12] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][12] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][12] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][12] ),
    .S0(net1382),
    .S1(net1378),
    .X(_2092_));
 sky130_fd_sc_hd__a22o_1 _4079_ (.A1(net812),
    .A2(net1089),
    .B1(net1086),
    .B2(net723),
    .X(_2093_));
 sky130_fd_sc_hd__or2_1 _4080_ (.A(_2090_),
    .B(_2093_),
    .X(net234));
 sky130_fd_sc_hd__mux4_2 _4081_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][13] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][13] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][13] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][13] ),
    .S0(net1351),
    .S1(net1344),
    .X(_2094_));
 sky130_fd_sc_hd__a22o_1 _4082_ (.A1(net1302),
    .A2(net1158),
    .B1(net1085),
    .B2(net805),
    .X(_2095_));
 sky130_fd_sc_hd__mux4_2 _4083_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][13] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][13] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][13] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][13] ),
    .S0(net1319),
    .S1(net1314),
    .X(_2096_));
 sky130_fd_sc_hd__mux4_2 _4084_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][13] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][13] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][13] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][13] ),
    .S0(net1380),
    .S1(net1376),
    .X(_2097_));
 sky130_fd_sc_hd__a22o_1 _4085_ (.A1(net812),
    .A2(net1084),
    .B1(net1082),
    .B2(net723),
    .X(_2098_));
 sky130_fd_sc_hd__or2_1 _4086_ (.A(_2095_),
    .B(_2098_),
    .X(net235));
 sky130_fd_sc_hd__mux4_2 _4087_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][14] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][14] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][14] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][14] ),
    .S0(net1349),
    .S1(net1345),
    .X(_2099_));
 sky130_fd_sc_hd__a22o_1 _4088_ (.A1(net1300),
    .A2(net1160),
    .B1(net1081),
    .B2(net805),
    .X(_2100_));
 sky130_fd_sc_hd__mux4_2 _4089_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][14] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][14] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][14] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][14] ),
    .S0(net1318),
    .S1(net1313),
    .X(_2101_));
 sky130_fd_sc_hd__mux4_2 _4090_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][14] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][14] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][14] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][14] ),
    .S0(net1381),
    .S1(net1377),
    .X(_2102_));
 sky130_fd_sc_hd__a22o_1 _4091_ (.A1(net812),
    .A2(net1080),
    .B1(net1078),
    .B2(net723),
    .X(_2103_));
 sky130_fd_sc_hd__or2_1 _4092_ (.A(_2100_),
    .B(_2103_),
    .X(net236));
 sky130_fd_sc_hd__mux4_2 _4093_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][15] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][15] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][15] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][15] ),
    .S0(net1320),
    .S1(net1315),
    .X(_2104_));
 sky130_fd_sc_hd__a22o_1 _4094_ (.A1(net1298),
    .A2(net1160),
    .B1(net1077),
    .B2(net812),
    .X(_2105_));
 sky130_fd_sc_hd__mux4_2 _4095_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][15] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][15] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][15] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][15] ),
    .S0(net1383),
    .S1(net1379),
    .X(_2106_));
 sky130_fd_sc_hd__mux4_1 _4096_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][15] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][15] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][15] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][15] ),
    .S0(net1349),
    .S1(net1345),
    .X(_2107_));
 sky130_fd_sc_hd__a22o_1 _4097_ (.A1(net721),
    .A2(net1075),
    .B1(net1073),
    .B2(net803),
    .X(_2108_));
 sky130_fd_sc_hd__or2_1 _4098_ (.A(_2105_),
    .B(_2108_),
    .X(net237));
 sky130_fd_sc_hd__mux4_2 _4099_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][16] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][16] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][16] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][16] ),
    .S0(net1349),
    .S1(net1345),
    .X(_2109_));
 sky130_fd_sc_hd__a22o_1 _4100_ (.A1(net1296),
    .A2(net1159),
    .B1(net1071),
    .B2(net805),
    .X(_2110_));
 sky130_fd_sc_hd__mux4_2 _4101_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][16] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][16] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][16] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][16] ),
    .S0(net1318),
    .S1(net1313),
    .X(_2111_));
 sky130_fd_sc_hd__mux4_2 _4102_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][16] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][16] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][16] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][16] ),
    .S0(net1380),
    .S1(net1376),
    .X(_2112_));
 sky130_fd_sc_hd__a22o_1 _4103_ (.A1(net811),
    .A2(net1070),
    .B1(net1068),
    .B2(net723),
    .X(_2113_));
 sky130_fd_sc_hd__or2_1 _4104_ (.A(_2110_),
    .B(_2113_),
    .X(net238));
 sky130_fd_sc_hd__mux4_1 _4105_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][17] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][17] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][17] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][17] ),
    .S0(net1348),
    .S1(net1344),
    .X(_2114_));
 sky130_fd_sc_hd__a22o_1 _4106_ (.A1(net1295),
    .A2(net1160),
    .B1(net1067),
    .B2(net805),
    .X(_2115_));
 sky130_fd_sc_hd__mux4_1 _4107_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][17] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][17] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][17] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][17] ),
    .S0(net1320),
    .S1(net1315),
    .X(_2116_));
 sky130_fd_sc_hd__mux4_2 _4108_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][17] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][17] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][17] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][17] ),
    .S0(net1382),
    .S1(net1378),
    .X(_2117_));
 sky130_fd_sc_hd__a22o_1 _4109_ (.A1(net812),
    .A2(net1066),
    .B1(net1064),
    .B2(net723),
    .X(_2118_));
 sky130_fd_sc_hd__or2_1 _4110_ (.A(_2115_),
    .B(_2118_),
    .X(net239));
 sky130_fd_sc_hd__mux4_1 _4111_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][18] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][18] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][18] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][18] ),
    .S0(net1322),
    .S1(net1316),
    .X(_2119_));
 sky130_fd_sc_hd__a22o_1 _4112_ (.A1(\u_reg.reg_rdata[18] ),
    .A2(net1158),
    .B1(net1063),
    .B2(net812),
    .X(_2120_));
 sky130_fd_sc_hd__mux4_2 _4113_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][18] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][18] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][18] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][18] ),
    .S0(net1383),
    .S1(net1379),
    .X(_2121_));
 sky130_fd_sc_hd__mux4_2 _4114_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][18] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][18] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][18] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][18] ),
    .S0(net1349),
    .S1(net1345),
    .X(_2122_));
 sky130_fd_sc_hd__a22o_1 _4115_ (.A1(net722),
    .A2(net1060),
    .B1(net1058),
    .B2(net804),
    .X(_2123_));
 sky130_fd_sc_hd__or2_1 _4116_ (.A(_2120_),
    .B(_2123_),
    .X(net240));
 sky130_fd_sc_hd__mux4_1 _4117_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][19] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][19] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][19] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][19] ),
    .S0(net1347),
    .S1(net1343),
    .X(_2124_));
 sky130_fd_sc_hd__a22o_1 _4118_ (.A1(\u_reg.reg_rdata[19] ),
    .A2(net1158),
    .B1(net1057),
    .B2(net804),
    .X(_2125_));
 sky130_fd_sc_hd__mux4_2 _4119_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][19] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][19] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][19] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][19] ),
    .S0(net1318),
    .S1(net1313),
    .X(_2126_));
 sky130_fd_sc_hd__mux4_2 _4120_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][19] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][19] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][19] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][19] ),
    .S0(net1380),
    .S1(net1376),
    .X(_2127_));
 sky130_fd_sc_hd__a22o_1 _4121_ (.A1(net809),
    .A2(_2126_),
    .B1(net1056),
    .B2(net722),
    .X(_2128_));
 sky130_fd_sc_hd__or2_1 _4122_ (.A(_2125_),
    .B(_2128_),
    .X(net241));
 sky130_fd_sc_hd__mux4_2 _4123_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][20] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][20] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][20] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][20] ),
    .S0(net1348),
    .S1(net1344),
    .X(_2129_));
 sky130_fd_sc_hd__a22o_1 _4124_ (.A1(net1293),
    .A2(net1161),
    .B1(net1055),
    .B2(net803),
    .X(_2130_));
 sky130_fd_sc_hd__mux4_2 _4125_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][20] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][20] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][20] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][20] ),
    .S0(net1318),
    .S1(net1313),
    .X(_2131_));
 sky130_fd_sc_hd__mux4_2 _4126_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][20] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][20] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][20] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][20] ),
    .S0(net1383),
    .S1(net1379),
    .X(_2132_));
 sky130_fd_sc_hd__a22o_1 _4127_ (.A1(net809),
    .A2(net1054),
    .B1(net1051),
    .B2(net721),
    .X(_2133_));
 sky130_fd_sc_hd__or2_1 _4128_ (.A(_2130_),
    .B(_2133_),
    .X(net243));
 sky130_fd_sc_hd__mux4_2 _4129_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][21] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][21] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][21] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][21] ),
    .S0(net1320),
    .S1(net1315),
    .X(_2134_));
 sky130_fd_sc_hd__a22o_1 _4130_ (.A1(net1291),
    .A2(net1161),
    .B1(net1050),
    .B2(net809),
    .X(_2135_));
 sky130_fd_sc_hd__mux4_2 _4131_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][21] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][21] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][21] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][21] ),
    .S0(net1380),
    .S1(net1376),
    .X(_2136_));
 sky130_fd_sc_hd__mux4_2 _4132_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][21] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][21] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][21] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][21] ),
    .S0(net1348),
    .S1(net1344),
    .X(_2137_));
 sky130_fd_sc_hd__a22o_1 _4133_ (.A1(net721),
    .A2(net1048),
    .B1(net1047),
    .B2(net803),
    .X(_2138_));
 sky130_fd_sc_hd__or2_1 _4134_ (.A(_2135_),
    .B(_2138_),
    .X(net244));
 sky130_fd_sc_hd__mux4_2 _4135_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][22] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][22] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][22] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][22] ),
    .S0(net1318),
    .S1(net1313),
    .X(_2139_));
 sky130_fd_sc_hd__a22o_1 _4136_ (.A1(net1290),
    .A2(net1161),
    .B1(net1046),
    .B2(net809),
    .X(_2140_));
 sky130_fd_sc_hd__mux4_2 _4137_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][22] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][22] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][22] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][22] ),
    .S0(net1381),
    .S1(net1377),
    .X(_2141_));
 sky130_fd_sc_hd__mux4_2 _4138_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][22] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][22] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][22] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][22] ),
    .S0(net1347),
    .S1(net1343),
    .X(_2142_));
 sky130_fd_sc_hd__a22o_1 _4139_ (.A1(net721),
    .A2(net1044),
    .B1(net1043),
    .B2(net803),
    .X(_2143_));
 sky130_fd_sc_hd__or2_1 _4140_ (.A(_2140_),
    .B(_2143_),
    .X(net245));
 sky130_fd_sc_hd__mux4_2 _4141_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][23] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][23] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][23] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][23] ),
    .S0(net1319),
    .S1(net1314),
    .X(_2144_));
 sky130_fd_sc_hd__a22o_1 _4142_ (.A1(\u_reg.reg_rdata[23] ),
    .A2(net1161),
    .B1(_2144_),
    .B2(net810),
    .X(_2145_));
 sky130_fd_sc_hd__mux4_1 _4143_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][23] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][23] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][23] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][23] ),
    .S0(net1383),
    .S1(net1379),
    .X(_2146_));
 sky130_fd_sc_hd__mux4_2 _4144_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][23] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][23] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][23] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][23] ),
    .S0(net1347),
    .S1(net1343),
    .X(_2147_));
 sky130_fd_sc_hd__a22o_1 _4145_ (.A1(net721),
    .A2(net1040),
    .B1(net1039),
    .B2(net803),
    .X(_2148_));
 sky130_fd_sc_hd__or2_1 _4146_ (.A(_2145_),
    .B(_2148_),
    .X(net246));
 sky130_fd_sc_hd__mux4_1 _4147_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][24] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][24] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][24] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][24] ),
    .S0(net1321),
    .S1(net1316),
    .X(_2149_));
 sky130_fd_sc_hd__a22o_1 _4148_ (.A1(net1289),
    .A2(net1158),
    .B1(net1038),
    .B2(net809),
    .X(_2150_));
 sky130_fd_sc_hd__mux4_2 _4149_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][24] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][24] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][24] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][24] ),
    .S0(net1381),
    .S1(net1377),
    .X(_2151_));
 sky130_fd_sc_hd__mux4_2 _4150_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][24] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][24] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][24] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][24] ),
    .S0(net1347),
    .S1(net1343),
    .X(_2152_));
 sky130_fd_sc_hd__a22o_1 _4151_ (.A1(net722),
    .A2(net1037),
    .B1(net1036),
    .B2(net804),
    .X(_2153_));
 sky130_fd_sc_hd__or2_1 _4152_ (.A(_2150_),
    .B(_2153_),
    .X(net247));
 sky130_fd_sc_hd__mux4_2 _4153_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][25] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][25] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][25] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][25] ),
    .S0(net1348),
    .S1(net1343),
    .X(_2154_));
 sky130_fd_sc_hd__a22o_1 _4154_ (.A1(net1288),
    .A2(net1158),
    .B1(net1035),
    .B2(net804),
    .X(_2155_));
 sky130_fd_sc_hd__mux4_2 _4155_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][25] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][25] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][25] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][25] ),
    .S0(net1321),
    .S1(net1316),
    .X(_2156_));
 sky130_fd_sc_hd__mux4_2 _4156_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][25] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][25] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][25] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][25] ),
    .S0(net1380),
    .S1(net1376),
    .X(_2157_));
 sky130_fd_sc_hd__a22o_1 _4157_ (.A1(net809),
    .A2(net1034),
    .B1(net1032),
    .B2(net722),
    .X(_2158_));
 sky130_fd_sc_hd__or2_1 _4158_ (.A(_2155_),
    .B(_2158_),
    .X(net248));
 sky130_fd_sc_hd__mux4_2 _4159_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][26] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][26] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][26] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][26] ),
    .S0(net1347),
    .S1(net1343),
    .X(_2159_));
 sky130_fd_sc_hd__a22o_1 _4160_ (.A1(net1286),
    .A2(net1161),
    .B1(net1031),
    .B2(net803),
    .X(_2160_));
 sky130_fd_sc_hd__mux4_2 _4161_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][26] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][26] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][26] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][26] ),
    .S0(net1318),
    .S1(net1313),
    .X(_2161_));
 sky130_fd_sc_hd__mux4_2 _4162_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][26] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][26] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][26] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][26] ),
    .S0(net1380),
    .S1(net1376),
    .X(_2162_));
 sky130_fd_sc_hd__a22o_1 _4163_ (.A1(net810),
    .A2(net1030),
    .B1(net1028),
    .B2(net721),
    .X(_2163_));
 sky130_fd_sc_hd__or2_1 _4164_ (.A(_2160_),
    .B(_2163_),
    .X(net249));
 sky130_fd_sc_hd__mux4_2 _4165_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][27] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][27] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][27] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][27] ),
    .S0(net1347),
    .S1(net1343),
    .X(_2164_));
 sky130_fd_sc_hd__a22o_1 _4166_ (.A1(net1285),
    .A2(net1161),
    .B1(net1027),
    .B2(net803),
    .X(_2165_));
 sky130_fd_sc_hd__mux4_2 _4167_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][27] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][27] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][27] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][27] ),
    .S0(net1319),
    .S1(net1314),
    .X(_2166_));
 sky130_fd_sc_hd__mux4_1 _4168_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][27] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][27] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][27] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][27] ),
    .S0(net1381),
    .S1(net1377),
    .X(_2167_));
 sky130_fd_sc_hd__a22o_1 _4169_ (.A1(net809),
    .A2(net1026),
    .B1(net1023),
    .B2(net721),
    .X(_2168_));
 sky130_fd_sc_hd__or2_1 _4170_ (.A(_2165_),
    .B(_2168_),
    .X(net250));
 sky130_fd_sc_hd__mux4_2 _4171_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][28] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][28] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][28] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][28] ),
    .S0(net1318),
    .S1(net1313),
    .X(_2169_));
 sky130_fd_sc_hd__a22o_1 _4172_ (.A1(net1284),
    .A2(net1158),
    .B1(net1022),
    .B2(net810),
    .X(_2170_));
 sky130_fd_sc_hd__mux4_2 _4173_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][28] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][28] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][28] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][28] ),
    .S0(net1381),
    .S1(net1377),
    .X(_2171_));
 sky130_fd_sc_hd__mux4_2 _4174_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][28] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][28] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][28] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][28] ),
    .S0(net1347),
    .S1(net1344),
    .X(_2172_));
 sky130_fd_sc_hd__a22o_1 _4175_ (.A1(net722),
    .A2(net1020),
    .B1(net1019),
    .B2(net804),
    .X(_2173_));
 sky130_fd_sc_hd__or2_1 _4176_ (.A(_2170_),
    .B(_2173_),
    .X(net251));
 sky130_fd_sc_hd__mux4_2 _4177_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][29] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][29] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][29] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][29] ),
    .S0(net1351),
    .S1(\u_s1.u_sync_wbb.u_resp_if.rd_ptr[1] ),
    .X(_2174_));
 sky130_fd_sc_hd__a22o_1 _4178_ (.A1(net1282),
    .A2(net1161),
    .B1(net1018),
    .B2(net803),
    .X(_2175_));
 sky130_fd_sc_hd__mux4_2 _4179_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][29] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][29] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][29] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][29] ),
    .S0(net1318),
    .S1(net1313),
    .X(_2176_));
 sky130_fd_sc_hd__mux4_2 _4180_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][29] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][29] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][29] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][29] ),
    .S0(net1380),
    .S1(net1376),
    .X(_2177_));
 sky130_fd_sc_hd__a22o_1 _4181_ (.A1(net809),
    .A2(net1017),
    .B1(net1015),
    .B2(net721),
    .X(_2178_));
 sky130_fd_sc_hd__or2_1 _4182_ (.A(_2175_),
    .B(_2178_),
    .X(net252));
 sky130_fd_sc_hd__mux4_2 _4183_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][30] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][30] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][30] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][30] ),
    .S0(net1347),
    .S1(net1343),
    .X(_2179_));
 sky130_fd_sc_hd__a22o_1 _4184_ (.A1(net1281),
    .A2(net1158),
    .B1(net1014),
    .B2(net804),
    .X(_2180_));
 sky130_fd_sc_hd__mux4_2 _4185_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][30] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][30] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][30] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][30] ),
    .S0(net1318),
    .S1(net1313),
    .X(_2181_));
 sky130_fd_sc_hd__mux4_2 _4186_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][30] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][30] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][30] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][30] ),
    .S0(net1380),
    .S1(net1376),
    .X(_2182_));
 sky130_fd_sc_hd__a22o_1 _4187_ (.A1(net810),
    .A2(net1013),
    .B1(net1011),
    .B2(net722),
    .X(_2183_));
 sky130_fd_sc_hd__or2_1 _4188_ (.A(_2180_),
    .B(_2183_),
    .X(net254));
 sky130_fd_sc_hd__mux4_1 _4189_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[0][31] ),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][31] ),
    .A2(\u_s0.u_sync_wbb.u_resp_if.mem[2][31] ),
    .A3(\u_s0.u_sync_wbb.u_resp_if.mem[3][31] ),
    .S0(net1321),
    .S1(net1316),
    .X(_2184_));
 sky130_fd_sc_hd__a22o_1 _4190_ (.A1(net1280),
    .A2(net1161),
    .B1(net1010),
    .B2(net809),
    .X(_2185_));
 sky130_fd_sc_hd__mux4_2 _4191_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[0][31] ),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][31] ),
    .A2(\u_s2.u_sync_wbb.u_resp_if.mem[2][31] ),
    .A3(\u_s2.u_sync_wbb.u_resp_if.mem[3][31] ),
    .S0(net1380),
    .S1(net1376),
    .X(_2186_));
 sky130_fd_sc_hd__mux4_2 _4192_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[0][31] ),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][31] ),
    .A2(\u_s1.u_sync_wbb.u_resp_if.mem[2][31] ),
    .A3(\u_s1.u_sync_wbb.u_resp_if.mem[3][31] ),
    .S0(net1348),
    .S1(net1343),
    .X(_2187_));
 sky130_fd_sc_hd__a22o_1 _4193_ (.A1(net721),
    .A2(net1008),
    .B1(net1007),
    .B2(net803),
    .X(_2188_));
 sky130_fd_sc_hd__or2_1 _4194_ (.A(_2185_),
    .B(_2188_),
    .X(net255));
 sky130_fd_sc_hd__and3b_2 _4195_ (.A_N(_1764_),
    .B(_1833_),
    .C(_1689_),
    .X(_2189_));
 sky130_fd_sc_hd__a22o_1 _4196_ (.A1(\u_reg.reg_ack ),
    .A2(net1164),
    .B1(net770),
    .B2(net1366),
    .X(_2190_));
 sky130_fd_sc_hd__a22o_1 _4197_ (.A1(\u_s0.u_sync_wbb.wbm_lack_o ),
    .A2(net735),
    .B1(net781),
    .B2(net1401),
    .X(_2191_));
 sky130_fd_sc_hd__or2_1 _4198_ (.A(_2190_),
    .B(_2191_),
    .X(net229));
 sky130_fd_sc_hd__a22o_1 _4199_ (.A1(\u_reg.reg_ack ),
    .A2(net1164),
    .B1(net770),
    .B2(net1367),
    .X(_2192_));
 sky130_fd_sc_hd__a22o_1 _4200_ (.A1(\u_s0.u_sync_wbb.wbm_ack_o ),
    .A2(net735),
    .B1(net781),
    .B2(net1402),
    .X(_2193_));
 sky130_fd_sc_hd__or2_1 _4201_ (.A(_2192_),
    .B(_2193_),
    .X(net196));
 sky130_fd_sc_hd__a22o_1 _4202_ (.A1(net1312),
    .A2(net1162),
    .B1(net1142),
    .B2(net733),
    .X(_2194_));
 sky130_fd_sc_hd__a22o_1 _4203_ (.A1(net779),
    .A2(net1140),
    .B1(net1138),
    .B2(net769),
    .X(_2195_));
 sky130_fd_sc_hd__or2_1 _4204_ (.A(_2194_),
    .B(_2195_),
    .X(net197));
 sky130_fd_sc_hd__a22o_1 _4205_ (.A1(\u_reg.reg_rdata[1] ),
    .A2(net1164),
    .B1(_2036_),
    .B2(net735),
    .X(_2196_));
 sky130_fd_sc_hd__a22o_1 _4206_ (.A1(net781),
    .A2(net1135),
    .B1(net770),
    .B2(net1137),
    .X(_2197_));
 sky130_fd_sc_hd__or2_1 _4207_ (.A(_2196_),
    .B(_2197_),
    .X(net208));
 sky130_fd_sc_hd__a22o_1 _4208_ (.A1(\u_reg.reg_rdata[2] ),
    .A2(net1164),
    .B1(net1129),
    .B2(net770),
    .X(_2198_));
 sky130_fd_sc_hd__a22o_1 _4209_ (.A1(net735),
    .A2(net1134),
    .B1(net1131),
    .B2(net781),
    .X(_2199_));
 sky130_fd_sc_hd__or2_1 _4210_ (.A(_2198_),
    .B(_2199_),
    .X(net219));
 sky130_fd_sc_hd__a22o_1 _4211_ (.A1(\u_reg.reg_rdata[3] ),
    .A2(net1164),
    .B1(net1128),
    .B2(net770),
    .X(_2200_));
 sky130_fd_sc_hd__a22o_1 _4212_ (.A1(net735),
    .A2(_2046_),
    .B1(net1126),
    .B2(net781),
    .X(_2201_));
 sky130_fd_sc_hd__or2_1 _4213_ (.A(_2200_),
    .B(_2201_),
    .X(net222));
 sky130_fd_sc_hd__a22o_1 _4214_ (.A1(net1311),
    .A2(net1164),
    .B1(net1122),
    .B2(net770),
    .X(_2202_));
 sky130_fd_sc_hd__a22o_1 _4215_ (.A1(net736),
    .A2(net1125),
    .B1(net1123),
    .B2(net782),
    .X(_2203_));
 sky130_fd_sc_hd__or2_1 _4216_ (.A(_2202_),
    .B(_2203_),
    .X(net223));
 sky130_fd_sc_hd__a22o_1 _4217_ (.A1(net1310),
    .A2(net1165),
    .B1(net1119),
    .B2(net736),
    .X(_2204_));
 sky130_fd_sc_hd__a22o_1 _4218_ (.A1(net782),
    .A2(net1116),
    .B1(net770),
    .B2(net1120),
    .X(_2205_));
 sky130_fd_sc_hd__or2_1 _4219_ (.A(_2204_),
    .B(_2205_),
    .X(net224));
 sky130_fd_sc_hd__a22o_1 _4220_ (.A1(\u_reg.reg_rdata[6] ),
    .A2(net1165),
    .B1(net1114),
    .B2(net736),
    .X(_2206_));
 sky130_fd_sc_hd__a22o_1 _4221_ (.A1(net782),
    .A2(net1112),
    .B1(net771),
    .B2(net1115),
    .X(_2207_));
 sky130_fd_sc_hd__or2_1 _4222_ (.A(_2206_),
    .B(_2207_),
    .X(net225));
 sky130_fd_sc_hd__a22o_1 _4223_ (.A1(net1309),
    .A2(net1163),
    .B1(net1111),
    .B2(net734),
    .X(_2208_));
 sky130_fd_sc_hd__a22o_1 _4224_ (.A1(net779),
    .A2(net1109),
    .B1(net1108),
    .B2(net769),
    .X(_2209_));
 sky130_fd_sc_hd__or2_1 _4225_ (.A(_2208_),
    .B(_2209_),
    .X(net226));
 sky130_fd_sc_hd__a22o_1 _4226_ (.A1(net1308),
    .A2(net1162),
    .B1(net1106),
    .B2(net769),
    .X(_2210_));
 sky130_fd_sc_hd__a22o_1 _4227_ (.A1(net735),
    .A2(_2071_),
    .B1(net1103),
    .B2(net781),
    .X(_2211_));
 sky130_fd_sc_hd__or2_1 _4228_ (.A(_2210_),
    .B(_2211_),
    .X(net227));
 sky130_fd_sc_hd__a22o_1 _4229_ (.A1(net1307),
    .A2(net1163),
    .B1(_2076_),
    .B2(net733),
    .X(_2212_));
 sky130_fd_sc_hd__a22o_1 _4230_ (.A1(net780),
    .A2(net1099),
    .B1(net769),
    .B2(net1102),
    .X(_2213_));
 sky130_fd_sc_hd__or2_1 _4231_ (.A(_2212_),
    .B(_2213_),
    .X(net228));
 sky130_fd_sc_hd__a22o_1 _4232_ (.A1(net1306),
    .A2(net1162),
    .B1(net1098),
    .B2(net769),
    .X(_2214_));
 sky130_fd_sc_hd__a22o_1 _4233_ (.A1(net733),
    .A2(_2081_),
    .B1(net1094),
    .B2(net779),
    .X(_2215_));
 sky130_fd_sc_hd__or2_1 _4234_ (.A(_2214_),
    .B(_2215_),
    .X(net198));
 sky130_fd_sc_hd__a22o_1 _4235_ (.A1(net1305),
    .A2(net1164),
    .B1(net1093),
    .B2(net735),
    .X(_2216_));
 sky130_fd_sc_hd__a22o_1 _4236_ (.A1(net781),
    .A2(net1092),
    .B1(net1091),
    .B2(net770),
    .X(_2217_));
 sky130_fd_sc_hd__or2_1 _4237_ (.A(_2216_),
    .B(_2217_),
    .X(net199));
 sky130_fd_sc_hd__a22o_1 _4238_ (.A1(net1304),
    .A2(net1162),
    .B1(net1090),
    .B2(net768),
    .X(_2218_));
 sky130_fd_sc_hd__a22o_1 _4239_ (.A1(net733),
    .A2(_2091_),
    .B1(net1086),
    .B2(net779),
    .X(_2219_));
 sky130_fd_sc_hd__or2_1 _4240_ (.A(_2218_),
    .B(_2219_),
    .X(net200));
 sky130_fd_sc_hd__a22o_1 _4241_ (.A1(net1302),
    .A2(net1164),
    .B1(net1085),
    .B2(net770),
    .X(_2220_));
 sky130_fd_sc_hd__a22o_1 _4242_ (.A1(net735),
    .A2(net1084),
    .B1(net1082),
    .B2(net781),
    .X(_2221_));
 sky130_fd_sc_hd__or2_1 _4243_ (.A(_2220_),
    .B(_2221_),
    .X(net201));
 sky130_fd_sc_hd__a22o_1 _4244_ (.A1(net1300),
    .A2(net1163),
    .B1(net1081),
    .B2(net768),
    .X(_2222_));
 sky130_fd_sc_hd__a22o_1 _4245_ (.A1(net733),
    .A2(_2101_),
    .B1(net1078),
    .B2(net779),
    .X(_2223_));
 sky130_fd_sc_hd__or2_1 _4246_ (.A(_2222_),
    .B(_2223_),
    .X(net202));
 sky130_fd_sc_hd__a22o_1 _4247_ (.A1(net1298),
    .A2(net1165),
    .B1(net1073),
    .B2(net771),
    .X(_2224_));
 sky130_fd_sc_hd__a22o_1 _4248_ (.A1(net736),
    .A2(net1077),
    .B1(net1075),
    .B2(net782),
    .X(_2225_));
 sky130_fd_sc_hd__or2_1 _4249_ (.A(_2224_),
    .B(_2225_),
    .X(net203));
 sky130_fd_sc_hd__a22o_1 _4250_ (.A1(net1296),
    .A2(net1163),
    .B1(net1071),
    .B2(net768),
    .X(_2226_));
 sky130_fd_sc_hd__a22o_1 _4251_ (.A1(net734),
    .A2(net1070),
    .B1(net1068),
    .B2(net780),
    .X(_2227_));
 sky130_fd_sc_hd__or2_1 _4252_ (.A(_2226_),
    .B(_2227_),
    .X(net204));
 sky130_fd_sc_hd__a22o_1 _4253_ (.A1(net1295),
    .A2(net1165),
    .B1(net1067),
    .B2(net771),
    .X(_2228_));
 sky130_fd_sc_hd__a22o_1 _4254_ (.A1(net735),
    .A2(net1066),
    .B1(net1064),
    .B2(net782),
    .X(_2229_));
 sky130_fd_sc_hd__or2_1 _4255_ (.A(_2228_),
    .B(_2229_),
    .X(net205));
 sky130_fd_sc_hd__a22o_1 _4256_ (.A1(\u_reg.reg_rdata[18] ),
    .A2(net1162),
    .B1(net1063),
    .B2(net733),
    .X(_2230_));
 sky130_fd_sc_hd__a22o_1 _4257_ (.A1(net779),
    .A2(net1060),
    .B1(net1058),
    .B2(net768),
    .X(_2231_));
 sky130_fd_sc_hd__or2_1 _4258_ (.A(_2230_),
    .B(_2231_),
    .X(net206));
 sky130_fd_sc_hd__a22o_1 _4259_ (.A1(\u_reg.reg_rdata[19] ),
    .A2(net1164),
    .B1(_2126_),
    .B2(net736),
    .X(_2232_));
 sky130_fd_sc_hd__a22o_1 _4260_ (.A1(net781),
    .A2(net1056),
    .B1(net771),
    .B2(net1057),
    .X(_2233_));
 sky130_fd_sc_hd__or2_1 _4261_ (.A(_2232_),
    .B(_2233_),
    .X(net207));
 sky130_fd_sc_hd__a22o_1 _4262_ (.A1(net1293),
    .A2(net1162),
    .B1(net1055),
    .B2(net769),
    .X(_2234_));
 sky130_fd_sc_hd__a22o_1 _4263_ (.A1(net734),
    .A2(net1054),
    .B1(net1051),
    .B2(net780),
    .X(_2235_));
 sky130_fd_sc_hd__or2_1 _4264_ (.A(_2234_),
    .B(_2235_),
    .X(net209));
 sky130_fd_sc_hd__a22o_1 _4265_ (.A1(net1291),
    .A2(net1162),
    .B1(net1050),
    .B2(net735),
    .X(_2236_));
 sky130_fd_sc_hd__a22o_1 _4266_ (.A1(net781),
    .A2(net1048),
    .B1(net1047),
    .B2(net770),
    .X(_2237_));
 sky130_fd_sc_hd__or2_1 _4267_ (.A(_2236_),
    .B(_2237_),
    .X(net210));
 sky130_fd_sc_hd__a22o_1 _4268_ (.A1(net1290),
    .A2(net1163),
    .B1(net1046),
    .B2(net734),
    .X(_2238_));
 sky130_fd_sc_hd__a22o_1 _4269_ (.A1(net780),
    .A2(net1044),
    .B1(net1043),
    .B2(net768),
    .X(_2239_));
 sky130_fd_sc_hd__or2_1 _4270_ (.A(_2238_),
    .B(_2239_),
    .X(net211));
 sky130_fd_sc_hd__a22o_1 _4271_ (.A1(\u_reg.reg_rdata[23] ),
    .A2(net1162),
    .B1(net1039),
    .B2(net768),
    .X(_2240_));
 sky130_fd_sc_hd__a22o_1 _4272_ (.A1(net733),
    .A2(_2144_),
    .B1(net1040),
    .B2(net779),
    .X(_2241_));
 sky130_fd_sc_hd__or2_1 _4273_ (.A(_2240_),
    .B(_2241_),
    .X(net212));
 sky130_fd_sc_hd__a22o_1 _4274_ (.A1(net1289),
    .A2(net1165),
    .B1(net1036),
    .B2(net771),
    .X(_2242_));
 sky130_fd_sc_hd__a22o_1 _4275_ (.A1(net736),
    .A2(net1038),
    .B1(net1037),
    .B2(net782),
    .X(_2243_));
 sky130_fd_sc_hd__or2_1 _4276_ (.A(_2242_),
    .B(_2243_),
    .X(net213));
 sky130_fd_sc_hd__a22o_1 _4277_ (.A1(net1288),
    .A2(net1165),
    .B1(net1034),
    .B2(net736),
    .X(_2244_));
 sky130_fd_sc_hd__a22o_1 _4278_ (.A1(net782),
    .A2(net1032),
    .B1(net771),
    .B2(net1035),
    .X(_2245_));
 sky130_fd_sc_hd__or2_1 _4279_ (.A(_2244_),
    .B(_2245_),
    .X(net214));
 sky130_fd_sc_hd__a22o_1 _4280_ (.A1(net1286),
    .A2(net1162),
    .B1(net1031),
    .B2(net769),
    .X(_2246_));
 sky130_fd_sc_hd__a22o_1 _4281_ (.A1(net733),
    .A2(net1030),
    .B1(net1028),
    .B2(net779),
    .X(_2247_));
 sky130_fd_sc_hd__or2_1 _4282_ (.A(_2246_),
    .B(_2247_),
    .X(net215));
 sky130_fd_sc_hd__a22o_1 _4283_ (.A1(net1285),
    .A2(net1163),
    .B1(net1026),
    .B2(net734),
    .X(_2248_));
 sky130_fd_sc_hd__a22o_1 _4284_ (.A1(net780),
    .A2(net1023),
    .B1(net768),
    .B2(net1027),
    .X(_2249_));
 sky130_fd_sc_hd__or2_1 _4285_ (.A(_2248_),
    .B(_2249_),
    .X(net216));
 sky130_fd_sc_hd__a22o_1 _4286_ (.A1(net1284),
    .A2(net1163),
    .B1(net1019),
    .B2(net768),
    .X(_2250_));
 sky130_fd_sc_hd__a22o_1 _4287_ (.A1(net733),
    .A2(net1022),
    .B1(net1020),
    .B2(net779),
    .X(_2251_));
 sky130_fd_sc_hd__or2_1 _4288_ (.A(_2250_),
    .B(_2251_),
    .X(net217));
 sky130_fd_sc_hd__a22o_1 _4289_ (.A1(net1282),
    .A2(net1163),
    .B1(net1018),
    .B2(net768),
    .X(_2252_));
 sky130_fd_sc_hd__a22o_1 _4290_ (.A1(net734),
    .A2(net1017),
    .B1(net1015),
    .B2(net780),
    .X(_2253_));
 sky130_fd_sc_hd__or2_1 _4291_ (.A(_2252_),
    .B(_2253_),
    .X(net218));
 sky130_fd_sc_hd__a22o_1 _4292_ (.A1(net1281),
    .A2(net1163),
    .B1(net1014),
    .B2(net768),
    .X(_2254_));
 sky130_fd_sc_hd__a22o_1 _4293_ (.A1(net734),
    .A2(net1013),
    .B1(net1011),
    .B2(net780),
    .X(_2255_));
 sky130_fd_sc_hd__or2_1 _4294_ (.A(_2254_),
    .B(_2255_),
    .X(net220));
 sky130_fd_sc_hd__a22o_1 _4295_ (.A1(net1280),
    .A2(net1162),
    .B1(net1007),
    .B2(net769),
    .X(_2256_));
 sky130_fd_sc_hd__a22o_1 _4296_ (.A1(net733),
    .A2(net1010),
    .B1(net1008),
    .B2(net779),
    .X(_2257_));
 sky130_fd_sc_hd__or2_1 _4297_ (.A(_2256_),
    .B(_2257_),
    .X(net221));
 sky130_fd_sc_hd__a22o_1 _4298_ (.A1(net1366),
    .A2(net801),
    .B1(net1147),
    .B2(\u_reg.reg_ack ),
    .X(_2258_));
 sky130_fd_sc_hd__and4bb_4 _4299_ (.A_N(_1684_),
    .B_N(_1752_),
    .C(net1173),
    .D(_1685_),
    .X(_2259_));
 sky130_fd_sc_hd__a22o_1 _4300_ (.A1(\u_s0.u_sync_wbb.wbm_lack_o ),
    .A2(net815),
    .B1(net766),
    .B2(net1401),
    .X(_2260_));
 sky130_fd_sc_hd__or2_4 _4301_ (.A(_2258_),
    .B(_2260_),
    .X(net195));
 sky130_fd_sc_hd__a22o_1 _4302_ (.A1(net1367),
    .A2(net802),
    .B1(net1145),
    .B2(\u_reg.reg_ack ),
    .X(_2261_));
 sky130_fd_sc_hd__a22o_1 _4303_ (.A1(\u_s0.u_sync_wbb.wbm_ack_o ),
    .A2(net815),
    .B1(net766),
    .B2(net1402),
    .X(_2262_));
 sky130_fd_sc_hd__or2_4 _4304_ (.A(_2261_),
    .B(_2262_),
    .X(net162));
 sky130_fd_sc_hd__a22o_1 _4305_ (.A1(net1312),
    .A2(net1143),
    .B1(net1142),
    .B2(net813),
    .X(_2263_));
 sky130_fd_sc_hd__a22o_1 _4306_ (.A1(net799),
    .A2(net1138),
    .B1(net764),
    .B2(net1140),
    .X(_2264_));
 sky130_fd_sc_hd__or2_4 _4307_ (.A(_2263_),
    .B(_2264_),
    .X(net163));
 sky130_fd_sc_hd__a22o_1 _4308_ (.A1(\u_reg.reg_rdata[1] ),
    .A2(net1145),
    .B1(net1137),
    .B2(net801),
    .X(_2265_));
 sky130_fd_sc_hd__a22o_1 _4309_ (.A1(net815),
    .A2(_2036_),
    .B1(net1135),
    .B2(net766),
    .X(_2266_));
 sky130_fd_sc_hd__or2_4 _4310_ (.A(_2265_),
    .B(_2266_),
    .X(net174));
 sky130_fd_sc_hd__a22o_1 _4311_ (.A1(\u_reg.reg_rdata[2] ),
    .A2(net1143),
    .B1(net1134),
    .B2(net813),
    .X(_2267_));
 sky130_fd_sc_hd__a22o_1 _4312_ (.A1(net799),
    .A2(net1129),
    .B1(net764),
    .B2(net1131),
    .X(_2268_));
 sky130_fd_sc_hd__or2_4 _4313_ (.A(_2267_),
    .B(_2268_),
    .X(net185));
 sky130_fd_sc_hd__a22o_1 _4314_ (.A1(\u_reg.reg_rdata[3] ),
    .A2(net1145),
    .B1(net1128),
    .B2(net801),
    .X(_2269_));
 sky130_fd_sc_hd__a22o_1 _4315_ (.A1(net815),
    .A2(_2046_),
    .B1(net1126),
    .B2(net766),
    .X(_2270_));
 sky130_fd_sc_hd__or2_4 _4316_ (.A(_2269_),
    .B(_2270_),
    .X(net188));
 sky130_fd_sc_hd__a22o_1 _4317_ (.A1(net1311),
    .A2(net1146),
    .B1(net1125),
    .B2(net816),
    .X(_2271_));
 sky130_fd_sc_hd__a22o_1 _4318_ (.A1(net802),
    .A2(net1122),
    .B1(net767),
    .B2(net1123),
    .X(_2272_));
 sky130_fd_sc_hd__or2_4 _4319_ (.A(_2271_),
    .B(_2272_),
    .X(net189));
 sky130_fd_sc_hd__a22o_1 _4320_ (.A1(net1310),
    .A2(net1145),
    .B1(net1119),
    .B2(net815),
    .X(_2273_));
 sky130_fd_sc_hd__a22o_1 _4321_ (.A1(net801),
    .A2(net1120),
    .B1(net1116),
    .B2(net766),
    .X(_2274_));
 sky130_fd_sc_hd__or2_4 _4322_ (.A(_2273_),
    .B(_2274_),
    .X(net190));
 sky130_fd_sc_hd__a22o_1 _4323_ (.A1(\u_reg.reg_rdata[6] ),
    .A2(net1145),
    .B1(net1115),
    .B2(net802),
    .X(_2275_));
 sky130_fd_sc_hd__a22o_1 _4324_ (.A1(net816),
    .A2(net1114),
    .B1(net1112),
    .B2(net767),
    .X(_2276_));
 sky130_fd_sc_hd__or2_4 _4325_ (.A(_2275_),
    .B(_2276_),
    .X(net191));
 sky130_fd_sc_hd__a22o_1 _4326_ (.A1(net1309),
    .A2(net1143),
    .B1(net1108),
    .B2(net799),
    .X(_2277_));
 sky130_fd_sc_hd__a22o_1 _4327_ (.A1(net814),
    .A2(net1111),
    .B1(net1109),
    .B2(net764),
    .X(_2278_));
 sky130_fd_sc_hd__or2_2 _4328_ (.A(_2277_),
    .B(_2278_),
    .X(net192));
 sky130_fd_sc_hd__a22o_1 _4329_ (.A1(net1308),
    .A2(net1145),
    .B1(_2071_),
    .B2(net815),
    .X(_2279_));
 sky130_fd_sc_hd__a22o_1 _4330_ (.A1(net801),
    .A2(net1106),
    .B1(net1103),
    .B2(net766),
    .X(_2280_));
 sky130_fd_sc_hd__or2_4 _4331_ (.A(_2279_),
    .B(_2280_),
    .X(net193));
 sky130_fd_sc_hd__a22o_1 _4332_ (.A1(net1307),
    .A2(net1143),
    .B1(net1102),
    .B2(net799),
    .X(_2281_));
 sky130_fd_sc_hd__a22o_1 _4333_ (.A1(net813),
    .A2(_2076_),
    .B1(net1099),
    .B2(net764),
    .X(_2282_));
 sky130_fd_sc_hd__or2_4 _4334_ (.A(_2281_),
    .B(_2282_),
    .X(net194));
 sky130_fd_sc_hd__a22o_1 _4335_ (.A1(net1306),
    .A2(net1143),
    .B1(_2081_),
    .B2(net813),
    .X(_2283_));
 sky130_fd_sc_hd__a22o_1 _4336_ (.A1(net799),
    .A2(net1098),
    .B1(net1094),
    .B2(net764),
    .X(_2284_));
 sky130_fd_sc_hd__or2_4 _4337_ (.A(_2283_),
    .B(_2284_),
    .X(net164));
 sky130_fd_sc_hd__a22o_1 _4338_ (.A1(net1305),
    .A2(net1146),
    .B1(net1091),
    .B2(net802),
    .X(_2285_));
 sky130_fd_sc_hd__a22o_1 _4339_ (.A1(net815),
    .A2(net1093),
    .B1(net1092),
    .B2(net766),
    .X(_2286_));
 sky130_fd_sc_hd__or2_4 _4340_ (.A(_2285_),
    .B(_2286_),
    .X(net165));
 sky130_fd_sc_hd__a22o_1 _4341_ (.A1(net1304),
    .A2(net1143),
    .B1(_2091_),
    .B2(net813),
    .X(_2287_));
 sky130_fd_sc_hd__a22o_1 _4342_ (.A1(net799),
    .A2(net1090),
    .B1(net1086),
    .B2(net764),
    .X(_2288_));
 sky130_fd_sc_hd__or2_4 _4343_ (.A(_2287_),
    .B(_2288_),
    .X(net166));
 sky130_fd_sc_hd__a22o_1 _4344_ (.A1(net1302),
    .A2(net1145),
    .B1(net1085),
    .B2(net801),
    .X(_2289_));
 sky130_fd_sc_hd__a22o_1 _4345_ (.A1(net815),
    .A2(_2096_),
    .B1(net1082),
    .B2(net766),
    .X(_2290_));
 sky130_fd_sc_hd__or2_4 _4346_ (.A(_2289_),
    .B(_2290_),
    .X(net167));
 sky130_fd_sc_hd__a22o_1 _4347_ (.A1(net1300),
    .A2(net1144),
    .B1(net1081),
    .B2(net800),
    .X(_2291_));
 sky130_fd_sc_hd__a22o_1 _4348_ (.A1(net814),
    .A2(_2101_),
    .B1(net1078),
    .B2(net765),
    .X(_2292_));
 sky130_fd_sc_hd__or2_2 _4349_ (.A(_2291_),
    .B(_2292_),
    .X(net168));
 sky130_fd_sc_hd__a22o_1 _4350_ (.A1(net1298),
    .A2(net1146),
    .B1(net1073),
    .B2(net802),
    .X(_2293_));
 sky130_fd_sc_hd__a22o_1 _4351_ (.A1(net816),
    .A2(_2104_),
    .B1(net1075),
    .B2(net767),
    .X(_2294_));
 sky130_fd_sc_hd__or2_4 _4352_ (.A(_2293_),
    .B(_2294_),
    .X(net169));
 sky130_fd_sc_hd__a22o_1 _4353_ (.A1(net1296),
    .A2(net1144),
    .B1(_2111_),
    .B2(net1777),
    .X(_2295_));
 sky130_fd_sc_hd__a22o_1 _4354_ (.A1(net800),
    .A2(net1071),
    .B1(net1068),
    .B2(net765),
    .X(_2296_));
 sky130_fd_sc_hd__or2_4 _4355_ (.A(_2295_),
    .B(_2296_),
    .X(net170));
 sky130_fd_sc_hd__a22o_1 _4356_ (.A1(net1295),
    .A2(net1145),
    .B1(net1066),
    .B2(net816),
    .X(_2297_));
 sky130_fd_sc_hd__a22o_1 _4357_ (.A1(net801),
    .A2(net1067),
    .B1(net1064),
    .B2(net766),
    .X(_2298_));
 sky130_fd_sc_hd__or2_4 _4358_ (.A(_2297_),
    .B(_2298_),
    .X(net171));
 sky130_fd_sc_hd__a22o_1 _4359_ (.A1(\u_reg.reg_rdata[18] ),
    .A2(net1144),
    .B1(net1058),
    .B2(net800),
    .X(_2299_));
 sky130_fd_sc_hd__a22o_1 _4360_ (.A1(net814),
    .A2(net1063),
    .B1(net1060),
    .B2(net765),
    .X(_2300_));
 sky130_fd_sc_hd__or2_1 _4361_ (.A(_2299_),
    .B(_2300_),
    .X(net172));
 sky130_fd_sc_hd__a22o_1 _4362_ (.A1(\u_reg.reg_rdata[19] ),
    .A2(net1146),
    .B1(net1057),
    .B2(net802),
    .X(_2301_));
 sky130_fd_sc_hd__a22o_1 _4363_ (.A1(net816),
    .A2(_2126_),
    .B1(net1056),
    .B2(net767),
    .X(_2302_));
 sky130_fd_sc_hd__or2_4 _4364_ (.A(_2301_),
    .B(_2302_),
    .X(net173));
 sky130_fd_sc_hd__a22o_1 _4365_ (.A1(net1293),
    .A2(net1143),
    .B1(_2131_),
    .B2(net813),
    .X(_2303_));
 sky130_fd_sc_hd__a22o_1 _4366_ (.A1(net799),
    .A2(net1055),
    .B1(net1051),
    .B2(net764),
    .X(_2304_));
 sky130_fd_sc_hd__or2_4 _4367_ (.A(_2303_),
    .B(_2304_),
    .X(net175));
 sky130_fd_sc_hd__a22o_1 _4368_ (.A1(net1291),
    .A2(net1145),
    .B1(net1050),
    .B2(net815),
    .X(_2305_));
 sky130_fd_sc_hd__a22o_1 _4369_ (.A1(net801),
    .A2(net1047),
    .B1(net766),
    .B2(net1048),
    .X(_2306_));
 sky130_fd_sc_hd__or2_4 _4370_ (.A(_2305_),
    .B(_2306_),
    .X(net176));
 sky130_fd_sc_hd__a22o_1 _4371_ (.A1(net1290),
    .A2(net1144),
    .B1(_2139_),
    .B2(net814),
    .X(_2307_));
 sky130_fd_sc_hd__a22o_1 _4372_ (.A1(net800),
    .A2(net1043),
    .B1(net765),
    .B2(net1044),
    .X(_2308_));
 sky130_fd_sc_hd__or2_1 _4373_ (.A(_2307_),
    .B(_2308_),
    .X(net177));
 sky130_fd_sc_hd__a22o_1 _4374_ (.A1(\u_reg.reg_rdata[23] ),
    .A2(net1143),
    .B1(net1039),
    .B2(net799),
    .X(_2309_));
 sky130_fd_sc_hd__a22o_1 _4375_ (.A1(net813),
    .A2(_2144_),
    .B1(net1040),
    .B2(net764),
    .X(_2310_));
 sky130_fd_sc_hd__or2_4 _4376_ (.A(_2309_),
    .B(_2310_),
    .X(net178));
 sky130_fd_sc_hd__a22o_1 _4377_ (.A1(net1289),
    .A2(net1145),
    .B1(net1038),
    .B2(net816),
    .X(_2311_));
 sky130_fd_sc_hd__a22o_1 _4378_ (.A1(net801),
    .A2(net1036),
    .B1(net767),
    .B2(net1037),
    .X(_2312_));
 sky130_fd_sc_hd__or2_4 _4379_ (.A(_2311_),
    .B(_2312_),
    .X(net179));
 sky130_fd_sc_hd__a22o_1 _4380_ (.A1(net1288),
    .A2(net1146),
    .B1(_2156_),
    .B2(net815),
    .X(_2313_));
 sky130_fd_sc_hd__a22o_1 _4381_ (.A1(net801),
    .A2(net1035),
    .B1(net1032),
    .B2(net767),
    .X(_2314_));
 sky130_fd_sc_hd__or2_4 _4382_ (.A(_2313_),
    .B(_2314_),
    .X(net180));
 sky130_fd_sc_hd__a22o_1 _4383_ (.A1(net1286),
    .A2(net1143),
    .B1(_2161_),
    .B2(net813),
    .X(_2315_));
 sky130_fd_sc_hd__a22o_1 _4384_ (.A1(net799),
    .A2(net1031),
    .B1(net1028),
    .B2(net764),
    .X(_2316_));
 sky130_fd_sc_hd__or2_4 _4385_ (.A(_2315_),
    .B(_2316_),
    .X(net181));
 sky130_fd_sc_hd__a22o_1 _4386_ (.A1(net1285),
    .A2(net1144),
    .B1(net1027),
    .B2(net800),
    .X(_2317_));
 sky130_fd_sc_hd__a22o_1 _4387_ (.A1(net1777),
    .A2(_2166_),
    .B1(net1023),
    .B2(net765),
    .X(_2318_));
 sky130_fd_sc_hd__or2_4 _4388_ (.A(_2317_),
    .B(_2318_),
    .X(net182));
 sky130_fd_sc_hd__a22o_1 _4389_ (.A1(net1284),
    .A2(net1143),
    .B1(_2169_),
    .B2(net813),
    .X(_2319_));
 sky130_fd_sc_hd__a22o_1 _4390_ (.A1(net799),
    .A2(net1019),
    .B1(net764),
    .B2(net1020),
    .X(_2320_));
 sky130_fd_sc_hd__or2_4 _4391_ (.A(_2319_),
    .B(_2320_),
    .X(net183));
 sky130_fd_sc_hd__a22o_1 _4392_ (.A1(net1282),
    .A2(net1144),
    .B1(net1018),
    .B2(net800),
    .X(_2321_));
 sky130_fd_sc_hd__a22o_1 _4393_ (.A1(net1777),
    .A2(_2176_),
    .B1(net1015),
    .B2(net765),
    .X(_2322_));
 sky130_fd_sc_hd__or2_4 _4394_ (.A(_2321_),
    .B(_2322_),
    .X(net184));
 sky130_fd_sc_hd__a22o_1 _4395_ (.A1(net1281),
    .A2(net1144),
    .B1(net1014),
    .B2(net800),
    .X(_2323_));
 sky130_fd_sc_hd__a22o_1 _4396_ (.A1(net1777),
    .A2(_2181_),
    .B1(net1011),
    .B2(net765),
    .X(_2324_));
 sky130_fd_sc_hd__or2_4 _4397_ (.A(_2323_),
    .B(_2324_),
    .X(net186));
 sky130_fd_sc_hd__a22o_1 _4398_ (.A1(net1280),
    .A2(net1144),
    .B1(net1007),
    .B2(net800),
    .X(_2325_));
 sky130_fd_sc_hd__a22o_1 _4399_ (.A1(net813),
    .A2(net1010),
    .B1(net1008),
    .B2(net765),
    .X(_2326_));
 sky130_fd_sc_hd__or2_4 _4400_ (.A(_2325_),
    .B(_2326_),
    .X(net187));
 sky130_fd_sc_hd__a31o_1 _4401_ (.A1(\u_dcg_s0.cfg_mode_ss[0] ),
    .A2(\u_dcg_s0.dst_idle_r ),
    .A3(net737),
    .B1(\u_dcg_s0.cfg_mode_ss[1] ),
    .X(_2327_));
 sky130_fd_sc_hd__o21ai_1 _4402_ (.A1(\u_dcg_s0.cfg_mode_ss[1] ),
    .A2(\u_dcg_s0.idle_his ),
    .B1(\u_dcg_s0.cfg_mode_ss[0] ),
    .Y(_2328_));
 sky130_fd_sc_hd__nand2_2 _4403_ (.A(_2327_),
    .B(_2328_),
    .Y(\u_dcg_s0.clk_enb ));
 sky130_fd_sc_hd__mux4_2 _4404_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][14] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][14] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][14] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][14] ),
    .S0(net1397),
    .S1(net1390),
    .X(_2329_));
 sky130_fd_sc_hd__mux2_1 _4405_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[14] ),
    .A1(_2329_),
    .S(net714),
    .X(net471));
 sky130_fd_sc_hd__mux4_2 _4406_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][15] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][15] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][15] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][15] ),
    .S0(net1398),
    .S1(net1391),
    .X(_2330_));
 sky130_fd_sc_hd__mux2_2 _4407_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[15] ),
    .A1(_2330_),
    .S(net717),
    .X(net472));
 sky130_fd_sc_hd__mux4_2 _4408_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][16] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][16] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][16] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][16] ),
    .S0(net1396),
    .S1(net1389),
    .X(_2331_));
 sky130_fd_sc_hd__mux2_1 _4409_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[16] ),
    .A1(_2331_),
    .S(net716),
    .X(net473));
 sky130_fd_sc_hd__mux4_2 _4410_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][17] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][17] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][17] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][17] ),
    .S0(net1393),
    .S1(net1386),
    .X(_2332_));
 sky130_fd_sc_hd__mux2_1 _4411_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[17] ),
    .A1(_2332_),
    .S(net713),
    .X(net474));
 sky130_fd_sc_hd__mux4_2 _4412_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][18] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][18] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][18] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][18] ),
    .S0(net1394),
    .S1(net1388),
    .X(_2333_));
 sky130_fd_sc_hd__mux2_1 _4413_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[18] ),
    .A1(_2333_),
    .S(net716),
    .X(net439));
 sky130_fd_sc_hd__mux4_2 _4414_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][19] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][19] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][19] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][19] ),
    .S0(net1395),
    .S1(net1388),
    .X(_2334_));
 sky130_fd_sc_hd__mux2_4 _4415_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[19] ),
    .A1(_2334_),
    .S(net717),
    .X(net450));
 sky130_fd_sc_hd__mux4_2 _4416_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][20] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][20] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][20] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][20] ),
    .S0(net1397),
    .S1(net1390),
    .X(_2335_));
 sky130_fd_sc_hd__mux2_2 _4417_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[20] ),
    .A1(_2335_),
    .S(net716),
    .X(net461));
 sky130_fd_sc_hd__mux4_1 _4418_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][21] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][21] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][21] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][21] ),
    .S0(net1394),
    .S1(net1387),
    .X(_2336_));
 sky130_fd_sc_hd__mux2_1 _4419_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[21] ),
    .A1(_2336_),
    .S(net715),
    .X(net464));
 sky130_fd_sc_hd__mux4_2 _4420_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][22] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][22] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][22] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][22] ),
    .S0(net1397),
    .S1(net1390),
    .X(_2337_));
 sky130_fd_sc_hd__mux2_4 _4421_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[22] ),
    .A1(_2337_),
    .S(net717),
    .X(net465));
 sky130_fd_sc_hd__mux4_2 _4422_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][23] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][23] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][23] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][23] ),
    .S0(net1395),
    .S1(net1388),
    .X(_2338_));
 sky130_fd_sc_hd__mux2_2 _4423_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[23] ),
    .A1(_2338_),
    .S(net716),
    .X(net466));
 sky130_fd_sc_hd__mux4_2 _4424_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][24] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][24] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][24] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][24] ),
    .S0(net1395),
    .S1(net1387),
    .X(_2339_));
 sky130_fd_sc_hd__mux2_1 _4425_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[24] ),
    .A1(_2339_),
    .S(net714),
    .X(net467));
 sky130_fd_sc_hd__mux4_2 _4426_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][25] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][25] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][25] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][25] ),
    .S0(net1397),
    .S1(net1390),
    .X(_2340_));
 sky130_fd_sc_hd__mux2_2 _4427_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[25] ),
    .A1(_2340_),
    .S(net716),
    .X(net468));
 sky130_fd_sc_hd__mux4_2 _4428_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][26] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][26] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][26] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][26] ),
    .S0(net1393),
    .S1(net1386),
    .X(_2341_));
 sky130_fd_sc_hd__mux2_1 _4429_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[26] ),
    .A1(_2341_),
    .S(net715),
    .X(net469));
 sky130_fd_sc_hd__mux4_2 _4430_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][27] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][27] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][27] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][27] ),
    .S0(net1394),
    .S1(net1387),
    .X(_2342_));
 sky130_fd_sc_hd__mux2_1 _4431_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[27] ),
    .A1(_2342_),
    .S(net714),
    .X(net470));
 sky130_fd_sc_hd__mux4_2 _4432_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][28] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][28] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][28] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][28] ),
    .S0(net1397),
    .S1(net1390),
    .X(_2343_));
 sky130_fd_sc_hd__mux2_4 _4433_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[28] ),
    .A1(_2343_),
    .S(net717),
    .X(net440));
 sky130_fd_sc_hd__mux4_2 _4434_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][29] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][29] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][29] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][29] ),
    .S0(net1393),
    .S1(net1386),
    .X(_2344_));
 sky130_fd_sc_hd__mux2_1 _4435_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[29] ),
    .A1(_2344_),
    .S(net714),
    .X(net441));
 sky130_fd_sc_hd__mux4_2 _4436_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][30] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][30] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][30] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][30] ),
    .S0(net1394),
    .S1(net1387),
    .X(_2345_));
 sky130_fd_sc_hd__mux2_1 _4437_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[30] ),
    .A1(_2345_),
    .S(net715),
    .X(net442));
 sky130_fd_sc_hd__mux4_2 _4438_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][31] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][31] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][31] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][31] ),
    .S0(net1392),
    .S1(net1385),
    .X(_2346_));
 sky130_fd_sc_hd__mux2_2 _4439_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[31] ),
    .A1(_2346_),
    .S(net713),
    .X(net443));
 sky130_fd_sc_hd__mux4_2 _4440_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][32] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][32] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][32] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][32] ),
    .S0(net1396),
    .S1(net1389),
    .X(_2347_));
 sky130_fd_sc_hd__mux2_1 _4441_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[32] ),
    .A1(_2347_),
    .S(net714),
    .X(net444));
 sky130_fd_sc_hd__mux4_2 _4442_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][33] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][33] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][33] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][33] ),
    .S0(net1396),
    .S1(net1389),
    .X(_2348_));
 sky130_fd_sc_hd__mux2_1 _4443_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[33] ),
    .A1(_2348_),
    .S(net716),
    .X(net445));
 sky130_fd_sc_hd__mux4_2 _4444_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][34] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][34] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][34] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][34] ),
    .S0(net1396),
    .S1(net1389),
    .X(_2349_));
 sky130_fd_sc_hd__mux2_1 _4445_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[34] ),
    .A1(_2349_),
    .S(net716),
    .X(net446));
 sky130_fd_sc_hd__mux4_2 _4446_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][35] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][35] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][35] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][35] ),
    .S0(net1396),
    .S1(net1389),
    .X(_2350_));
 sky130_fd_sc_hd__mux2_1 _4447_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[35] ),
    .A1(_2350_),
    .S(net717),
    .X(net447));
 sky130_fd_sc_hd__mux4_2 _4448_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][36] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][36] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][36] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][36] ),
    .S0(net1397),
    .S1(net1390),
    .X(_2351_));
 sky130_fd_sc_hd__mux2_2 _4449_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[36] ),
    .A1(_2351_),
    .S(net717),
    .X(net448));
 sky130_fd_sc_hd__mux4_2 _4450_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][37] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][37] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][37] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][37] ),
    .S0(net1397),
    .S1(net1390),
    .X(_2352_));
 sky130_fd_sc_hd__mux2_1 _4451_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[37] ),
    .A1(_2352_),
    .S(net714),
    .X(net449));
 sky130_fd_sc_hd__mux4_2 _4452_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][38] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][38] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][38] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][38] ),
    .S0(net1392),
    .S1(net1385),
    .X(_2353_));
 sky130_fd_sc_hd__mux2_1 _4453_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[38] ),
    .A1(_2353_),
    .S(net714),
    .X(net451));
 sky130_fd_sc_hd__mux4_2 _4454_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][39] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][39] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][39] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][39] ),
    .S0(net1392),
    .S1(net1385),
    .X(_2354_));
 sky130_fd_sc_hd__mux2_2 _4455_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[39] ),
    .A1(_2354_),
    .S(net713),
    .X(net452));
 sky130_fd_sc_hd__mux4_2 _4456_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][40] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][40] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][40] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][40] ),
    .S0(net1393),
    .S1(net1386),
    .X(_2355_));
 sky130_fd_sc_hd__mux2_1 _4457_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[40] ),
    .A1(_2355_),
    .S(net718),
    .X(net453));
 sky130_fd_sc_hd__mux4_2 _4458_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][41] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][41] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][41] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][41] ),
    .S0(net1392),
    .S1(net1385),
    .X(_2356_));
 sky130_fd_sc_hd__mux2_1 _4459_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[41] ),
    .A1(_2356_),
    .S(net714),
    .X(net454));
 sky130_fd_sc_hd__mux4_2 _4460_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][42] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][42] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][42] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][42] ),
    .S0(net1393),
    .S1(net1386),
    .X(_2357_));
 sky130_fd_sc_hd__mux2_2 _4461_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[42] ),
    .A1(_2357_),
    .S(net713),
    .X(net455));
 sky130_fd_sc_hd__mux4_2 _4462_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][43] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][43] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][43] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][43] ),
    .S0(net1395),
    .S1(net1388),
    .X(_2358_));
 sky130_fd_sc_hd__mux2_1 _4463_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[43] ),
    .A1(_2358_),
    .S(net713),
    .X(net456));
 sky130_fd_sc_hd__mux4_2 _4464_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][44] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][44] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][44] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][44] ),
    .S0(net1398),
    .S1(net1390),
    .X(_2359_));
 sky130_fd_sc_hd__mux2_2 _4465_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[44] ),
    .A1(_2359_),
    .S(net718),
    .X(net457));
 sky130_fd_sc_hd__mux4_2 _4466_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][45] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][45] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][45] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][45] ),
    .S0(net1399),
    .S1(net1391),
    .X(_2360_));
 sky130_fd_sc_hd__mux2_1 _4467_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[45] ),
    .A1(_2360_),
    .S(net714),
    .X(net458));
 sky130_fd_sc_hd__mux4_2 _4468_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][46] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][46] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][46] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][46] ),
    .S0(net1392),
    .S1(net1385),
    .X(_2361_));
 sky130_fd_sc_hd__mux2_1 _4469_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[46] ),
    .A1(_2361_),
    .S(net713),
    .X(net459));
 sky130_fd_sc_hd__mux4_2 _4470_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][47] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][47] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][47] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][47] ),
    .S0(net1392),
    .S1(net1385),
    .X(_2362_));
 sky130_fd_sc_hd__mux2_1 _4471_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[47] ),
    .A1(_2362_),
    .S(net715),
    .X(net460));
 sky130_fd_sc_hd__mux4_2 _4472_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][48] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][48] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][48] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][48] ),
    .S0(net1394),
    .S1(net1387),
    .X(_2363_));
 sky130_fd_sc_hd__mux2_1 _4473_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[48] ),
    .A1(_2363_),
    .S(net714),
    .X(net462));
 sky130_fd_sc_hd__mux4_2 _4474_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][49] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][49] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][49] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][49] ),
    .S0(net1392),
    .S1(net1386),
    .X(_2364_));
 sky130_fd_sc_hd__mux2_1 _4475_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[49] ),
    .A1(_2364_),
    .S(net715),
    .X(net463));
 sky130_fd_sc_hd__mux4_2 _4476_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][53] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][53] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][53] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][53] ),
    .S0(net1394),
    .S1(net1387),
    .X(_2365_));
 sky130_fd_sc_hd__mux2_2 _4477_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[53] ),
    .A1(_2365_),
    .S(net716),
    .X(net430));
 sky130_fd_sc_hd__mux4_2 _4478_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][54] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][54] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][54] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][54] ),
    .S0(net1394),
    .S1(net1387),
    .X(_2366_));
 sky130_fd_sc_hd__mux2_1 _4479_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[54] ),
    .A1(_2366_),
    .S(net715),
    .X(net431));
 sky130_fd_sc_hd__mux4_2 _4480_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][55] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][55] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][55] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][55] ),
    .S0(net1394),
    .S1(net1387),
    .X(_2367_));
 sky130_fd_sc_hd__mux2_2 _4481_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[55] ),
    .A1(_2367_),
    .S(net716),
    .X(net432));
 sky130_fd_sc_hd__mux4_2 _4482_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][56] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][56] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][56] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][56] ),
    .S0(net1393),
    .S1(net1386),
    .X(_2368_));
 sky130_fd_sc_hd__mux2_2 _4483_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[56] ),
    .A1(_2368_),
    .S(net713),
    .X(net433));
 sky130_fd_sc_hd__mux4_2 _4484_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][57] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][57] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][57] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][57] ),
    .S0(net1395),
    .S1(net1388),
    .X(_2369_));
 sky130_fd_sc_hd__mux2_1 _4485_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[57] ),
    .A1(_2369_),
    .S(net713),
    .X(net434));
 sky130_fd_sc_hd__mux4_2 _4486_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][58] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][58] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][58] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][58] ),
    .S0(net1392),
    .S1(net1385),
    .X(_2370_));
 sky130_fd_sc_hd__mux2_2 _4487_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[58] ),
    .A1(_2370_),
    .S(net713),
    .X(net435));
 sky130_fd_sc_hd__mux4_2 _4488_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][59] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][59] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][59] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][59] ),
    .S0(net1394),
    .S1(net1387),
    .X(_2371_));
 sky130_fd_sc_hd__mux2_4 _4489_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[59] ),
    .A1(_2371_),
    .S(net718),
    .X(net436));
 sky130_fd_sc_hd__mux4_2 _4490_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][60] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][60] ),
    .A2(net1788),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][60] ),
    .S0(net1393),
    .S1(net1385),
    .X(_2372_));
 sky130_fd_sc_hd__mux2_1 _4491_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[60] ),
    .A1(_2372_),
    .S(net718),
    .X(net437));
 sky130_fd_sc_hd__mux4_2 _4492_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][61] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][61] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][61] ),
    .A3(net1785),
    .S0(net1392),
    .S1(net1385),
    .X(_2373_));
 sky130_fd_sc_hd__mux2_2 _4493_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[61] ),
    .A1(_2373_),
    .S(net713),
    .X(net429));
 sky130_fd_sc_hd__mux4_2 _4494_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][14] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][14] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][14] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][14] ),
    .S0(net1364),
    .S1(net1357),
    .X(_2374_));
 sky130_fd_sc_hd__mux2_2 _4495_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[14] ),
    .A1(_2374_),
    .S(net775),
    .X(net422));
 sky130_fd_sc_hd__mux4_2 _4496_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][15] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][15] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][15] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][15] ),
    .S0(net1360),
    .S1(net1353),
    .X(_2375_));
 sky130_fd_sc_hd__mux2_1 _4497_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[15] ),
    .A1(_2375_),
    .S(net773),
    .X(net423));
 sky130_fd_sc_hd__mux4_1 _4498_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][16] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][16] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][16] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][16] ),
    .S0(net1362),
    .S1(net1355),
    .X(_2376_));
 sky130_fd_sc_hd__mux2_2 _4499_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[16] ),
    .A1(_2376_),
    .S(net775),
    .X(net424));
 sky130_fd_sc_hd__mux4_1 _4500_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][17] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][17] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][17] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][17] ),
    .S0(net1363),
    .S1(net1356),
    .X(_2377_));
 sky130_fd_sc_hd__mux2_4 _4501_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[17] ),
    .A1(_2377_),
    .S(net775),
    .X(net425));
 sky130_fd_sc_hd__mux4_2 _4502_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][18] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][18] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][18] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][18] ),
    .S0(net1364),
    .S1(net1357),
    .X(_2378_));
 sky130_fd_sc_hd__mux2_1 _4503_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[18] ),
    .A1(_2378_),
    .S(net773),
    .X(net390));
 sky130_fd_sc_hd__mux4_2 _4504_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][19] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][19] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][19] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][19] ),
    .S0(net1363),
    .S1(net1356),
    .X(_2379_));
 sky130_fd_sc_hd__mux2_1 _4505_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[19] ),
    .A1(_2379_),
    .S(net774),
    .X(net401));
 sky130_fd_sc_hd__mux4_1 _4506_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][20] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][20] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][20] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][20] ),
    .S0(net1362),
    .S1(net1355),
    .X(_2380_));
 sky130_fd_sc_hd__mux2_2 _4507_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[20] ),
    .A1(_2380_),
    .S(net776),
    .X(net412));
 sky130_fd_sc_hd__mux4_1 _4508_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][21] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][21] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][21] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][21] ),
    .S0(net1362),
    .S1(net1355),
    .X(_2381_));
 sky130_fd_sc_hd__mux2_2 _4509_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[21] ),
    .A1(_2381_),
    .S(net775),
    .X(net415));
 sky130_fd_sc_hd__mux4_2 _4510_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][22] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][22] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][22] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][22] ),
    .S0(net1364),
    .S1(net1357),
    .X(_2382_));
 sky130_fd_sc_hd__mux2_2 _4511_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[22] ),
    .A1(_2382_),
    .S(net776),
    .X(net416));
 sky130_fd_sc_hd__mux4_2 _4512_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][23] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][23] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][23] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][23] ),
    .S0(net1363),
    .S1(net1356),
    .X(_2383_));
 sky130_fd_sc_hd__mux2_1 _4513_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[23] ),
    .A1(_2383_),
    .S(net778),
    .X(net417));
 sky130_fd_sc_hd__mux4_1 _4514_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][24] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][24] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][24] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][24] ),
    .S0(net1360),
    .S1(net1353),
    .X(_2384_));
 sky130_fd_sc_hd__mux2_1 _4515_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[24] ),
    .A1(_2384_),
    .S(net774),
    .X(net418));
 sky130_fd_sc_hd__mux4_1 _4516_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][25] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][25] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][25] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][25] ),
    .S0(net1364),
    .S1(net1357),
    .X(_2385_));
 sky130_fd_sc_hd__mux2_4 _4517_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[25] ),
    .A1(_2385_),
    .S(net777),
    .X(net419));
 sky130_fd_sc_hd__mux4_2 _4518_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][26] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][26] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][26] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][26] ),
    .S0(net1363),
    .S1(net1356),
    .X(_2386_));
 sky130_fd_sc_hd__mux2_2 _4519_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[26] ),
    .A1(_2386_),
    .S(net776),
    .X(net420));
 sky130_fd_sc_hd__mux4_2 _4520_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][27] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][27] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][27] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][27] ),
    .S0(net1364),
    .S1(net1357),
    .X(_2387_));
 sky130_fd_sc_hd__mux2_2 _4521_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[27] ),
    .A1(_2387_),
    .S(net776),
    .X(net421));
 sky130_fd_sc_hd__mux4_1 _4522_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][28] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][28] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][28] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][28] ),
    .S0(net1364),
    .S1(net1357),
    .X(_2388_));
 sky130_fd_sc_hd__mux2_4 _4523_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[28] ),
    .A1(_2388_),
    .S(net777),
    .X(net391));
 sky130_fd_sc_hd__mux4_2 _4524_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][29] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][29] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][29] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][29] ),
    .S0(net1364),
    .S1(net1357),
    .X(_2389_));
 sky130_fd_sc_hd__mux2_2 _4525_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[29] ),
    .A1(_2389_),
    .S(net775),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 _4526_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][30] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][30] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][30] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][30] ),
    .S0(net1364),
    .S1(net1358),
    .X(_2390_));
 sky130_fd_sc_hd__mux2_4 _4527_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[30] ),
    .A1(_2390_),
    .S(net777),
    .X(net393));
 sky130_fd_sc_hd__mux4_1 _4528_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][31] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][31] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][31] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][31] ),
    .S0(net1360),
    .S1(net1353),
    .X(_2391_));
 sky130_fd_sc_hd__mux2_1 _4529_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[31] ),
    .A1(_2391_),
    .S(net774),
    .X(net394));
 sky130_fd_sc_hd__mux4_2 _4530_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][32] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][32] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][32] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][32] ),
    .S0(net1362),
    .S1(net1355),
    .X(_2392_));
 sky130_fd_sc_hd__mux2_1 _4531_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[32] ),
    .A1(_2392_),
    .S(net774),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 _4532_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][33] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][33] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][33] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][33] ),
    .S0(net1359),
    .S1(net1352),
    .X(_2393_));
 sky130_fd_sc_hd__mux2_1 _4533_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[33] ),
    .A1(_2393_),
    .S(net772),
    .X(net396));
 sky130_fd_sc_hd__mux4_2 _4534_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][34] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][34] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][34] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][34] ),
    .S0(net1363),
    .S1(net1356),
    .X(_2394_));
 sky130_fd_sc_hd__mux2_2 _4535_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[34] ),
    .A1(_2394_),
    .S(net778),
    .X(net397));
 sky130_fd_sc_hd__mux4_2 _4536_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][35] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][35] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][35] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][35] ),
    .S0(net1364),
    .S1(net1357),
    .X(_2395_));
 sky130_fd_sc_hd__mux2_2 _4537_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[35] ),
    .A1(_2395_),
    .S(net776),
    .X(net398));
 sky130_fd_sc_hd__mux4_1 _4538_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][36] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][36] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][36] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][36] ),
    .S0(net1359),
    .S1(net1352),
    .X(_2396_));
 sky130_fd_sc_hd__mux2_1 _4539_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[36] ),
    .A1(_2396_),
    .S(net772),
    .X(net399));
 sky130_fd_sc_hd__mux4_2 _4540_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][37] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][37] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][37] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][37] ),
    .S0(net1363),
    .S1(net1356),
    .X(_2397_));
 sky130_fd_sc_hd__mux2_1 _4541_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[37] ),
    .A1(_2397_),
    .S(net773),
    .X(net400));
 sky130_fd_sc_hd__mux4_1 _4542_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][38] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][38] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][38] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][38] ),
    .S0(net1362),
    .S1(net1355),
    .X(_2398_));
 sky130_fd_sc_hd__mux2_2 _4543_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[38] ),
    .A1(_2398_),
    .S(net775),
    .X(net402));
 sky130_fd_sc_hd__mux4_2 _4544_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][39] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][39] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][39] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][39] ),
    .S0(net1359),
    .S1(net1352),
    .X(_2399_));
 sky130_fd_sc_hd__mux2_1 _4545_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[39] ),
    .A1(_2399_),
    .S(net772),
    .X(net403));
 sky130_fd_sc_hd__mux4_1 _4546_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][40] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][40] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][40] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][40] ),
    .S0(net1361),
    .S1(net1354),
    .X(_2400_));
 sky130_fd_sc_hd__mux2_1 _4547_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[40] ),
    .A1(_2400_),
    .S(net772),
    .X(net404));
 sky130_fd_sc_hd__mux4_1 _4548_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][41] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][41] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][41] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][41] ),
    .S0(net1362),
    .S1(net1355),
    .X(_2401_));
 sky130_fd_sc_hd__mux2_2 _4549_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[41] ),
    .A1(_2401_),
    .S(net776),
    .X(net405));
 sky130_fd_sc_hd__mux4_2 _4550_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][42] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][42] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][42] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][42] ),
    .S0(net1363),
    .S1(net1356),
    .X(_2402_));
 sky130_fd_sc_hd__mux2_1 _4551_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[42] ),
    .A1(_2402_),
    .S(net772),
    .X(net406));
 sky130_fd_sc_hd__mux4_2 _4552_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][43] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][43] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][43] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][43] ),
    .S0(net1360),
    .S1(net1353),
    .X(_2403_));
 sky130_fd_sc_hd__mux2_1 _4553_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[43] ),
    .A1(_2403_),
    .S(net774),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 _4554_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][44] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][44] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][44] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][44] ),
    .S0(net1359),
    .S1(net1352),
    .X(_2404_));
 sky130_fd_sc_hd__mux2_1 _4555_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[44] ),
    .A1(_2404_),
    .S(net772),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 _4556_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][45] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][45] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][45] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][45] ),
    .S0(net1365),
    .S1(net1358),
    .X(_2405_));
 sky130_fd_sc_hd__mux2_4 _4557_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[45] ),
    .A1(_2405_),
    .S(net777),
    .X(net409));
 sky130_fd_sc_hd__mux4_2 _4558_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][46] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][46] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][46] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][46] ),
    .S0(net1365),
    .S1(net1358),
    .X(_2406_));
 sky130_fd_sc_hd__mux2_2 _4559_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[46] ),
    .A1(_2406_),
    .S(net775),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 _4560_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][47] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][47] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][47] ),
    .A3(net1951),
    .S0(net1359),
    .S1(net1352),
    .X(_2407_));
 sky130_fd_sc_hd__mux2_1 _4561_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[47] ),
    .A1(_2407_),
    .S(net772),
    .X(net411));
 sky130_fd_sc_hd__mux4_2 _4562_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][48] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][48] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][48] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][48] ),
    .S0(net1359),
    .S1(net1352),
    .X(_2408_));
 sky130_fd_sc_hd__mux2_1 _4563_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[48] ),
    .A1(_2408_),
    .S(net772),
    .X(net413));
 sky130_fd_sc_hd__mux4_1 _4564_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][49] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][49] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][49] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][49] ),
    .S0(net1359),
    .S1(net1352),
    .X(_2409_));
 sky130_fd_sc_hd__mux2_1 _4565_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[49] ),
    .A1(_2409_),
    .S(net772),
    .X(net414));
 sky130_fd_sc_hd__mux4_1 _4566_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][53] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][53] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][53] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][53] ),
    .S0(net1361),
    .S1(net1354),
    .X(_2410_));
 sky130_fd_sc_hd__mux2_1 _4567_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[53] ),
    .A1(_2410_),
    .S(net773),
    .X(net382));
 sky130_fd_sc_hd__mux4_1 _4568_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][54] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][54] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][54] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][54] ),
    .S0(net1360),
    .S1(net1353),
    .X(_2411_));
 sky130_fd_sc_hd__mux2_2 _4569_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[54] ),
    .A1(_2411_),
    .S(net774),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 _4570_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][55] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][55] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][55] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][55] ),
    .S0(net1360),
    .S1(net1353),
    .X(_2412_));
 sky130_fd_sc_hd__mux2_2 _4571_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[55] ),
    .A1(_2412_),
    .S(net774),
    .X(net384));
 sky130_fd_sc_hd__mux4_1 _4572_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][56] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][56] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][56] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][56] ),
    .S0(net1361),
    .S1(net1354),
    .X(_2413_));
 sky130_fd_sc_hd__mux2_2 _4573_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[56] ),
    .A1(_2413_),
    .S(net774),
    .X(net385));
 sky130_fd_sc_hd__mux4_2 _4574_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][57] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][57] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][57] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][57] ),
    .S0(net1361),
    .S1(net1354),
    .X(_2414_));
 sky130_fd_sc_hd__mux2_1 _4575_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[57] ),
    .A1(_2414_),
    .S(net772),
    .X(net386));
 sky130_fd_sc_hd__mux4_1 _4576_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][58] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][58] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][58] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][58] ),
    .S0(net1360),
    .S1(net1353),
    .X(_2415_));
 sky130_fd_sc_hd__mux2_2 _4577_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[58] ),
    .A1(_2415_),
    .S(net774),
    .X(net387));
 sky130_fd_sc_hd__mux4_1 _4578_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][59] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][59] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][59] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][59] ),
    .S0(net1361),
    .S1(net1354),
    .X(_2416_));
 sky130_fd_sc_hd__mux2_1 _4579_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[59] ),
    .A1(_2416_),
    .S(net773),
    .X(net388));
 sky130_fd_sc_hd__and2b_1 _4580_ (.A_N(_1719_),
    .B(net712),
    .X(_2417_));
 sky130_fd_sc_hd__mux2_1 _4581_ (.A0(s0_wbd_lack_i),
    .A1(s0_wbd_ack_i),
    .S(_2417_),
    .X(_2418_));
 sky130_fd_sc_hd__inv_2 _4582_ (.A(net570),
    .Y(_2419_));
 sky130_fd_sc_hd__nand2_1 _4583_ (.A(_1721_),
    .B(net380),
    .Y(_2420_));
 sky130_fd_sc_hd__a211o_1 _4584_ (.A1(_1715_),
    .A2(_2419_),
    .B1(_2420_),
    .C1(_1722_),
    .X(_2421_));
 sky130_fd_sc_hd__nand3_1 _4585_ (.A(_1812_),
    .B(_1815_),
    .C(_1817_),
    .Y(_2422_));
 sky130_fd_sc_hd__or3b_4 _4586_ (.A(net738),
    .B(net712),
    .C_N(net2049),
    .X(_2423_));
 sky130_fd_sc_hd__inv_2 _4587_ (.A(_2423_),
    .Y(_2424_));
 sky130_fd_sc_hd__or4_1 _4588_ (.A(_1815_),
    .B(_1816_),
    .C(_1817_),
    .D(_2423_),
    .X(_2425_));
 sky130_fd_sc_hd__o211a_4 _4589_ (.A1(net712),
    .A2(_2422_),
    .B1(_2425_),
    .C1(_2421_),
    .X(net341));
 sky130_fd_sc_hd__mux4_2 _4590_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][0] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][0] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][0] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][0] ),
    .S0(net1338),
    .S1(net1328),
    .X(_2426_));
 sky130_fd_sc_hd__mux2_2 _4591_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[0] ),
    .A1(_2426_),
    .S(net829),
    .X(net331));
 sky130_fd_sc_hd__mux4_2 _4592_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][14] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][14] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][14] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][14] ),
    .S0(net1342),
    .S1(net1332),
    .X(_2427_));
 sky130_fd_sc_hd__mux2_2 _4593_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[14] ),
    .A1(_2427_),
    .S(net829),
    .X(net375));
 sky130_fd_sc_hd__mux4_2 _4594_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][15] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][15] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][15] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][15] ),
    .S0(net1334),
    .S1(net1324),
    .X(_2428_));
 sky130_fd_sc_hd__mux2_1 _4595_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[15] ),
    .A1(_2428_),
    .S(net826),
    .X(net376));
 sky130_fd_sc_hd__mux4_2 _4596_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][16] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][16] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][16] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][16] ),
    .S0(net1335),
    .S1(net1325),
    .X(_2429_));
 sky130_fd_sc_hd__mux2_1 _4597_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[16] ),
    .A1(_2429_),
    .S(net825),
    .X(net377));
 sky130_fd_sc_hd__mux4_1 _4598_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][17] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][17] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][17] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][17] ),
    .S0(net1335),
    .S1(net1325),
    .X(_2430_));
 sky130_fd_sc_hd__mux2_1 _4599_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[17] ),
    .A1(_2430_),
    .S(net824),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 _4600_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][18] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][18] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][18] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][18] ),
    .S0(net1340),
    .S1(net1330),
    .X(_2431_));
 sky130_fd_sc_hd__mux2_4 _4601_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[18] ),
    .A1(_2431_),
    .S(net831),
    .X(net343));
 sky130_fd_sc_hd__mux4_1 _4602_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][19] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][19] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][19] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][19] ),
    .S0(net1340),
    .S1(net1330),
    .X(_2432_));
 sky130_fd_sc_hd__mux2_4 _4603_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[19] ),
    .A1(_2432_),
    .S(net832),
    .X(net354));
 sky130_fd_sc_hd__mux4_1 _4604_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][20] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][20] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][20] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][20] ),
    .S0(net1341),
    .S1(net1331),
    .X(_2433_));
 sky130_fd_sc_hd__mux2_4 _4605_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[20] ),
    .A1(_2433_),
    .S(net831),
    .X(net365));
 sky130_fd_sc_hd__mux4_2 _4606_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][21] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][21] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][21] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][21] ),
    .S0(net1340),
    .S1(net1330),
    .X(_2434_));
 sky130_fd_sc_hd__mux2_4 _4607_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[21] ),
    .A1(_2434_),
    .S(net832),
    .X(net368));
 sky130_fd_sc_hd__mux4_1 _4608_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][22] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][22] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][22] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][22] ),
    .S0(net1338),
    .S1(net1328),
    .X(_2435_));
 sky130_fd_sc_hd__mux2_2 _4609_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[22] ),
    .A1(_2435_),
    .S(net832),
    .X(net369));
 sky130_fd_sc_hd__mux4_2 _4610_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][23] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][23] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][23] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][23] ),
    .S0(net1339),
    .S1(net1329),
    .X(_2436_));
 sky130_fd_sc_hd__mux2_2 _4611_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[23] ),
    .A1(_2436_),
    .S(net829),
    .X(net370));
 sky130_fd_sc_hd__mux4_1 _4612_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][24] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][24] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][24] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][24] ),
    .S0(net1339),
    .S1(net1329),
    .X(_2437_));
 sky130_fd_sc_hd__mux2_4 _4613_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[24] ),
    .A1(_2437_),
    .S(net832),
    .X(net371));
 sky130_fd_sc_hd__mux4_2 _4614_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][25] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][25] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][25] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][25] ),
    .S0(net1337),
    .S1(net1327),
    .X(_2438_));
 sky130_fd_sc_hd__mux2_1 _4615_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[25] ),
    .A1(_2438_),
    .S(net827),
    .X(net372));
 sky130_fd_sc_hd__mux4_2 _4616_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][26] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][26] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][26] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][26] ),
    .S0(net1339),
    .S1(net1329),
    .X(_2439_));
 sky130_fd_sc_hd__mux2_2 _4617_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[26] ),
    .A1(_2439_),
    .S(net829),
    .X(net373));
 sky130_fd_sc_hd__mux4_1 _4618_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][27] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][27] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][27] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][27] ),
    .S0(net1341),
    .S1(net1331),
    .X(_2440_));
 sky130_fd_sc_hd__mux2_4 _4619_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[27] ),
    .A1(_2440_),
    .S(net831),
    .X(net374));
 sky130_fd_sc_hd__mux4_2 _4620_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][28] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][28] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][28] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][28] ),
    .S0(net1340),
    .S1(net1330),
    .X(_2441_));
 sky130_fd_sc_hd__mux2_2 _4621_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[28] ),
    .A1(_2441_),
    .S(net829),
    .X(net344));
 sky130_fd_sc_hd__mux4_1 _4622_ (.A0(net1957),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][29] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][29] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][29] ),
    .S0(net1341),
    .S1(net1331),
    .X(_2442_));
 sky130_fd_sc_hd__mux2_1 _4623_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[29] ),
    .A1(_2442_),
    .S(net831),
    .X(net345));
 sky130_fd_sc_hd__mux4_1 _4624_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][30] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][30] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][30] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][30] ),
    .S0(net1334),
    .S1(net1324),
    .X(_2443_));
 sky130_fd_sc_hd__mux2_1 _4625_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[30] ),
    .A1(_2443_),
    .S(net827),
    .X(net346));
 sky130_fd_sc_hd__mux4_1 _4626_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][31] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][31] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][31] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][31] ),
    .S0(net1336),
    .S1(net1326),
    .X(_2444_));
 sky130_fd_sc_hd__mux2_1 _4627_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[31] ),
    .A1(_2444_),
    .S(net830),
    .X(net347));
 sky130_fd_sc_hd__mux4_1 _4628_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][32] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][32] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][32] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][32] ),
    .S0(net1341),
    .S1(net1331),
    .X(_2445_));
 sky130_fd_sc_hd__mux2_1 _4629_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[32] ),
    .A1(_2445_),
    .S(net831),
    .X(net348));
 sky130_fd_sc_hd__mux4_2 _4630_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][33] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][33] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][33] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][33] ),
    .S0(net1338),
    .S1(net1328),
    .X(_2446_));
 sky130_fd_sc_hd__mux2_2 _4631_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[33] ),
    .A1(_2446_),
    .S(net829),
    .X(net349));
 sky130_fd_sc_hd__mux4_2 _4632_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][34] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][34] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][34] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][34] ),
    .S0(net1336),
    .S1(net1326),
    .X(_2447_));
 sky130_fd_sc_hd__mux2_1 _4633_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[34] ),
    .A1(_2447_),
    .S(net827),
    .X(net350));
 sky130_fd_sc_hd__mux4_2 _4634_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][35] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][35] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][35] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][35] ),
    .S0(net1340),
    .S1(net1330),
    .X(_2448_));
 sky130_fd_sc_hd__mux2_1 _4635_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[35] ),
    .A1(_2448_),
    .S(net830),
    .X(net351));
 sky130_fd_sc_hd__mux4_1 _4636_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][36] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][36] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][36] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][36] ),
    .S0(net1334),
    .S1(net1324),
    .X(_2449_));
 sky130_fd_sc_hd__mux2_1 _4637_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[36] ),
    .A1(_2449_),
    .S(net828),
    .X(net352));
 sky130_fd_sc_hd__mux4_1 _4638_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][37] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][37] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][37] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][37] ),
    .S0(net1338),
    .S1(net1328),
    .X(_2450_));
 sky130_fd_sc_hd__mux2_4 _4639_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[37] ),
    .A1(_2450_),
    .S(net832),
    .X(net353));
 sky130_fd_sc_hd__mux4_1 _4640_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][38] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][38] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][38] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][38] ),
    .S0(net1334),
    .S1(net1324),
    .X(_2451_));
 sky130_fd_sc_hd__mux2_1 _4641_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[38] ),
    .A1(_2451_),
    .S(net827),
    .X(net355));
 sky130_fd_sc_hd__mux4_1 _4642_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][39] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][39] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][39] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][39] ),
    .S0(net1339),
    .S1(net1329),
    .X(_2452_));
 sky130_fd_sc_hd__mux2_4 _4643_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[39] ),
    .A1(_2452_),
    .S(net832),
    .X(net356));
 sky130_fd_sc_hd__mux4_1 _4644_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][40] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][40] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][40] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][40] ),
    .S0(net1336),
    .S1(net1326),
    .X(_2453_));
 sky130_fd_sc_hd__mux2_1 _4645_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[40] ),
    .A1(_2453_),
    .S(net828),
    .X(net357));
 sky130_fd_sc_hd__mux4_2 _4646_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][41] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][41] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][41] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][41] ),
    .S0(net1339),
    .S1(net1329),
    .X(_2454_));
 sky130_fd_sc_hd__mux2_1 _4647_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[41] ),
    .A1(_2454_),
    .S(net827),
    .X(net358));
 sky130_fd_sc_hd__mux4_2 _4648_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][42] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][42] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][42] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][42] ),
    .S0(net1337),
    .S1(net1327),
    .X(_2455_));
 sky130_fd_sc_hd__mux2_1 _4649_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[42] ),
    .A1(_2455_),
    .S(net830),
    .X(net359));
 sky130_fd_sc_hd__mux4_2 _4650_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][43] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][43] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][43] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][43] ),
    .S0(net1338),
    .S1(net1328),
    .X(_2456_));
 sky130_fd_sc_hd__mux2_2 _4651_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[43] ),
    .A1(_2456_),
    .S(net829),
    .X(net360));
 sky130_fd_sc_hd__mux4_1 _4652_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][44] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][44] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][44] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][44] ),
    .S0(net1337),
    .S1(net1327),
    .X(_2457_));
 sky130_fd_sc_hd__mux2_2 _4653_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[44] ),
    .A1(_2457_),
    .S(net830),
    .X(net361));
 sky130_fd_sc_hd__mux4_2 _4654_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][45] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][45] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][45] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][45] ),
    .S0(net1337),
    .S1(net1327),
    .X(_2458_));
 sky130_fd_sc_hd__mux2_2 _4655_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[45] ),
    .A1(_2458_),
    .S(net830),
    .X(net362));
 sky130_fd_sc_hd__mux4_1 _4656_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][46] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][46] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][46] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][46] ),
    .S0(net1335),
    .S1(net1325),
    .X(_2459_));
 sky130_fd_sc_hd__mux2_1 _4657_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[46] ),
    .A1(_2459_),
    .S(net826),
    .X(net363));
 sky130_fd_sc_hd__mux4_2 _4658_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][47] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][47] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][47] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][47] ),
    .S0(net1337),
    .S1(net1327),
    .X(_2460_));
 sky130_fd_sc_hd__mux2_2 _4659_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[47] ),
    .A1(_2460_),
    .S(net830),
    .X(net364));
 sky130_fd_sc_hd__mux4_2 _4660_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][48] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][48] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][48] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][48] ),
    .S0(net1338),
    .S1(net1328),
    .X(_2461_));
 sky130_fd_sc_hd__mux2_2 _4661_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[48] ),
    .A1(_2461_),
    .S(net832),
    .X(net366));
 sky130_fd_sc_hd__mux4_2 _4662_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][49] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][49] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][49] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][49] ),
    .S0(net1335),
    .S1(net1325),
    .X(_2462_));
 sky130_fd_sc_hd__mux2_1 _4663_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[49] ),
    .A1(_2462_),
    .S(net827),
    .X(net367));
 sky130_fd_sc_hd__mux4_2 _4664_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][53] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][53] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][53] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][53] ),
    .S0(net1338),
    .S1(net1328),
    .X(_2463_));
 sky130_fd_sc_hd__mux2_1 _4665_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[53] ),
    .A1(_2463_),
    .S(net827),
    .X(net321));
 sky130_fd_sc_hd__mux4_2 _4666_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][54] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][54] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][54] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][54] ),
    .S0(net1342),
    .S1(net1327),
    .X(_2464_));
 sky130_fd_sc_hd__mux2_2 _4667_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[54] ),
    .A1(_2464_),
    .S(net830),
    .X(net324));
 sky130_fd_sc_hd__mux4_2 _4668_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][55] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][55] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][55] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][55] ),
    .S0(net1338),
    .S1(net1328),
    .X(_2465_));
 sky130_fd_sc_hd__mux2_2 _4669_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[55] ),
    .A1(_2465_),
    .S(net829),
    .X(net325));
 sky130_fd_sc_hd__mux4_2 _4670_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][56] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][56] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][56] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][56] ),
    .S0(net1337),
    .S1(net1327),
    .X(_2466_));
 sky130_fd_sc_hd__mux2_2 _4671_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[56] ),
    .A1(_2466_),
    .S(net829),
    .X(net326));
 sky130_fd_sc_hd__mux4_1 _4672_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][57] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][57] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][57] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][57] ),
    .S0(net1335),
    .S1(net1325),
    .X(_2467_));
 sky130_fd_sc_hd__mux2_1 _4673_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[57] ),
    .A1(_2467_),
    .S(net828),
    .X(net327));
 sky130_fd_sc_hd__mux4_1 _4674_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][58] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][58] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][58] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][58] ),
    .S0(net1333),
    .S1(net1325),
    .X(_2468_));
 sky130_fd_sc_hd__mux2_1 _4675_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[58] ),
    .A1(_2468_),
    .S(net824),
    .X(net328));
 sky130_fd_sc_hd__mux4_2 _4676_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][59] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][59] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][59] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][59] ),
    .S0(net1337),
    .S1(net1327),
    .X(_2469_));
 sky130_fd_sc_hd__mux2_2 _4677_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[59] ),
    .A1(_2469_),
    .S(net829),
    .X(net329));
 sky130_fd_sc_hd__mux4_2 _4678_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][60] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][60] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][60] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][60] ),
    .S0(net1336),
    .S1(net1326),
    .X(_2470_));
 sky130_fd_sc_hd__mux2_1 _4679_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[60] ),
    .A1(_2470_),
    .S(net825),
    .X(net330));
 sky130_fd_sc_hd__mux4_2 _4680_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][61] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][61] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][61] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][61] ),
    .S0(net1337),
    .S1(net1327),
    .X(_2471_));
 sky130_fd_sc_hd__mux2_1 _4681_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[61] ),
    .A1(_2471_),
    .S(net825),
    .X(net301));
 sky130_fd_sc_hd__mux4_2 _4682_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][62] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][62] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][62] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][62] ),
    .S0(net1334),
    .S1(net1324),
    .X(_2472_));
 sky130_fd_sc_hd__mux2_1 _4683_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[62] ),
    .A1(_2472_),
    .S(net825),
    .X(net302));
 sky130_fd_sc_hd__mux4_2 _4684_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][63] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][63] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][63] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][63] ),
    .S0(net1336),
    .S1(net1326),
    .X(_2473_));
 sky130_fd_sc_hd__mux2_1 _4685_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[63] ),
    .A1(_2473_),
    .S(net825),
    .X(net303));
 sky130_fd_sc_hd__mux4_2 _4686_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][64] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][64] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][64] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][64] ),
    .S0(net1336),
    .S1(net1326),
    .X(_2474_));
 sky130_fd_sc_hd__mux2_2 _4687_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[64] ),
    .A1(_2474_),
    .S(net833),
    .X(net304));
 sky130_fd_sc_hd__mux4_2 _4688_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][65] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][65] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][65] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][65] ),
    .S0(net1333),
    .S1(net1323),
    .X(_2475_));
 sky130_fd_sc_hd__mux2_1 _4689_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[65] ),
    .A1(_2475_),
    .S(net826),
    .X(net305));
 sky130_fd_sc_hd__mux4_2 _4690_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][66] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][66] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][66] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][66] ),
    .S0(net1333),
    .S1(net1323),
    .X(_2476_));
 sky130_fd_sc_hd__mux2_1 _4691_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[66] ),
    .A1(_2476_),
    .S(net824),
    .X(net306));
 sky130_fd_sc_hd__mux4_2 _4692_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][67] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][67] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][67] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][67] ),
    .S0(net1336),
    .S1(net1326),
    .X(_2477_));
 sky130_fd_sc_hd__mux2_1 _4693_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[67] ),
    .A1(_2477_),
    .S(net826),
    .X(net307));
 sky130_fd_sc_hd__mux4_2 _4694_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][68] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][68] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][68] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][68] ),
    .S0(net1336),
    .S1(net1326),
    .X(_2478_));
 sky130_fd_sc_hd__mux2_1 _4695_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[68] ),
    .A1(_2478_),
    .S(net826),
    .X(net308));
 sky130_fd_sc_hd__mux4_2 _4696_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][69] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][69] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][69] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][69] ),
    .S0(net1333),
    .S1(net1323),
    .X(_2479_));
 sky130_fd_sc_hd__mux2_1 _4697_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[69] ),
    .A1(_2479_),
    .S(net826),
    .X(net309));
 sky130_fd_sc_hd__mux4_1 _4698_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][70] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][70] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][70] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][70] ),
    .S0(net1333),
    .S1(net1323),
    .X(_2480_));
 sky130_fd_sc_hd__mux2_1 _4699_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[70] ),
    .A1(_2480_),
    .S(net824),
    .X(net310));
 sky130_fd_sc_hd__mux4_2 _4700_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][71] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][71] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][71] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][71] ),
    .S0(net1336),
    .S1(net1326),
    .X(_2481_));
 sky130_fd_sc_hd__mux2_1 _4701_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[71] ),
    .A1(_2481_),
    .S(net825),
    .X(net311));
 sky130_fd_sc_hd__mux4_2 _4702_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][72] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][72] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][72] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][72] ),
    .S0(net1334),
    .S1(net1324),
    .X(_2482_));
 sky130_fd_sc_hd__mux2_1 _4703_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[72] ),
    .A1(_2482_),
    .S(net828),
    .X(net312));
 sky130_fd_sc_hd__mux4_2 _4704_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][73] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][73] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][73] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][73] ),
    .S0(net1336),
    .S1(net1326),
    .X(_2483_));
 sky130_fd_sc_hd__mux2_2 _4705_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[73] ),
    .A1(_2483_),
    .S(net830),
    .X(net313));
 sky130_fd_sc_hd__mux4_2 _4706_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][74] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][74] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][74] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][74] ),
    .S0(net1333),
    .S1(net1323),
    .X(_2484_));
 sky130_fd_sc_hd__mux2_1 _4707_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[74] ),
    .A1(_2484_),
    .S(net824),
    .X(net314));
 sky130_fd_sc_hd__mux4_2 _4708_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][75] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][75] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][75] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][75] ),
    .S0(net1334),
    .S1(net1324),
    .X(_2485_));
 sky130_fd_sc_hd__mux2_1 _4709_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[75] ),
    .A1(_2485_),
    .S(net825),
    .X(net315));
 sky130_fd_sc_hd__mux4_2 _4710_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][76] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][76] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][76] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][76] ),
    .S0(net1334),
    .S1(net1324),
    .X(_2486_));
 sky130_fd_sc_hd__mux2_1 _4711_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[76] ),
    .A1(_2486_),
    .S(net824),
    .X(net316));
 sky130_fd_sc_hd__mux4_2 _4712_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][77] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][77] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][77] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][77] ),
    .S0(net1333),
    .S1(net1323),
    .X(_2487_));
 sky130_fd_sc_hd__mux2_1 _4713_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[77] ),
    .A1(_2487_),
    .S(net824),
    .X(net317));
 sky130_fd_sc_hd__mux4_2 _4714_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][78] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][78] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][78] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][78] ),
    .S0(net1333),
    .S1(net1323),
    .X(_2488_));
 sky130_fd_sc_hd__mux2_1 _4715_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[78] ),
    .A1(_2488_),
    .S(net825),
    .X(net318));
 sky130_fd_sc_hd__mux4_2 _4716_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][79] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][79] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][79] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][79] ),
    .S0(net1334),
    .S1(net1324),
    .X(_2489_));
 sky130_fd_sc_hd__mux2_1 _4717_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[79] ),
    .A1(_2489_),
    .S(net824),
    .X(net319));
 sky130_fd_sc_hd__mux4_2 _4718_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][80] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][80] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][80] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][80] ),
    .S0(net1333),
    .S1(net1323),
    .X(_2490_));
 sky130_fd_sc_hd__mux2_1 _4719_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[80] ),
    .A1(_2490_),
    .S(net824),
    .X(net320));
 sky130_fd_sc_hd__mux4_2 _4720_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][81] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][81] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][81] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][81] ),
    .S0(net1333),
    .S1(net1323),
    .X(_2491_));
 sky130_fd_sc_hd__mux2_1 _4721_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[81] ),
    .A1(_2491_),
    .S(net824),
    .X(net322));
 sky130_fd_sc_hd__mux4_2 _4722_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[0][82] ),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[1][82] ),
    .A2(\u_s0.u_sync_wbb.u_cmd_if.mem[2][82] ),
    .A3(\u_s0.u_sync_wbb.u_cmd_if.mem[3][82] ),
    .S0(net1335),
    .S1(net1323),
    .X(_2492_));
 sky130_fd_sc_hd__mux2_1 _4723_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[82] ),
    .A1(_2492_),
    .S(net825),
    .X(net323));
 sky130_fd_sc_hd__nand2_1 _4724_ (.A(\u_s0.u_sync_wbb.wbm_lack_o ),
    .B(net1208),
    .Y(_2493_));
 sky130_fd_sc_hd__and3_1 _4725_ (.A(_1741_),
    .B(_1743_),
    .C(_2493_),
    .X(_2494_));
 sky130_fd_sc_hd__and2_1 _4726_ (.A(net1179),
    .B(_1958_),
    .X(_2495_));
 sky130_fd_sc_hd__nand2_1 _4727_ (.A(net1366),
    .B(net1185),
    .Y(_2496_));
 sky130_fd_sc_hd__a22o_1 _4728_ (.A1(_1741_),
    .A2(_1743_),
    .B1(net1157),
    .B2(\u_reg.reg_ack ),
    .X(_2497_));
 sky130_fd_sc_hd__a31o_1 _4729_ (.A1(net1366),
    .A2(net1185),
    .A3(_1853_),
    .B1(_2497_),
    .X(_2498_));
 sky130_fd_sc_hd__a21oi_1 _4730_ (.A1(net1401),
    .A2(net763),
    .B1(_2498_),
    .Y(_2499_));
 sky130_fd_sc_hd__nand2_1 _4731_ (.A(net1401),
    .B(net1179),
    .Y(_2500_));
 sky130_fd_sc_hd__and2_1 _4732_ (.A(net1185),
    .B(_1853_),
    .X(_2501_));
 sky130_fd_sc_hd__nor2_2 _4733_ (.A(_2494_),
    .B(_2499_),
    .Y(net297));
 sky130_fd_sc_hd__a22o_1 _4734_ (.A1(\u_reg.reg_ack ),
    .A2(net1154),
    .B1(net759),
    .B2(net1367),
    .X(_2502_));
 sky130_fd_sc_hd__a22o_1 _4735_ (.A1(\u_s0.u_sync_wbb.wbm_ack_o ),
    .A2(net817),
    .B1(net761),
    .B2(net1402),
    .X(_2503_));
 sky130_fd_sc_hd__or2_1 _4736_ (.A(_2502_),
    .B(_2503_),
    .X(net264));
 sky130_fd_sc_hd__a22o_1 _4737_ (.A1(net1312),
    .A2(net1157),
    .B1(net1142),
    .B2(net818),
    .X(_2504_));
 sky130_fd_sc_hd__a22o_1 _4738_ (.A1(net1141),
    .A2(net761),
    .B1(net757),
    .B2(net1139),
    .X(_2505_));
 sky130_fd_sc_hd__or2_1 _4739_ (.A(_2504_),
    .B(_2505_),
    .X(net265));
 sky130_fd_sc_hd__a22o_1 _4740_ (.A1(\u_reg.reg_rdata[1] ),
    .A2(net1157),
    .B1(net1137),
    .B2(net756),
    .X(_2506_));
 sky130_fd_sc_hd__a22o_1 _4741_ (.A1(net818),
    .A2(_2036_),
    .B1(net1135),
    .B2(net763),
    .X(_2507_));
 sky130_fd_sc_hd__or2_1 _4742_ (.A(_2506_),
    .B(_2507_),
    .X(net276));
 sky130_fd_sc_hd__a22o_1 _4743_ (.A1(\u_reg.reg_rdata[2] ),
    .A2(net1153),
    .B1(net1134),
    .B2(net818),
    .X(_2508_));
 sky130_fd_sc_hd__a22o_1 _4744_ (.A1(net1132),
    .A2(net762),
    .B1(net757),
    .B2(net1130),
    .X(_2509_));
 sky130_fd_sc_hd__or2_1 _4745_ (.A(_2508_),
    .B(_2509_),
    .X(net287));
 sky130_fd_sc_hd__a22o_1 _4746_ (.A1(\u_reg.reg_rdata[3] ),
    .A2(net1153),
    .B1(_2046_),
    .B2(net818),
    .X(_2510_));
 sky130_fd_sc_hd__a22o_1 _4747_ (.A1(net1126),
    .A2(net761),
    .B1(net756),
    .B2(net1128),
    .X(_2511_));
 sky130_fd_sc_hd__or2_1 _4748_ (.A(_2510_),
    .B(_2511_),
    .X(net290));
 sky130_fd_sc_hd__a22o_1 _4749_ (.A1(net1311),
    .A2(net1153),
    .B1(net1122),
    .B2(net757),
    .X(_2512_));
 sky130_fd_sc_hd__a22o_1 _4750_ (.A1(net817),
    .A2(net1125),
    .B1(net1123),
    .B2(net760),
    .X(_2513_));
 sky130_fd_sc_hd__or2_1 _4751_ (.A(_2512_),
    .B(_2513_),
    .X(net291));
 sky130_fd_sc_hd__a22o_1 _4752_ (.A1(\u_reg.reg_rdata[5] ),
    .A2(net1155),
    .B1(net1121),
    .B2(net758),
    .X(_2514_));
 sky130_fd_sc_hd__a22o_1 _4753_ (.A1(net819),
    .A2(_2056_),
    .B1(net1117),
    .B2(net762),
    .X(_2515_));
 sky130_fd_sc_hd__or2_1 _4754_ (.A(_2514_),
    .B(_2515_),
    .X(net292));
 sky130_fd_sc_hd__a22o_1 _4755_ (.A1(\u_reg.reg_rdata[6] ),
    .A2(net1154),
    .B1(net1114),
    .B2(net817),
    .X(_2516_));
 sky130_fd_sc_hd__a22o_1 _4756_ (.A1(net1112),
    .A2(net761),
    .B1(net756),
    .B2(net1115),
    .X(_2517_));
 sky130_fd_sc_hd__or2_1 _4757_ (.A(_2516_),
    .B(_2517_),
    .X(net293));
 sky130_fd_sc_hd__a22o_1 _4758_ (.A1(\u_reg.reg_rdata[7] ),
    .A2(net1155),
    .B1(_2064_),
    .B2(net820),
    .X(_2518_));
 sky130_fd_sc_hd__a22o_1 _4759_ (.A1(net1110),
    .A2(net762),
    .B1(net758),
    .B2(_2067_),
    .X(_2519_));
 sky130_fd_sc_hd__or2_1 _4760_ (.A(_2518_),
    .B(_2519_),
    .X(net294));
 sky130_fd_sc_hd__a22o_1 _4761_ (.A1(\u_reg.reg_rdata[8] ),
    .A2(net1155),
    .B1(net1107),
    .B2(net757),
    .X(_2520_));
 sky130_fd_sc_hd__a22o_1 _4762_ (.A1(net819),
    .A2(_2071_),
    .B1(net1104),
    .B2(net761),
    .X(_2521_));
 sky130_fd_sc_hd__or2_1 _4763_ (.A(_2520_),
    .B(_2521_),
    .X(net295));
 sky130_fd_sc_hd__a22o_1 _4764_ (.A1(\u_reg.reg_rdata[9] ),
    .A2(net1156),
    .B1(_2074_),
    .B2(net758),
    .X(_2522_));
 sky130_fd_sc_hd__a22o_1 _4765_ (.A1(net819),
    .A2(net1101),
    .B1(net1100),
    .B2(net762),
    .X(_2523_));
 sky130_fd_sc_hd__or2_1 _4766_ (.A(_2522_),
    .B(_2523_),
    .X(net296));
 sky130_fd_sc_hd__a22o_1 _4767_ (.A1(\u_reg.reg_rdata[10] ),
    .A2(net1155),
    .B1(_2079_),
    .B2(net758),
    .X(_2524_));
 sky130_fd_sc_hd__a22o_1 _4768_ (.A1(net819),
    .A2(net1097),
    .B1(net1095),
    .B2(net761),
    .X(_2525_));
 sky130_fd_sc_hd__or2_1 _4769_ (.A(_2524_),
    .B(_2525_),
    .X(net266));
 sky130_fd_sc_hd__a22o_1 _4770_ (.A1(net1305),
    .A2(net1153),
    .B1(net1091),
    .B2(net756),
    .X(_2526_));
 sky130_fd_sc_hd__a22o_1 _4771_ (.A1(net818),
    .A2(net1093),
    .B1(net1092),
    .B2(net760),
    .X(_2527_));
 sky130_fd_sc_hd__or2_1 _4772_ (.A(_2526_),
    .B(_2527_),
    .X(net267));
 sky130_fd_sc_hd__a22o_1 _4773_ (.A1(\u_reg.reg_rdata[12] ),
    .A2(net1156),
    .B1(_2089_),
    .B2(net758),
    .X(_2528_));
 sky130_fd_sc_hd__a22o_1 _4774_ (.A1(net820),
    .A2(net1089),
    .B1(net1087),
    .B2(net763),
    .X(_2529_));
 sky130_fd_sc_hd__or2_1 _4775_ (.A(_2528_),
    .B(_2529_),
    .X(net268));
 sky130_fd_sc_hd__a22o_1 _4776_ (.A1(net1303),
    .A2(net1155),
    .B1(_2094_),
    .B2(net757),
    .X(_2530_));
 sky130_fd_sc_hd__a22o_1 _4777_ (.A1(net819),
    .A2(net1084),
    .B1(net1083),
    .B2(net761),
    .X(_2531_));
 sky130_fd_sc_hd__or2_1 _4778_ (.A(_2530_),
    .B(_2531_),
    .X(net269));
 sky130_fd_sc_hd__a22o_1 _4779_ (.A1(net1301),
    .A2(net1156),
    .B1(_2099_),
    .B2(net758),
    .X(_2532_));
 sky130_fd_sc_hd__a22o_1 _4780_ (.A1(net820),
    .A2(net1080),
    .B1(net1079),
    .B2(net762),
    .X(_2533_));
 sky130_fd_sc_hd__or2_1 _4781_ (.A(_2532_),
    .B(_2533_),
    .X(net270));
 sky130_fd_sc_hd__a22o_1 _4782_ (.A1(net1299),
    .A2(net1155),
    .B1(net1077),
    .B2(net819),
    .X(_2534_));
 sky130_fd_sc_hd__a22o_1 _4783_ (.A1(net1076),
    .A2(net763),
    .B1(net757),
    .B2(net1074),
    .X(_2535_));
 sky130_fd_sc_hd__or2_1 _4784_ (.A(_2534_),
    .B(_2535_),
    .X(net271));
 sky130_fd_sc_hd__a22o_1 _4785_ (.A1(net1297),
    .A2(net1155),
    .B1(net1072),
    .B2(net758),
    .X(_2536_));
 sky130_fd_sc_hd__a22o_1 _4786_ (.A1(net819),
    .A2(net1070),
    .B1(net1069),
    .B2(net761),
    .X(_2537_));
 sky130_fd_sc_hd__or2_1 _4787_ (.A(_2536_),
    .B(_2537_),
    .X(net272));
 sky130_fd_sc_hd__a22o_1 _4788_ (.A1(net1295),
    .A2(net1155),
    .B1(net1067),
    .B2(net757),
    .X(_2538_));
 sky130_fd_sc_hd__a22o_1 _4789_ (.A1(net819),
    .A2(net1066),
    .B1(net1064),
    .B2(net761),
    .X(_2539_));
 sky130_fd_sc_hd__or2_1 _4790_ (.A(_2538_),
    .B(_2539_),
    .X(net273));
 sky130_fd_sc_hd__a22o_1 _4791_ (.A1(\u_reg.reg_rdata[18] ),
    .A2(net1157),
    .B1(net1063),
    .B2(_1747_),
    .X(_2540_));
 sky130_fd_sc_hd__a22o_1 _4792_ (.A1(net1061),
    .A2(net760),
    .B1(net756),
    .B2(net1059),
    .X(_2541_));
 sky130_fd_sc_hd__or2_1 _4793_ (.A(_2540_),
    .B(_2541_),
    .X(net274));
 sky130_fd_sc_hd__a22o_1 _4794_ (.A1(\u_reg.reg_rdata[19] ),
    .A2(net1157),
    .B1(_2126_),
    .B2(net818),
    .X(_2542_));
 sky130_fd_sc_hd__a22o_1 _4795_ (.A1(net1056),
    .A2(net762),
    .B1(net758),
    .B2(net1057),
    .X(_2543_));
 sky130_fd_sc_hd__or2_1 _4796_ (.A(_2542_),
    .B(_2543_),
    .X(net275));
 sky130_fd_sc_hd__a22o_1 _4797_ (.A1(net1294),
    .A2(net1153),
    .B1(_2129_),
    .B2(net756),
    .X(_2544_));
 sky130_fd_sc_hd__a22o_1 _4798_ (.A1(net817),
    .A2(net1054),
    .B1(net1052),
    .B2(net760),
    .X(_2545_));
 sky130_fd_sc_hd__or2_1 _4799_ (.A(_2544_),
    .B(_2545_),
    .X(net277));
 sky130_fd_sc_hd__a22o_1 _4800_ (.A1(net1292),
    .A2(net1154),
    .B1(_2137_),
    .B2(net759),
    .X(_2546_));
 sky130_fd_sc_hd__a22o_1 _4801_ (.A1(net817),
    .A2(_2134_),
    .B1(net1049),
    .B2(net760),
    .X(_2547_));
 sky130_fd_sc_hd__or2_1 _4802_ (.A(_2546_),
    .B(_2547_),
    .X(net278));
 sky130_fd_sc_hd__a22o_1 _4803_ (.A1(\u_reg.reg_rdata[22] ),
    .A2(net1154),
    .B1(_2142_),
    .B2(net756),
    .X(_2548_));
 sky130_fd_sc_hd__a22o_1 _4804_ (.A1(net817),
    .A2(net1046),
    .B1(net1045),
    .B2(net763),
    .X(_2549_));
 sky130_fd_sc_hd__or2_1 _4805_ (.A(_2548_),
    .B(_2549_),
    .X(net279));
 sky130_fd_sc_hd__a22o_2 _4806_ (.A1(\u_reg.reg_rdata[23] ),
    .A2(net1157),
    .B1(_2144_),
    .B2(_1747_),
    .X(_2550_));
 sky130_fd_sc_hd__a22o_1 _4807_ (.A1(net1041),
    .A2(net762),
    .B1(net757),
    .B2(_2147_),
    .X(_2551_));
 sky130_fd_sc_hd__or2_1 _4808_ (.A(_2550_),
    .B(_2551_),
    .X(net280));
 sky130_fd_sc_hd__a22o_1 _4809_ (.A1(net1289),
    .A2(net1155),
    .B1(_2152_),
    .B2(net757),
    .X(_2552_));
 sky130_fd_sc_hd__a22o_1 _4810_ (.A1(net819),
    .A2(net1038),
    .B1(net1037),
    .B2(net762),
    .X(_2553_));
 sky130_fd_sc_hd__or2_1 _4811_ (.A(_2552_),
    .B(_2553_),
    .X(net281));
 sky130_fd_sc_hd__a22o_1 _4812_ (.A1(\u_reg.reg_rdata[25] ),
    .A2(net1155),
    .B1(_2154_),
    .B2(net758),
    .X(_2554_));
 sky130_fd_sc_hd__a22o_1 _4813_ (.A1(net819),
    .A2(net1034),
    .B1(net1033),
    .B2(net762),
    .X(_2555_));
 sky130_fd_sc_hd__or2_2 _4814_ (.A(_2554_),
    .B(_2555_),
    .X(net282));
 sky130_fd_sc_hd__a22o_1 _4815_ (.A1(net1287),
    .A2(net1153),
    .B1(net1030),
    .B2(net817),
    .X(_2556_));
 sky130_fd_sc_hd__a22o_1 _4816_ (.A1(net1029),
    .A2(net760),
    .B1(net759),
    .B2(_2159_),
    .X(_2557_));
 sky130_fd_sc_hd__or2_1 _4817_ (.A(_2556_),
    .B(_2557_),
    .X(net283));
 sky130_fd_sc_hd__a22o_1 _4818_ (.A1(\u_reg.reg_rdata[27] ),
    .A2(net1153),
    .B1(net1026),
    .B2(net817),
    .X(_2558_));
 sky130_fd_sc_hd__a22o_1 _4819_ (.A1(net1024),
    .A2(net760),
    .B1(net756),
    .B2(_2164_),
    .X(_2559_));
 sky130_fd_sc_hd__or2_1 _4820_ (.A(_2558_),
    .B(_2559_),
    .X(net284));
 sky130_fd_sc_hd__a22o_1 _4821_ (.A1(\u_reg.reg_rdata[28] ),
    .A2(net1153),
    .B1(_2172_),
    .B2(net757),
    .X(_2560_));
 sky130_fd_sc_hd__a22o_1 _4822_ (.A1(net817),
    .A2(net1022),
    .B1(net1021),
    .B2(net761),
    .X(_2561_));
 sky130_fd_sc_hd__or2_1 _4823_ (.A(_2560_),
    .B(_2561_),
    .X(net285));
 sky130_fd_sc_hd__a22o_1 _4824_ (.A1(net1283),
    .A2(net1154),
    .B1(_2174_),
    .B2(net759),
    .X(_2562_));
 sky130_fd_sc_hd__a22o_1 _4825_ (.A1(net818),
    .A2(net1017),
    .B1(net1016),
    .B2(net760),
    .X(_2563_));
 sky130_fd_sc_hd__or2_1 _4826_ (.A(_2562_),
    .B(_2563_),
    .X(net286));
 sky130_fd_sc_hd__a22o_1 _4827_ (.A1(\u_reg.reg_rdata[30] ),
    .A2(net1153),
    .B1(_2179_),
    .B2(net756),
    .X(_2564_));
 sky130_fd_sc_hd__a22o_1 _4828_ (.A1(net818),
    .A2(net1013),
    .B1(net1012),
    .B2(net760),
    .X(_2565_));
 sky130_fd_sc_hd__or2_1 _4829_ (.A(_2564_),
    .B(_2565_),
    .X(net288));
 sky130_fd_sc_hd__a22o_1 _4830_ (.A1(net1280),
    .A2(net1153),
    .B1(net1010),
    .B2(net817),
    .X(_2566_));
 sky130_fd_sc_hd__a22o_1 _4831_ (.A1(net1009),
    .A2(net760),
    .B1(net756),
    .B2(_2187_),
    .X(_2567_));
 sky130_fd_sc_hd__or2_1 _4832_ (.A(_2566_),
    .B(_2567_),
    .X(net289));
 sky130_fd_sc_hd__mux4_1 _4833_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][1] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][1] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][1] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][1] ),
    .S0(net1397),
    .S1(net1390),
    .X(_2568_));
 sky130_fd_sc_hd__mux2_1 _4834_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[1] ),
    .A1(_2568_),
    .S(net1502),
    .X(_0010_));
 sky130_fd_sc_hd__mux4_1 _4835_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][2] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][2] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][2] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][2] ),
    .S0(net1396),
    .S1(net1391),
    .X(_2569_));
 sky130_fd_sc_hd__mux2_1 _4836_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[2] ),
    .A1(_2569_),
    .S(net1501),
    .X(_0011_));
 sky130_fd_sc_hd__mux4_1 _4837_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][3] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][3] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][3] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][3] ),
    .S0(net1398),
    .S1(net1391),
    .X(_2570_));
 sky130_fd_sc_hd__mux2_1 _4838_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[3] ),
    .A1(_2570_),
    .S(net1501),
    .X(_0012_));
 sky130_fd_sc_hd__mux4_2 _4839_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][4] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][4] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][4] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][4] ),
    .S0(net1398),
    .S1(net1391),
    .X(_2571_));
 sky130_fd_sc_hd__mux2_1 _4840_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[4] ),
    .A1(_2571_),
    .S(net1501),
    .X(_0013_));
 sky130_fd_sc_hd__mux4_2 _4841_ (.A0(net1815),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][5] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][5] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][5] ),
    .S0(net1392),
    .S1(net1385),
    .X(_2572_));
 sky130_fd_sc_hd__mux2_1 _4842_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[5] ),
    .A1(net1816),
    .S(net1501),
    .X(_0014_));
 sky130_fd_sc_hd__mux4_2 _4843_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][6] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][6] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][6] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][6] ),
    .S0(net1396),
    .S1(net1389),
    .X(_2573_));
 sky130_fd_sc_hd__mux2_1 _4844_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[6] ),
    .A1(_2573_),
    .S(net1501),
    .X(_0015_));
 sky130_fd_sc_hd__mux4_2 _4845_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][7] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][7] ),
    .A2(net1803),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][7] ),
    .S0(net1393),
    .S1(net1386),
    .X(_2574_));
 sky130_fd_sc_hd__mux2_1 _4846_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[7] ),
    .A1(net1804),
    .S(net1502),
    .X(_0016_));
 sky130_fd_sc_hd__mux4_2 _4847_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][8] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][8] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][8] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][8] ),
    .S0(net1394),
    .S1(net1387),
    .X(_2575_));
 sky130_fd_sc_hd__mux2_1 _4848_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[8] ),
    .A1(_2575_),
    .S(net1501),
    .X(_0017_));
 sky130_fd_sc_hd__mux4_2 _4849_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[0][9] ),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[1][9] ),
    .A2(\u_s2.u_sync_wbb.u_cmd_if.mem[2][9] ),
    .A3(\u_s2.u_sync_wbb.u_cmd_if.mem[3][9] ),
    .S0(net1396),
    .S1(net1389),
    .X(_2576_));
 sky130_fd_sc_hd__mux2_1 _4850_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[9] ),
    .A1(_2576_),
    .S(net1499),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _4851_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[14] ),
    .A1(_2329_),
    .S(net1496),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _4852_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[15] ),
    .A1(_2330_),
    .S(net1502),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _4853_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[16] ),
    .A1(_2331_),
    .S(net1500),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _4854_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[17] ),
    .A1(_2332_),
    .S(net1495),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _4855_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[18] ),
    .A1(_2333_),
    .S(net1499),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _4856_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[19] ),
    .A1(_2334_),
    .S(net1502),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _4857_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[20] ),
    .A1(_2335_),
    .S(net1500),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _4858_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[21] ),
    .A1(_2336_),
    .S(net1496),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _4859_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[22] ),
    .A1(_2337_),
    .S(net1502),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _4860_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[23] ),
    .A1(_2338_),
    .S(net1499),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _4861_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[24] ),
    .A1(_2339_),
    .S(net1497),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _4862_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[25] ),
    .A1(_2340_),
    .S(net1500),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _4863_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[26] ),
    .A1(_2341_),
    .S(net1496),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _4864_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[27] ),
    .A1(_2342_),
    .S(net1497),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _4865_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[28] ),
    .A1(_2343_),
    .S(net1501),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _4866_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[29] ),
    .A1(_2344_),
    .S(net1496),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _4867_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[30] ),
    .A1(_2345_),
    .S(net1496),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _4868_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[31] ),
    .A1(_2346_),
    .S(net1495),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _4869_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[32] ),
    .A1(_2347_),
    .S(net1497),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _4870_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[33] ),
    .A1(_2348_),
    .S(net1500),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _4871_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[34] ),
    .A1(_2349_),
    .S(net1499),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _4872_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[35] ),
    .A1(_2350_),
    .S(net1500),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _4873_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[36] ),
    .A1(_2351_),
    .S(net1500),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _4874_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[37] ),
    .A1(_2352_),
    .S(net1496),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _4875_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[38] ),
    .A1(_2353_),
    .S(net1500),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _4876_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[39] ),
    .A1(_2354_),
    .S(net1495),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _4877_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[40] ),
    .A1(_2355_),
    .S(net1498),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _4878_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[41] ),
    .A1(_2356_),
    .S(net1496),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _4879_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[42] ),
    .A1(_2357_),
    .S(net1495),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _4880_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[43] ),
    .A1(_2358_),
    .S(net1495),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _4881_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[44] ),
    .A1(_2359_),
    .S(net1500),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _4882_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[45] ),
    .A1(_2360_),
    .S(net1497),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _4883_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[46] ),
    .A1(_2361_),
    .S(net1495),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _4884_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[47] ),
    .A1(_2362_),
    .S(net1497),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _4885_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[48] ),
    .A1(_2363_),
    .S(net1496),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _4886_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[49] ),
    .A1(_2364_),
    .S(net1496),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _4887_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[50] ),
    .A1(_2004_),
    .S(net1499),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _4888_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[53] ),
    .A1(_2365_),
    .S(net1499),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _4889_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[54] ),
    .A1(_2366_),
    .S(net1496),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _4890_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[55] ),
    .A1(_2367_),
    .S(net1499),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _4891_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[56] ),
    .A1(_2368_),
    .S(net1495),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _4892_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[57] ),
    .A1(_2369_),
    .S(net1495),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _4893_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[58] ),
    .A1(_2370_),
    .S(net1495),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _4894_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[59] ),
    .A1(_2371_),
    .S(net1499),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _4895_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[60] ),
    .A1(net1789),
    .S(net1498),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _4896_ (.A0(\u_s2.u_sync_wbb.s_cmd_rd_data_l[61] ),
    .A1(net1786),
    .S(net1495),
    .X(_0064_));
 sky130_fd_sc_hd__a22o_1 _4897_ (.A1(net1180),
    .A2(_1964_),
    .B1(_1965_),
    .B2(net1409),
    .X(_2577_));
 sky130_fd_sc_hd__nand2_1 _4898_ (.A(net1407),
    .B(_1968_),
    .Y(_2578_));
 sky130_fd_sc_hd__or4b_4 _4899_ (.A(_1690_),
    .B(_1768_),
    .C(net1176),
    .D_N(_1760_),
    .X(_2579_));
 sky130_fd_sc_hd__a21oi_1 _4900_ (.A1(net1407),
    .A2(_1968_),
    .B1(_2579_),
    .Y(_2580_));
 sky130_fd_sc_hd__a21o_1 _4901_ (.A1(_1962_),
    .A2(_2577_),
    .B1(_2580_),
    .X(_2581_));
 sky130_fd_sc_hd__o21a_1 _4902_ (.A1(net1409),
    .A2(_1965_),
    .B1(net1224),
    .X(_2582_));
 sky130_fd_sc_hd__a31o_1 _4903_ (.A1(m3_wbd_stb_i),
    .A2(_1958_),
    .A3(_2582_),
    .B1(_2581_),
    .X(_2583_));
 sky130_fd_sc_hd__a21o_1 _4904_ (.A1(_1967_),
    .A2(_1970_),
    .B1(net1401),
    .X(_2584_));
 sky130_fd_sc_hd__mux2_1 _4905_ (.A0(net1409),
    .A1(_2583_),
    .S(_2584_),
    .X(_0065_));
 sky130_fd_sc_hd__o2bb2a_1 _4906_ (.A1_N(net1224),
    .A2_N(_1965_),
    .B1(_1962_),
    .B2(net1232),
    .X(_2585_));
 sky130_fd_sc_hd__a21o_1 _4907_ (.A1(_1964_),
    .A2(_2500_),
    .B1(_2585_),
    .X(_2586_));
 sky130_fd_sc_hd__and3_1 _4908_ (.A(_2578_),
    .B(_2579_),
    .C(_2586_),
    .X(_2587_));
 sky130_fd_sc_hd__mux2_1 _4909_ (.A0(net1407),
    .A1(_2587_),
    .S(_2584_),
    .X(_0066_));
 sky130_fd_sc_hd__nand2_1 _4910_ (.A(\u_s0.u_sync_wbb.m_state[1] ),
    .B(_1820_),
    .Y(_2588_));
 sky130_fd_sc_hd__nor2_4 _4911_ (.A(\u_s0.u_sync_wbb.m_state[1] ),
    .B(\u_s0.u_sync_wbb.m_state[2] ),
    .Y(_2589_));
 sky130_fd_sc_hd__or2_1 _4912_ (.A(\u_s0.u_sync_wbb.m_state[1] ),
    .B(\u_s0.u_sync_wbb.m_state[2] ),
    .X(_2590_));
 sky130_fd_sc_hd__nor2_1 _4913_ (.A(\u_s0.u_sync_wbb.m_state[0] ),
    .B(net1005),
    .Y(_2591_));
 sky130_fd_sc_hd__a221o_1 _4914_ (.A1(\u_s0.u_sync_wbb.m_state[1] ),
    .A2(_1820_),
    .B1(_1829_),
    .B2(net1005),
    .C1(_2591_),
    .X(_2592_));
 sky130_fd_sc_hd__a221o_2 _4915_ (.A1(\u_s0.u_sync_wbb.m_state[2] ),
    .A2(_1735_),
    .B1(_1784_),
    .B2(\u_s0.u_sync_wbb.m_state[0] ),
    .C1(_2592_),
    .X(_2593_));
 sky130_fd_sc_hd__nand2_1 _4916_ (.A(_1786_),
    .B(net580),
    .Y(_2594_));
 sky130_fd_sc_hd__o21a_1 _4917_ (.A1(_1786_),
    .A2(net580),
    .B1(_2589_),
    .X(_2595_));
 sky130_fd_sc_hd__a221o_1 _4918_ (.A1(\u_s0.u_sync_wbb.m_bl_cnt[0] ),
    .A2(net1005),
    .B1(_2594_),
    .B2(_2595_),
    .C1(net513),
    .X(_2596_));
 sky130_fd_sc_hd__a21bo_1 _4919_ (.A1(\u_s0.u_sync_wbb.m_bl_cnt[0] ),
    .A2(net513),
    .B1_N(_2596_),
    .X(_0067_));
 sky130_fd_sc_hd__o21ai_1 _4920_ (.A1(_1786_),
    .A2(net580),
    .B1(_1789_),
    .Y(_2597_));
 sky130_fd_sc_hd__or2_2 _4921_ (.A(_1786_),
    .B(_1789_),
    .X(_2598_));
 sky130_fd_sc_hd__o211a_1 _4922_ (.A1(net580),
    .A2(_2598_),
    .B1(_2597_),
    .C1(_2589_),
    .X(_2599_));
 sky130_fd_sc_hd__nand2_1 _4923_ (.A(\u_s0.u_sync_wbb.m_bl_cnt[0] ),
    .B(\u_s0.u_sync_wbb.m_bl_cnt[1] ),
    .Y(_2600_));
 sky130_fd_sc_hd__or2_1 _4924_ (.A(\u_s0.u_sync_wbb.m_bl_cnt[0] ),
    .B(\u_s0.u_sync_wbb.m_bl_cnt[1] ),
    .X(_2601_));
 sky130_fd_sc_hd__a31o_1 _4925_ (.A1(net1005),
    .A2(_2600_),
    .A3(_2601_),
    .B1(net513),
    .X(_2602_));
 sky130_fd_sc_hd__a2bb2o_1 _4926_ (.A1_N(_2599_),
    .A2_N(_2602_),
    .B1(\u_s0.u_sync_wbb.m_bl_cnt[1] ),
    .B2(net513),
    .X(_0068_));
 sky130_fd_sc_hd__o21ai_1 _4927_ (.A1(net580),
    .A2(_2598_),
    .B1(_1792_),
    .Y(_2603_));
 sky130_fd_sc_hd__or3_1 _4928_ (.A(_1792_),
    .B(net580),
    .C(_2598_),
    .X(_2604_));
 sky130_fd_sc_hd__and3_1 _4929_ (.A(_2589_),
    .B(_2603_),
    .C(_2604_),
    .X(_2605_));
 sky130_fd_sc_hd__nand2_1 _4930_ (.A(\u_s0.u_sync_wbb.m_bl_cnt[2] ),
    .B(_2601_),
    .Y(_2606_));
 sky130_fd_sc_hd__or3_1 _4931_ (.A(\u_s0.u_sync_wbb.m_bl_cnt[0] ),
    .B(\u_s0.u_sync_wbb.m_bl_cnt[1] ),
    .C(\u_s0.u_sync_wbb.m_bl_cnt[2] ),
    .X(_2607_));
 sky130_fd_sc_hd__a31o_1 _4932_ (.A1(net1005),
    .A2(_2606_),
    .A3(_2607_),
    .B1(net513),
    .X(_2608_));
 sky130_fd_sc_hd__a2bb2o_1 _4933_ (.A1_N(_2605_),
    .A2_N(_2608_),
    .B1(\u_s0.u_sync_wbb.m_bl_cnt[2] ),
    .B2(net513),
    .X(_0069_));
 sky130_fd_sc_hd__o31ai_1 _4934_ (.A1(_1792_),
    .A2(net580),
    .A3(_2598_),
    .B1(_1794_),
    .Y(_2609_));
 sky130_fd_sc_hd__o31a_1 _4935_ (.A1(_1795_),
    .A2(net580),
    .A3(_2598_),
    .B1(_2589_),
    .X(_2610_));
 sky130_fd_sc_hd__nand2_1 _4936_ (.A(\u_s0.u_sync_wbb.m_bl_cnt[3] ),
    .B(_2607_),
    .Y(_2611_));
 sky130_fd_sc_hd__or2_2 _4937_ (.A(\u_s0.u_sync_wbb.m_bl_cnt[3] ),
    .B(_2607_),
    .X(_2612_));
 sky130_fd_sc_hd__and3_1 _4938_ (.A(net1005),
    .B(_2611_),
    .C(_2612_),
    .X(_2613_));
 sky130_fd_sc_hd__a21oi_1 _4939_ (.A1(_2609_),
    .A2(_2610_),
    .B1(_2613_),
    .Y(_2614_));
 sky130_fd_sc_hd__mux2_1 _4940_ (.A0(_2614_),
    .A1(\u_s0.u_sync_wbb.m_bl_cnt[3] ),
    .S(net513),
    .X(_0070_));
 sky130_fd_sc_hd__o31a_1 _4941_ (.A1(_1795_),
    .A2(net581),
    .A3(_2598_),
    .B1(_1793_),
    .X(_2615_));
 sky130_fd_sc_hd__or3_4 _4942_ (.A(_1793_),
    .B(_1795_),
    .C(_2598_),
    .X(_2616_));
 sky130_fd_sc_hd__nor2_1 _4943_ (.A(net581),
    .B(_2616_),
    .Y(_2617_));
 sky130_fd_sc_hd__nor2_1 _4944_ (.A(\u_s0.u_sync_wbb.m_bl_cnt[4] ),
    .B(_2612_),
    .Y(_2618_));
 sky130_fd_sc_hd__a211o_1 _4945_ (.A1(\u_s0.u_sync_wbb.m_bl_cnt[4] ),
    .A2(_2612_),
    .B1(_2618_),
    .C1(_2589_),
    .X(_2619_));
 sky130_fd_sc_hd__o31a_1 _4946_ (.A1(net1005),
    .A2(_2615_),
    .A3(_2617_),
    .B1(_2619_),
    .X(_2620_));
 sky130_fd_sc_hd__mux2_1 _4947_ (.A0(_2620_),
    .A1(\u_s0.u_sync_wbb.m_bl_cnt[4] ),
    .S(net513),
    .X(_0071_));
 sky130_fd_sc_hd__or3_1 _4948_ (.A(net808),
    .B(net581),
    .C(_2616_),
    .X(_2621_));
 sky130_fd_sc_hd__o21ai_1 _4949_ (.A1(_1998_),
    .A2(_2616_),
    .B1(net808),
    .Y(_2622_));
 sky130_fd_sc_hd__and3_1 _4950_ (.A(_2589_),
    .B(_2621_),
    .C(_2622_),
    .X(_2623_));
 sky130_fd_sc_hd__o21ai_1 _4951_ (.A1(\u_s0.u_sync_wbb.m_bl_cnt[4] ),
    .A2(_2612_),
    .B1(\u_s0.u_sync_wbb.m_bl_cnt[5] ),
    .Y(_2624_));
 sky130_fd_sc_hd__or3_2 _4952_ (.A(\u_s0.u_sync_wbb.m_bl_cnt[5] ),
    .B(\u_s0.u_sync_wbb.m_bl_cnt[4] ),
    .C(_2612_),
    .X(_2625_));
 sky130_fd_sc_hd__a31o_1 _4953_ (.A1(net1006),
    .A2(_2624_),
    .A3(_2625_),
    .B1(net513),
    .X(_2626_));
 sky130_fd_sc_hd__a2bb2o_1 _4954_ (.A1_N(_2623_),
    .A2_N(_2626_),
    .B1(\u_s0.u_sync_wbb.m_bl_cnt[5] ),
    .B2(net513),
    .X(_0072_));
 sky130_fd_sc_hd__o31ai_1 _4955_ (.A1(net808),
    .A2(net581),
    .A3(_2616_),
    .B1(_1797_),
    .Y(_2627_));
 sky130_fd_sc_hd__or4_1 _4956_ (.A(_1797_),
    .B(net808),
    .C(net581),
    .D(_2616_),
    .X(_2628_));
 sky130_fd_sc_hd__and3_1 _4957_ (.A(_2589_),
    .B(_2627_),
    .C(_2628_),
    .X(_2629_));
 sky130_fd_sc_hd__or2_1 _4958_ (.A(\u_s0.u_sync_wbb.m_bl_cnt[6] ),
    .B(_2625_),
    .X(_2630_));
 sky130_fd_sc_hd__nand2_1 _4959_ (.A(\u_s0.u_sync_wbb.m_bl_cnt[6] ),
    .B(_2625_),
    .Y(_2631_));
 sky130_fd_sc_hd__a31o_1 _4960_ (.A1(net1005),
    .A2(_2630_),
    .A3(_2631_),
    .B1(net514),
    .X(_2632_));
 sky130_fd_sc_hd__a2bb2o_1 _4961_ (.A1_N(_2629_),
    .A2_N(_2632_),
    .B1(\u_s0.u_sync_wbb.m_bl_cnt[6] ),
    .B2(net514),
    .X(_0073_));
 sky130_fd_sc_hd__o41a_1 _4962_ (.A1(_1797_),
    .A2(net808),
    .A3(net581),
    .A4(_2616_),
    .B1(_1796_),
    .X(_2633_));
 sky130_fd_sc_hd__nor4_1 _4963_ (.A(_1798_),
    .B(_1800_),
    .C(net581),
    .D(_2616_),
    .Y(_2634_));
 sky130_fd_sc_hd__or4_1 _4964_ (.A(_1798_),
    .B(_1800_),
    .C(net581),
    .D(_2616_),
    .X(_2635_));
 sky130_fd_sc_hd__nor2_1 _4965_ (.A(\u_s0.u_sync_wbb.m_bl_cnt[7] ),
    .B(_2630_),
    .Y(_2636_));
 sky130_fd_sc_hd__a21o_1 _4966_ (.A1(\u_s0.u_sync_wbb.m_bl_cnt[7] ),
    .A2(_2630_),
    .B1(_2589_),
    .X(_2637_));
 sky130_fd_sc_hd__o32a_1 _4967_ (.A1(net1005),
    .A2(_2633_),
    .A3(_2634_),
    .B1(_2636_),
    .B2(_2637_),
    .X(_2638_));
 sky130_fd_sc_hd__mux2_1 _4968_ (.A0(_2638_),
    .A1(\u_s0.u_sync_wbb.m_bl_cnt[7] ),
    .S(net514),
    .X(_0074_));
 sky130_fd_sc_hd__a221o_1 _4969_ (.A1(_1801_),
    .A2(_2617_),
    .B1(_2635_),
    .B2(_1799_),
    .C1(net1006),
    .X(_2639_));
 sky130_fd_sc_hd__or3_1 _4970_ (.A(\u_s0.u_sync_wbb.m_bl_cnt[7] ),
    .B(\u_s0.u_sync_wbb.m_bl_cnt[8] ),
    .C(_2630_),
    .X(_2640_));
 sky130_fd_sc_hd__a21oi_1 _4971_ (.A1(net1006),
    .A2(_2640_),
    .B1(net514),
    .Y(_2641_));
 sky130_fd_sc_hd__o21ai_1 _4972_ (.A1(\u_s0.u_sync_wbb.m_bl_cnt[7] ),
    .A2(_2630_),
    .B1(\u_s0.u_sync_wbb.m_bl_cnt[8] ),
    .Y(_2642_));
 sky130_fd_sc_hd__a31oi_1 _4973_ (.A1(net1006),
    .A2(_2640_),
    .A3(_2642_),
    .B1(net514),
    .Y(_2643_));
 sky130_fd_sc_hd__a22o_1 _4974_ (.A1(\u_s0.u_sync_wbb.m_bl_cnt[8] ),
    .A2(net514),
    .B1(_2639_),
    .B2(_2643_),
    .X(_0075_));
 sky130_fd_sc_hd__o31a_1 _4975_ (.A1(_1802_),
    .A2(_1998_),
    .A3(_2616_),
    .B1(_1787_),
    .X(_2644_));
 sky130_fd_sc_hd__nor4_1 _4976_ (.A(_1787_),
    .B(_1802_),
    .C(net581),
    .D(_2616_),
    .Y(_2645_));
 sky130_fd_sc_hd__or3b_1 _4977_ (.A(_2589_),
    .B(_2640_),
    .C_N(\u_s0.u_sync_wbb.m_bl_cnt[9] ),
    .X(_2646_));
 sky130_fd_sc_hd__o31a_1 _4978_ (.A1(net1006),
    .A2(_2644_),
    .A3(_2645_),
    .B1(_2646_),
    .X(_2647_));
 sky130_fd_sc_hd__o22a_1 _4979_ (.A1(\u_s0.u_sync_wbb.m_bl_cnt[9] ),
    .A2(_2641_),
    .B1(_2647_),
    .B2(net514),
    .X(_0076_));
 sky130_fd_sc_hd__nor2_2 _4980_ (.A(net1223),
    .B(net1275),
    .Y(_2648_));
 sky130_fd_sc_hd__and3b_1 _4981_ (.A_N(net1275),
    .B(m1_wbd_adr_i[3]),
    .C(net1276),
    .X(_2649_));
 sky130_fd_sc_hd__and3_1 _4982_ (.A(net1276),
    .B(net1275),
    .C(m3_wbd_adr_i[3]),
    .X(_2650_));
 sky130_fd_sc_hd__and2b_1 _4983_ (.A_N(net1276),
    .B(m2_wbd_adr_i[3]),
    .X(_2651_));
 sky130_fd_sc_hd__or3_1 _4984_ (.A(net1276),
    .B(\u_wbi_arb.gnt[1] ),
    .C(net1597),
    .X(_2652_));
 sky130_fd_sc_hd__o41a_4 _4985_ (.A1(_2019_),
    .A2(_2649_),
    .A3(_2650_),
    .A4(_2651_),
    .B1(_2652_),
    .X(_2653_));
 sky130_fd_sc_hd__and3_1 _4986_ (.A(net1219),
    .B(net1274),
    .C(m2_wbd_adr_i[4]),
    .X(_2654_));
 sky130_fd_sc_hd__a221o_1 _4987_ (.A1(net1210),
    .A2(m1_wbd_adr_i[4]),
    .B1(_2013_),
    .B2(m3_wbd_adr_i[4]),
    .C1(_2019_),
    .X(_2655_));
 sky130_fd_sc_hd__o22ai_4 _4988_ (.A1(net1596),
    .A2(net1148),
    .B1(_2654_),
    .B2(_2655_),
    .Y(_2656_));
 sky130_fd_sc_hd__nand3b_2 _4989_ (.A_N(net1274),
    .B(m1_wbd_adr_i[2]),
    .C(net1277),
    .Y(_2657_));
 sky130_fd_sc_hd__nand3_2 _4990_ (.A(net1277),
    .B(net1274),
    .C(m3_wbd_adr_i[2]),
    .Y(_2658_));
 sky130_fd_sc_hd__nand2b_1 _4991_ (.A_N(net1277),
    .B(m2_wbd_adr_i[2]),
    .Y(_2659_));
 sky130_fd_sc_hd__nor3_2 _4992_ (.A(net1276),
    .B(net1274),
    .C(net1598),
    .Y(_2660_));
 sky130_fd_sc_hd__a41oi_4 _4993_ (.A1(net1152),
    .A2(_2657_),
    .A3(_2658_),
    .A4(_2659_),
    .B1(_2660_),
    .Y(_2661_));
 sky130_fd_sc_hd__a41o_4 _4994_ (.A1(net1152),
    .A2(_2657_),
    .A3(_2658_),
    .A4(_2659_),
    .B1(_2660_),
    .X(_2662_));
 sky130_fd_sc_hd__nor3_1 _4995_ (.A(_2653_),
    .B(_2656_),
    .C(_2662_),
    .Y(_2663_));
 sky130_fd_sc_hd__mux4_2 _4996_ (.A0(m0_wbd_we_i),
    .A1(m1_wbd_we_i),
    .A2(m2_wbd_we_i),
    .A3(m3_wbd_we_i),
    .S0(net1276),
    .S1(net1274),
    .X(_2664_));
 sky130_fd_sc_hd__nand2b_1 _4997_ (.A_N(net711),
    .B(_2664_),
    .Y(_2665_));
 sky130_fd_sc_hd__and2_1 _4998_ (.A(m1_wbd_sel_i[2]),
    .B(_2648_),
    .X(_2666_));
 sky130_fd_sc_hd__a221o_1 _4999_ (.A1(net1219),
    .A2(m2_wbd_sel_i[2]),
    .B1(_2013_),
    .B2(m3_wbd_sel_i[2]),
    .C1(_2019_),
    .X(_2667_));
 sky130_fd_sc_hd__o22a_1 _5000_ (.A1(m0_wbd_sel_i[2]),
    .A2(net1148),
    .B1(_2666_),
    .B2(_2667_),
    .X(_2668_));
 sky130_fd_sc_hd__and4b_4 _5001_ (.A_N(net711),
    .B(net621),
    .C(_2664_),
    .D(net617),
    .X(_2669_));
 sky130_fd_sc_hd__or2_1 _5002_ (.A(net1586),
    .B(net1149),
    .X(_2670_));
 sky130_fd_sc_hd__a21o_1 _5003_ (.A1(net1215),
    .A2(net1555),
    .B1(net1220),
    .X(_2671_));
 sky130_fd_sc_hd__o211a_1 _5004_ (.A1(net1216),
    .A2(net1529),
    .B1(_2670_),
    .C1(_2671_),
    .X(_2672_));
 sky130_fd_sc_hd__mux2_1 _5005_ (.A0(\u_reg.reg_5[16] ),
    .A1(net708),
    .S(net561),
    .X(_0077_));
 sky130_fd_sc_hd__or2_1 _5006_ (.A(net1585),
    .B(net1150),
    .X(_2673_));
 sky130_fd_sc_hd__a21o_1 _5007_ (.A1(net1216),
    .A2(net1554),
    .B1(net1220),
    .X(_2674_));
 sky130_fd_sc_hd__o211a_1 _5008_ (.A1(net1216),
    .A2(net1528),
    .B1(_2673_),
    .C1(_2674_),
    .X(_2675_));
 sky130_fd_sc_hd__mux2_1 _5009_ (.A0(\u_reg.reg_5[17] ),
    .A1(net707),
    .S(net561),
    .X(_0078_));
 sky130_fd_sc_hd__or2_1 _5010_ (.A(net1584),
    .B(net1152),
    .X(_2676_));
 sky130_fd_sc_hd__a21o_1 _5011_ (.A1(net1222),
    .A2(m2_wbd_dat_i[18]),
    .B1(net1211),
    .X(_2677_));
 sky130_fd_sc_hd__o211a_4 _5012_ (.A1(net1222),
    .A2(net1553),
    .B1(_2676_),
    .C1(_2677_),
    .X(_2678_));
 sky130_fd_sc_hd__mux2_1 _5013_ (.A0(\u_reg.reg_5[18] ),
    .A1(_2678_),
    .S(_2669_),
    .X(_0079_));
 sky130_fd_sc_hd__or2_1 _5014_ (.A(net1583),
    .B(net1149),
    .X(_2679_));
 sky130_fd_sc_hd__a21o_1 _5015_ (.A1(net1221),
    .A2(net1527),
    .B1(net1213),
    .X(_2680_));
 sky130_fd_sc_hd__o211a_2 _5016_ (.A1(net1221),
    .A2(net1552),
    .B1(_2679_),
    .C1(_2680_),
    .X(_2681_));
 sky130_fd_sc_hd__mux2_1 _5017_ (.A0(\u_reg.reg_5[19] ),
    .A1(_2681_),
    .S(_2669_),
    .X(_0080_));
 sky130_fd_sc_hd__or2_1 _5018_ (.A(net1581),
    .B(net1149),
    .X(_2682_));
 sky130_fd_sc_hd__a21o_1 _5019_ (.A1(net1213),
    .A2(net1550),
    .B1(net1221),
    .X(_2683_));
 sky130_fd_sc_hd__o211a_1 _5020_ (.A1(net1213),
    .A2(net1526),
    .B1(_2682_),
    .C1(_2683_),
    .X(_2684_));
 sky130_fd_sc_hd__mux2_1 _5021_ (.A0(\u_reg.reg_5[20] ),
    .A1(net706),
    .S(net561),
    .X(_0081_));
 sky130_fd_sc_hd__a21o_1 _5022_ (.A1(net1211),
    .A2(net1549),
    .B1(net1222),
    .X(_2685_));
 sky130_fd_sc_hd__o221a_1 _5023_ (.A1(net1211),
    .A2(net1525),
    .B1(net1580),
    .B2(net1151),
    .C1(_2685_),
    .X(_2686_));
 sky130_fd_sc_hd__mux2_1 _5024_ (.A0(\u_reg.reg_5[21] ),
    .A1(net705),
    .S(net561),
    .X(_0082_));
 sky130_fd_sc_hd__a21o_1 _5025_ (.A1(net1211),
    .A2(net1548),
    .B1(net1222),
    .X(_2687_));
 sky130_fd_sc_hd__o221a_4 _5026_ (.A1(net1211),
    .A2(net2051),
    .B1(net1579),
    .B2(net1151),
    .C1(_2687_),
    .X(_2688_));
 sky130_fd_sc_hd__mux2_1 _5027_ (.A0(\u_reg.reg_5[22] ),
    .A1(_2688_),
    .S(_2669_),
    .X(_0083_));
 sky130_fd_sc_hd__a21o_1 _5028_ (.A1(net1212),
    .A2(net1547),
    .B1(net1222),
    .X(_2689_));
 sky130_fd_sc_hd__o221a_1 _5029_ (.A1(net1212),
    .A2(net1524),
    .B1(net1578),
    .B2(net1151),
    .C1(_2689_),
    .X(_2690_));
 sky130_fd_sc_hd__mux2_1 _5030_ (.A0(\u_reg.reg_5[23] ),
    .A1(net704),
    .S(_2669_),
    .X(_0084_));
 sky130_fd_sc_hd__nor3b_1 _5031_ (.A(_2661_),
    .B(_2656_),
    .C_N(_2653_),
    .Y(_2691_));
 sky130_fd_sc_hd__and3_1 _5032_ (.A(net1276),
    .B(net1274),
    .C(m3_wbd_sel_i[0]),
    .X(_2692_));
 sky130_fd_sc_hd__a221o_1 _5033_ (.A1(net1219),
    .A2(m2_wbd_sel_i[0]),
    .B1(m1_wbd_sel_i[0]),
    .B2(_2648_),
    .C1(_2019_),
    .X(_2693_));
 sky130_fd_sc_hd__o22a_4 _5034_ (.A1(net1565),
    .A2(net1148),
    .B1(_2692_),
    .B2(_2693_),
    .X(_2694_));
 sky130_fd_sc_hd__and3b_4 _5035_ (.A_N(net618),
    .B(net610),
    .C(_2694_),
    .X(_2695_));
 sky130_fd_sc_hd__a21o_1 _5036_ (.A1(net1211),
    .A2(net1562),
    .B1(net1222),
    .X(_2696_));
 sky130_fd_sc_hd__o221a_4 _5037_ (.A1(net1211),
    .A2(net2050),
    .B1(net1593),
    .B2(net1148),
    .C1(_2696_),
    .X(_2697_));
 sky130_fd_sc_hd__mux2_1 _5038_ (.A0(\u_reg.reg_6[0] ),
    .A1(_2697_),
    .S(_2695_),
    .X(_0085_));
 sky130_fd_sc_hd__or2_1 _5039_ (.A(net1582),
    .B(net1152),
    .X(_2698_));
 sky130_fd_sc_hd__a21o_1 _5040_ (.A1(net1218),
    .A2(net1551),
    .B1(net1223),
    .X(_2699_));
 sky130_fd_sc_hd__o211a_2 _5041_ (.A1(net1218),
    .A2(m2_wbd_dat_i[1]),
    .B1(_2698_),
    .C1(_2699_),
    .X(_2700_));
 sky130_fd_sc_hd__mux2_1 _5042_ (.A0(\u_reg.reg_6[1] ),
    .A1(_2700_),
    .S(_2695_),
    .X(_0086_));
 sky130_fd_sc_hd__or2_1 _5043_ (.A(net1574),
    .B(net1151),
    .X(_2701_));
 sky130_fd_sc_hd__a21o_1 _5044_ (.A1(net1211),
    .A2(net1543),
    .B1(net1222),
    .X(_2702_));
 sky130_fd_sc_hd__o211a_2 _5045_ (.A1(net1211),
    .A2(m2_wbd_dat_i[2]),
    .B1(_2701_),
    .C1(_2702_),
    .X(_2703_));
 sky130_fd_sc_hd__mux2_1 _5046_ (.A0(\u_reg.reg_6[2] ),
    .A1(_2703_),
    .S(_2695_),
    .X(_0087_));
 sky130_fd_sc_hd__a21o_1 _5047_ (.A1(net1210),
    .A2(m1_wbd_dat_i[3]),
    .B1(net1219),
    .X(_2704_));
 sky130_fd_sc_hd__o221a_4 _5048_ (.A1(net1210),
    .A2(net2088),
    .B1(m0_wbd_dat_i[3]),
    .B2(net1148),
    .C1(_2704_),
    .X(_2705_));
 sky130_fd_sc_hd__mux2_1 _5049_ (.A0(\u_reg.reg_6[3] ),
    .A1(_2705_),
    .S(_2695_),
    .X(_0088_));
 sky130_fd_sc_hd__a21o_1 _5050_ (.A1(net1213),
    .A2(net1540),
    .B1(net1221),
    .X(_2706_));
 sky130_fd_sc_hd__o221a_4 _5051_ (.A1(net1213),
    .A2(net1518),
    .B1(net1571),
    .B2(net1149),
    .C1(_2706_),
    .X(_2707_));
 sky130_fd_sc_hd__mux2_1 _5052_ (.A0(\u_reg.reg_6[4] ),
    .A1(_2707_),
    .S(_2695_),
    .X(_0089_));
 sky130_fd_sc_hd__a21o_1 _5053_ (.A1(net1213),
    .A2(net1539),
    .B1(net1221),
    .X(_2708_));
 sky130_fd_sc_hd__o221a_4 _5054_ (.A1(net1213),
    .A2(net1517),
    .B1(net1570),
    .B2(net1149),
    .C1(_2708_),
    .X(_2709_));
 sky130_fd_sc_hd__mux2_1 _5055_ (.A0(\u_reg.reg_6[5] ),
    .A1(_2709_),
    .S(_2695_),
    .X(_0090_));
 sky130_fd_sc_hd__or2_1 _5056_ (.A(net1569),
    .B(net1150),
    .X(_2710_));
 sky130_fd_sc_hd__a21o_1 _5057_ (.A1(net1217),
    .A2(net1538),
    .B1(net1220),
    .X(_2711_));
 sky130_fd_sc_hd__o211a_2 _5058_ (.A1(net1217),
    .A2(net1516),
    .B1(_2710_),
    .C1(_2711_),
    .X(_2712_));
 sky130_fd_sc_hd__mux2_1 _5059_ (.A0(\u_reg.reg_6[6] ),
    .A1(_2712_),
    .S(_2695_),
    .X(_0091_));
 sky130_fd_sc_hd__a21o_1 _5060_ (.A1(net1215),
    .A2(net1537),
    .B1(net1220),
    .X(_2713_));
 sky130_fd_sc_hd__o221a_4 _5061_ (.A1(net1215),
    .A2(net1515),
    .B1(net1568),
    .B2(net1149),
    .C1(_2713_),
    .X(_2714_));
 sky130_fd_sc_hd__mux2_1 _5062_ (.A0(\u_reg.reg_6[7] ),
    .A1(_2714_),
    .S(_2695_),
    .X(_0092_));
 sky130_fd_sc_hd__and3_1 _5063_ (.A(net1276),
    .B(net1274),
    .C(m3_wbd_sel_i[1]),
    .X(_2715_));
 sky130_fd_sc_hd__a221o_1 _5064_ (.A1(net1219),
    .A2(m2_wbd_sel_i[1]),
    .B1(m1_wbd_sel_i[1]),
    .B2(_2648_),
    .C1(_2019_),
    .X(_2716_));
 sky130_fd_sc_hd__o22a_1 _5065_ (.A1(m0_wbd_sel_i[1]),
    .A2(net1148),
    .B1(_2715_),
    .B2(_2716_),
    .X(_2717_));
 sky130_fd_sc_hd__and3b_4 _5066_ (.A_N(net619),
    .B(net611),
    .C(net609),
    .X(_2718_));
 sky130_fd_sc_hd__or2_1 _5067_ (.A(net1567),
    .B(net1150),
    .X(_2719_));
 sky130_fd_sc_hd__a21o_1 _5068_ (.A1(net1220),
    .A2(net1514),
    .B1(net1215),
    .X(_2720_));
 sky130_fd_sc_hd__o211a_4 _5069_ (.A1(net1220),
    .A2(net1536),
    .B1(_2719_),
    .C1(_2720_),
    .X(_2721_));
 sky130_fd_sc_hd__mux2_1 _5070_ (.A0(\u_reg.reg_6[8] ),
    .A1(_2721_),
    .S(_2718_),
    .X(_0093_));
 sky130_fd_sc_hd__a21o_1 _5071_ (.A1(net1215),
    .A2(net1535),
    .B1(net1223),
    .X(_2722_));
 sky130_fd_sc_hd__o221a_4 _5072_ (.A1(net1215),
    .A2(net1513),
    .B1(net1566),
    .B2(net1150),
    .C1(_2722_),
    .X(_2723_));
 sky130_fd_sc_hd__mux2_1 _5073_ (.A0(\u_reg.reg_6[9] ),
    .A1(_2723_),
    .S(_2718_),
    .X(_0094_));
 sky130_fd_sc_hd__a21o_1 _5074_ (.A1(net1214),
    .A2(net1561),
    .B1(net1220),
    .X(_2724_));
 sky130_fd_sc_hd__o221a_4 _5075_ (.A1(net1213),
    .A2(net1534),
    .B1(net1592),
    .B2(net1149),
    .C1(_2724_),
    .X(_2725_));
 sky130_fd_sc_hd__mux2_1 _5076_ (.A0(\u_reg.reg_6[10] ),
    .A1(_2725_),
    .S(_2718_),
    .X(_0095_));
 sky130_fd_sc_hd__a21o_1 _5077_ (.A1(net1214),
    .A2(net1560),
    .B1(net1221),
    .X(_2726_));
 sky130_fd_sc_hd__o221a_1 _5078_ (.A1(net1213),
    .A2(net1533),
    .B1(net1591),
    .B2(net1149),
    .C1(_2726_),
    .X(_2727_));
 sky130_fd_sc_hd__mux2_1 _5079_ (.A0(\u_reg.reg_6[11] ),
    .A1(net702),
    .S(_2718_),
    .X(_0096_));
 sky130_fd_sc_hd__a21o_1 _5080_ (.A1(net1216),
    .A2(net1559),
    .B1(net1220),
    .X(_2728_));
 sky130_fd_sc_hd__o221a_1 _5081_ (.A1(net1216),
    .A2(net1532),
    .B1(net1590),
    .B2(net1150),
    .C1(_2728_),
    .X(_2729_));
 sky130_fd_sc_hd__mux2_1 _5082_ (.A0(\u_reg.reg_6[12] ),
    .A1(net701),
    .S(_2718_),
    .X(_0097_));
 sky130_fd_sc_hd__a21o_1 _5083_ (.A1(net1212),
    .A2(net1558),
    .B1(net1222),
    .X(_2730_));
 sky130_fd_sc_hd__o221a_1 _5084_ (.A1(net1212),
    .A2(m2_wbd_dat_i[13]),
    .B1(net1589),
    .B2(net1151),
    .C1(_2730_),
    .X(_2731_));
 sky130_fd_sc_hd__mux2_1 _5085_ (.A0(\u_reg.reg_6[13] ),
    .A1(net700),
    .S(_2718_),
    .X(_0098_));
 sky130_fd_sc_hd__a21o_1 _5086_ (.A1(net1212),
    .A2(net1557),
    .B1(net1222),
    .X(_2732_));
 sky130_fd_sc_hd__o221a_2 _5087_ (.A1(net1212),
    .A2(net1531),
    .B1(net1588),
    .B2(net1151),
    .C1(_2732_),
    .X(_2733_));
 sky130_fd_sc_hd__mux2_1 _5088_ (.A0(\u_reg.reg_6[14] ),
    .A1(net699),
    .S(_2718_),
    .X(_0099_));
 sky130_fd_sc_hd__a21o_1 _5089_ (.A1(net1212),
    .A2(net1556),
    .B1(net1222),
    .X(_2734_));
 sky130_fd_sc_hd__o221a_1 _5090_ (.A1(net1212),
    .A2(net1530),
    .B1(net1587),
    .B2(net1151),
    .C1(_2734_),
    .X(_2735_));
 sky130_fd_sc_hd__mux2_1 _5091_ (.A0(\u_reg.reg_6[15] ),
    .A1(net697),
    .S(_2718_),
    .X(_0100_));
 sky130_fd_sc_hd__and3b_2 _5092_ (.A_N(net620),
    .B(net617),
    .C(net616),
    .X(_2736_));
 sky130_fd_sc_hd__mux2_1 _5093_ (.A0(\u_reg.reg_6[16] ),
    .A1(net708),
    .S(net560),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _5094_ (.A0(\u_reg.reg_6[17] ),
    .A1(net707),
    .S(net560),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _5095_ (.A0(\u_reg.reg_6[18] ),
    .A1(_2678_),
    .S(_2736_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _5096_ (.A0(\u_reg.reg_6[19] ),
    .A1(_2681_),
    .S(_2736_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _5097_ (.A0(\u_reg.reg_6[20] ),
    .A1(net706),
    .S(net560),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _5098_ (.A0(\u_reg.reg_6[21] ),
    .A1(net705),
    .S(net560),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _5099_ (.A0(\u_reg.reg_6[22] ),
    .A1(_2688_),
    .S(_2736_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _5100_ (.A0(\u_reg.reg_6[23] ),
    .A1(net704),
    .S(net560),
    .X(_0108_));
 sky130_fd_sc_hd__nand2_1 _5101_ (.A(_2653_),
    .B(_2661_),
    .Y(_2737_));
 sky130_fd_sc_hd__nor2_1 _5102_ (.A(_2656_),
    .B(_2737_),
    .Y(_2738_));
 sky130_fd_sc_hd__and3b_4 _5103_ (.A_N(net618),
    .B(_2694_),
    .C(net603),
    .X(_2739_));
 sky130_fd_sc_hd__mux2_1 _5104_ (.A0(\u_reg.reg_7[0] ),
    .A1(_2697_),
    .S(_2739_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _5105_ (.A0(\u_reg.reg_7[1] ),
    .A1(_2700_),
    .S(_2739_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _5106_ (.A0(\u_reg.reg_7[2] ),
    .A1(_2703_),
    .S(_2739_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _5107_ (.A0(\u_reg.reg_7[3] ),
    .A1(_2705_),
    .S(_2739_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _5108_ (.A0(\u_reg.reg_7[4] ),
    .A1(_2707_),
    .S(_2739_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _5109_ (.A0(\u_reg.reg_7[5] ),
    .A1(_2709_),
    .S(_2739_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _5110_ (.A0(\u_reg.reg_7[6] ),
    .A1(_2712_),
    .S(_2739_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _5111_ (.A0(\u_reg.reg_7[7] ),
    .A1(_2714_),
    .S(_2739_),
    .X(_0116_));
 sky130_fd_sc_hd__and3b_4 _5112_ (.A_N(net620),
    .B(net609),
    .C(net608),
    .X(_2740_));
 sky130_fd_sc_hd__mux2_1 _5113_ (.A0(\u_reg.reg_7[8] ),
    .A1(_2721_),
    .S(_2740_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _5114_ (.A0(\u_reg.reg_7[9] ),
    .A1(net703),
    .S(net559),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _5115_ (.A0(\u_reg.reg_7[10] ),
    .A1(_2725_),
    .S(_2740_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _5116_ (.A0(\u_reg.reg_7[11] ),
    .A1(net702),
    .S(net559),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _5117_ (.A0(\u_reg.reg_7[12] ),
    .A1(net701),
    .S(net559),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _5118_ (.A0(\u_reg.reg_7[13] ),
    .A1(net700),
    .S(_2740_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _5119_ (.A0(\u_reg.reg_7[14] ),
    .A1(net699),
    .S(net559),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _5120_ (.A0(\u_reg.reg_7[15] ),
    .A1(net697),
    .S(net559),
    .X(_0124_));
 sky130_fd_sc_hd__and3b_2 _5121_ (.A_N(net618),
    .B(net617),
    .C(net603),
    .X(_2741_));
 sky130_fd_sc_hd__mux2_1 _5122_ (.A0(\u_reg.reg_7[16] ),
    .A1(net708),
    .S(net558),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _5123_ (.A0(\u_reg.reg_7[17] ),
    .A1(net707),
    .S(net558),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _5124_ (.A0(\u_reg.reg_7[18] ),
    .A1(_2678_),
    .S(_2741_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _5125_ (.A0(\u_reg.reg_7[19] ),
    .A1(_2681_),
    .S(_2741_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _5126_ (.A0(\u_reg.reg_7[20] ),
    .A1(net706),
    .S(net558),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _5127_ (.A0(\u_reg.reg_7[21] ),
    .A1(net705),
    .S(net558),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _5128_ (.A0(\u_reg.reg_7[22] ),
    .A1(_2688_),
    .S(_2741_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _5129_ (.A0(\u_reg.reg_7[23] ),
    .A1(net704),
    .S(net558),
    .X(_0132_));
 sky130_fd_sc_hd__and4b_1 _5130_ (.A_N(net711),
    .B(net622),
    .C(_2664_),
    .D(net609),
    .X(_2742_));
 sky130_fd_sc_hd__mux2_1 _5131_ (.A0(\u_reg.reg_5[8] ),
    .A1(_2721_),
    .S(_2742_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _5132_ (.A0(\u_reg.reg_5[9] ),
    .A1(_2723_),
    .S(net557),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _5133_ (.A0(\u_reg.reg_5[10] ),
    .A1(_2725_),
    .S(net557),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _5134_ (.A0(\u_reg.reg_5[11] ),
    .A1(net702),
    .S(net557),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _5135_ (.A0(\u_reg.reg_5[12] ),
    .A1(net701),
    .S(net557),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _5136_ (.A0(\u_reg.reg_5[13] ),
    .A1(net700),
    .S(net557),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _5137_ (.A0(\u_reg.reg_5[14] ),
    .A1(net699),
    .S(net557),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _5138_ (.A0(\u_reg.reg_5[15] ),
    .A1(net697),
    .S(net557),
    .X(_0140_));
 sky130_fd_sc_hd__and4b_1 _5139_ (.A_N(net711),
    .B(net621),
    .C(_2664_),
    .D(_2694_),
    .X(_2743_));
 sky130_fd_sc_hd__mux2_1 _5140_ (.A0(\u_reg.reg_5[0] ),
    .A1(_2697_),
    .S(net556),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _5141_ (.A0(\u_reg.reg_5[1] ),
    .A1(_2700_),
    .S(net556),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _5142_ (.A0(\u_reg.reg_5[2] ),
    .A1(_2703_),
    .S(_2743_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _5143_ (.A0(\u_reg.reg_5[3] ),
    .A1(_2705_),
    .S(_2743_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _5144_ (.A0(\u_reg.reg_5[4] ),
    .A1(_2707_),
    .S(net556),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _5145_ (.A0(\u_reg.reg_5[5] ),
    .A1(_2709_),
    .S(net556),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _5146_ (.A0(\u_reg.reg_5[6] ),
    .A1(_2712_),
    .S(net556),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _5147_ (.A0(\u_reg.reg_5[7] ),
    .A1(_2714_),
    .S(net556),
    .X(_0148_));
 sky130_fd_sc_hd__nor3_2 _5148_ (.A(_2653_),
    .B(_2656_),
    .C(_2661_),
    .Y(_2744_));
 sky130_fd_sc_hd__and3b_4 _5149_ (.A_N(net618),
    .B(net617),
    .C(net598),
    .X(_2745_));
 sky130_fd_sc_hd__mux2_1 _5150_ (.A0(\u_reg.reg_4[16] ),
    .A1(net708),
    .S(net555),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _5151_ (.A0(\u_reg.reg_4[17] ),
    .A1(net707),
    .S(net555),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _5152_ (.A0(\u_reg.reg_4[18] ),
    .A1(_2678_),
    .S(_2745_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _5153_ (.A0(\u_reg.reg_4[19] ),
    .A1(_2681_),
    .S(_2745_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _5154_ (.A0(\u_reg.reg_4[20] ),
    .A1(net706),
    .S(net555),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _5155_ (.A0(\u_reg.reg_4[21] ),
    .A1(net705),
    .S(net555),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _5156_ (.A0(\u_reg.reg_4[22] ),
    .A1(_2688_),
    .S(_2745_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _5157_ (.A0(\u_reg.reg_4[23] ),
    .A1(net704),
    .S(_2745_),
    .X(_0156_));
 sky130_fd_sc_hd__and3b_4 _5158_ (.A_N(net619),
    .B(net609),
    .C(net599),
    .X(_2746_));
 sky130_fd_sc_hd__mux2_1 _5159_ (.A0(\u_reg.reg_4[8] ),
    .A1(_2721_),
    .S(_2746_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _5160_ (.A0(\u_reg.reg_4[9] ),
    .A1(net703),
    .S(net554),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _5161_ (.A0(\u_reg.reg_4[10] ),
    .A1(_2725_),
    .S(_2746_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _5162_ (.A0(\u_reg.reg_4[11] ),
    .A1(net702),
    .S(net554),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _5163_ (.A0(\u_reg.reg_4[12] ),
    .A1(net701),
    .S(net554),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _5164_ (.A0(\u_reg.reg_4[13] ),
    .A1(net700),
    .S(_2746_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _5165_ (.A0(\u_reg.reg_4[14] ),
    .A1(net699),
    .S(net554),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _5166_ (.A0(\u_reg.reg_4[15] ),
    .A1(net697),
    .S(net554),
    .X(_0164_));
 sky130_fd_sc_hd__and3b_4 _5167_ (.A_N(net618),
    .B(_2694_),
    .C(net598),
    .X(_2747_));
 sky130_fd_sc_hd__mux2_1 _5168_ (.A0(\u_reg.reg_4[0] ),
    .A1(_2697_),
    .S(_2747_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _5169_ (.A0(\u_reg.reg_4[1] ),
    .A1(_2700_),
    .S(_2747_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _5170_ (.A0(\u_reg.reg_4[2] ),
    .A1(_2703_),
    .S(_2747_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _5171_ (.A0(\u_reg.reg_4[3] ),
    .A1(_2705_),
    .S(_2747_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _5172_ (.A0(\u_reg.reg_4[4] ),
    .A1(_2707_),
    .S(_2747_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _5173_ (.A0(\u_reg.reg_4[5] ),
    .A1(_2709_),
    .S(_2747_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _5174_ (.A0(\u_reg.reg_4[6] ),
    .A1(_2712_),
    .S(_2747_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _5175_ (.A0(\u_reg.reg_4[7] ),
    .A1(_2714_),
    .S(_2747_),
    .X(_0172_));
 sky130_fd_sc_hd__and3_1 _5176_ (.A(_2653_),
    .B(_2656_),
    .C(_2661_),
    .X(_2748_));
 sky130_fd_sc_hd__and3_1 _5177_ (.A(net1223),
    .B(net1275),
    .C(m2_wbd_sel_i[3]),
    .X(_2749_));
 sky130_fd_sc_hd__a221o_1 _5178_ (.A1(m3_wbd_sel_i[3]),
    .A2(_2013_),
    .B1(_2648_),
    .B2(m1_wbd_sel_i[3]),
    .C1(_2749_),
    .X(_2750_));
 sky130_fd_sc_hd__mux2_1 _5179_ (.A0(m0_wbd_sel_i[3]),
    .A1(_2750_),
    .S(net1148),
    .X(_2751_));
 sky130_fd_sc_hd__and3b_1 _5180_ (.A_N(net619),
    .B(net596),
    .C(net592),
    .X(_2752_));
 sky130_fd_sc_hd__or2_1 _5181_ (.A(m0_wbd_dat_i[24]),
    .B(net1148),
    .X(_2753_));
 sky130_fd_sc_hd__a21o_1 _5182_ (.A1(net1210),
    .A2(m1_wbd_dat_i[24]),
    .B1(net1219),
    .X(_2754_));
 sky130_fd_sc_hd__o211a_2 _5183_ (.A1(net1210),
    .A2(m2_wbd_dat_i[24]),
    .B1(_2753_),
    .C1(_2754_),
    .X(_2755_));
 sky130_fd_sc_hd__mux2_1 _5184_ (.A0(\u_reg.reg_3[24] ),
    .A1(net695),
    .S(net553),
    .X(_0173_));
 sky130_fd_sc_hd__a21o_1 _5185_ (.A1(net1210),
    .A2(m1_wbd_dat_i[25]),
    .B1(net1219),
    .X(_2756_));
 sky130_fd_sc_hd__o221a_2 _5186_ (.A1(net1218),
    .A2(m2_wbd_dat_i[25]),
    .B1(m0_wbd_dat_i[25]),
    .B2(net1148),
    .C1(_2756_),
    .X(_2757_));
 sky130_fd_sc_hd__mux2_1 _5187_ (.A0(\u_reg.reg_3[25] ),
    .A1(net693),
    .S(net553),
    .X(_0174_));
 sky130_fd_sc_hd__a21o_1 _5188_ (.A1(net1215),
    .A2(net1546),
    .B1(net1220),
    .X(_2758_));
 sky130_fd_sc_hd__o221a_1 _5189_ (.A1(net1215),
    .A2(net1523),
    .B1(net1577),
    .B2(net1150),
    .C1(_2758_),
    .X(_2759_));
 sky130_fd_sc_hd__mux2_1 _5190_ (.A0(\u_reg.reg_3[26] ),
    .A1(net692),
    .S(net553),
    .X(_0175_));
 sky130_fd_sc_hd__a21o_1 _5191_ (.A1(net1215),
    .A2(net1545),
    .B1(net1220),
    .X(_2760_));
 sky130_fd_sc_hd__o221a_2 _5192_ (.A1(net1215),
    .A2(net1522),
    .B1(net1576),
    .B2(net1150),
    .C1(_2760_),
    .X(_2761_));
 sky130_fd_sc_hd__mux2_1 _5193_ (.A0(\u_reg.reg_3[27] ),
    .A1(net691),
    .S(net553),
    .X(_0176_));
 sky130_fd_sc_hd__or2_1 _5194_ (.A(m0_wbd_dat_i[28]),
    .B(net1148),
    .X(_2762_));
 sky130_fd_sc_hd__a21o_1 _5195_ (.A1(net1210),
    .A2(m1_wbd_dat_i[28]),
    .B1(net1219),
    .X(_2763_));
 sky130_fd_sc_hd__o211a_2 _5196_ (.A1(net1210),
    .A2(net1895),
    .B1(_2762_),
    .C1(_2763_),
    .X(_2764_));
 sky130_fd_sc_hd__mux2_1 _5197_ (.A0(\u_reg.reg_3[28] ),
    .A1(net690),
    .S(net553),
    .X(_0177_));
 sky130_fd_sc_hd__or2_1 _5198_ (.A(net1575),
    .B(net1149),
    .X(_2765_));
 sky130_fd_sc_hd__a21o_1 _5199_ (.A1(net1221),
    .A2(net1521),
    .B1(net1214),
    .X(_2766_));
 sky130_fd_sc_hd__o211a_1 _5200_ (.A1(net1221),
    .A2(net1544),
    .B1(_2765_),
    .C1(_2766_),
    .X(_2767_));
 sky130_fd_sc_hd__mux2_1 _5201_ (.A0(\u_reg.reg_3[29] ),
    .A1(net689),
    .S(net553),
    .X(_0178_));
 sky130_fd_sc_hd__a21o_1 _5202_ (.A1(net1212),
    .A2(net1542),
    .B1(net1221),
    .X(_2768_));
 sky130_fd_sc_hd__o221a_4 _5203_ (.A1(net1211),
    .A2(net1520),
    .B1(net1573),
    .B2(net1151),
    .C1(_2768_),
    .X(_2769_));
 sky130_fd_sc_hd__mux2_1 _5204_ (.A0(\u_reg.reg_3[30] ),
    .A1(net688),
    .S(net553),
    .X(_0179_));
 sky130_fd_sc_hd__or2_1 _5205_ (.A(net1572),
    .B(net1149),
    .X(_2770_));
 sky130_fd_sc_hd__a21o_1 _5206_ (.A1(net1213),
    .A2(net1541),
    .B1(net1221),
    .X(_2771_));
 sky130_fd_sc_hd__o211a_1 _5207_ (.A1(net1214),
    .A2(net1519),
    .B1(_2770_),
    .C1(_2771_),
    .X(_2772_));
 sky130_fd_sc_hd__mux2_1 _5208_ (.A0(\u_reg.reg_3[31] ),
    .A1(net687),
    .S(_2752_),
    .X(_0180_));
 sky130_fd_sc_hd__and3b_2 _5209_ (.A_N(net619),
    .B(net609),
    .C(net594),
    .X(_2773_));
 sky130_fd_sc_hd__mux2_1 _5210_ (.A0(\u_reg.reg_3[8] ),
    .A1(_2721_),
    .S(_2773_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _5211_ (.A0(\u_reg.reg_3[9] ),
    .A1(net703),
    .S(net552),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _5212_ (.A0(\u_reg.reg_3[10] ),
    .A1(_2725_),
    .S(_2773_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _5213_ (.A0(\u_reg.reg_3[11] ),
    .A1(net702),
    .S(net552),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _5214_ (.A0(\u_reg.reg_3[12] ),
    .A1(net701),
    .S(net552),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _5215_ (.A0(\u_reg.reg_3[13] ),
    .A1(net700),
    .S(net552),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _5216_ (.A0(\u_reg.reg_3[14] ),
    .A1(net699),
    .S(net552),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _5217_ (.A0(\u_reg.reg_3[15] ),
    .A1(net697),
    .S(net552),
    .X(_0188_));
 sky130_fd_sc_hd__and3b_4 _5218_ (.A_N(net618),
    .B(_2694_),
    .C(net593),
    .X(_2774_));
 sky130_fd_sc_hd__mux2_1 _5219_ (.A0(\u_reg.reg_3[0] ),
    .A1(_2697_),
    .S(_2774_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _5220_ (.A0(\u_reg.reg_3[1] ),
    .A1(_2700_),
    .S(_2774_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _5221_ (.A0(\u_reg.reg_3[2] ),
    .A1(_2703_),
    .S(_2774_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _5222_ (.A0(\u_reg.reg_3[3] ),
    .A1(_2705_),
    .S(_2774_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _5223_ (.A0(\u_reg.reg_3[4] ),
    .A1(_2707_),
    .S(_2774_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _5224_ (.A0(\u_reg.reg_3[5] ),
    .A1(_2709_),
    .S(_2774_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _5225_ (.A0(\u_reg.reg_3[6] ),
    .A1(_2712_),
    .S(_2774_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _5226_ (.A0(\u_reg.reg_3[7] ),
    .A1(_2714_),
    .S(_2774_),
    .X(_0196_));
 sky130_fd_sc_hd__and3_1 _5227_ (.A(_2653_),
    .B(_2656_),
    .C(_2662_),
    .X(_2775_));
 sky130_fd_sc_hd__and3b_4 _5228_ (.A_N(net619),
    .B(net609),
    .C(net586),
    .X(_2776_));
 sky130_fd_sc_hd__mux2_1 _5229_ (.A0(\u_reg.reg_2[8] ),
    .A1(_2721_),
    .S(_2776_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _5230_ (.A0(\u_reg.reg_2[9] ),
    .A1(_2723_),
    .S(_2776_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _5231_ (.A0(\u_reg.reg_2[10] ),
    .A1(_2725_),
    .S(_2776_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _5232_ (.A0(\u_reg.reg_2[11] ),
    .A1(net702),
    .S(_2776_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _5233_ (.A0(\u_reg.reg_2[12] ),
    .A1(net701),
    .S(_2776_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _5234_ (.A0(\u_reg.reg_2[13] ),
    .A1(net700),
    .S(_2776_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _5235_ (.A0(\u_reg.reg_2[14] ),
    .A1(net699),
    .S(_2776_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _5236_ (.A0(\u_reg.reg_2[15] ),
    .A1(net698),
    .S(_2776_),
    .X(_0204_));
 sky130_fd_sc_hd__and3b_2 _5237_ (.A_N(net618),
    .B(net617),
    .C(net586),
    .X(_2777_));
 sky130_fd_sc_hd__mux2_1 _5238_ (.A0(\u_reg.reg_2[16] ),
    .A1(net708),
    .S(net551),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _5239_ (.A0(\u_reg.reg_2[17] ),
    .A1(net707),
    .S(net551),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _5240_ (.A0(\u_reg.reg_2[18] ),
    .A1(_2678_),
    .S(_2777_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _5241_ (.A0(\u_reg.reg_2[19] ),
    .A1(_2681_),
    .S(_2777_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _5242_ (.A0(\u_reg.reg_2[20] ),
    .A1(net706),
    .S(net551),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _5243_ (.A0(\u_reg.reg_2[21] ),
    .A1(net705),
    .S(net551),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _5244_ (.A0(\u_reg.reg_2[22] ),
    .A1(_2688_),
    .S(_2777_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _5245_ (.A0(\u_reg.reg_2[23] ),
    .A1(net704),
    .S(net551),
    .X(_0212_));
 sky130_fd_sc_hd__and3b_1 _5246_ (.A_N(net619),
    .B(net592),
    .C(net588),
    .X(_2778_));
 sky130_fd_sc_hd__mux2_1 _5247_ (.A0(\u_reg.reg_2[24] ),
    .A1(net695),
    .S(net550),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _5248_ (.A0(\u_reg.reg_2[25] ),
    .A1(net693),
    .S(net550),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _5249_ (.A0(\u_reg.reg_2[26] ),
    .A1(net692),
    .S(net550),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _5250_ (.A0(\u_reg.reg_2[27] ),
    .A1(net691),
    .S(net550),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _5251_ (.A0(\u_reg.reg_2[28] ),
    .A1(net690),
    .S(_2778_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _5252_ (.A0(\u_reg.reg_2[29] ),
    .A1(net689),
    .S(net550),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _5253_ (.A0(\u_reg.reg_2[30] ),
    .A1(net688),
    .S(net550),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _5254_ (.A0(\u_reg.reg_2[31] ),
    .A1(net687),
    .S(_2778_),
    .X(_0220_));
 sky130_fd_sc_hd__and2b_4 _5255_ (.A_N(_2653_),
    .B(_2656_),
    .X(_2779_));
 sky130_fd_sc_hd__and2_1 _5256_ (.A(_2661_),
    .B(_2779_),
    .X(_2780_));
 sky130_fd_sc_hd__and3b_2 _5257_ (.A_N(net619),
    .B(net609),
    .C(net546),
    .X(_2781_));
 sky130_fd_sc_hd__mux2_1 _5258_ (.A0(\u_dcg_riscv.cfg_mode[0] ),
    .A1(_2721_),
    .S(_2781_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _5259_ (.A0(\u_dcg_riscv.cfg_mode[1] ),
    .A1(net703),
    .S(net512),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _5260_ (.A0(\u_reg.cfg_dcg_ctrl[10] ),
    .A1(_2725_),
    .S(_2781_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _5261_ (.A0(\u_reg.cfg_dcg_ctrl[11] ),
    .A1(net702),
    .S(net512),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _5262_ (.A0(\u_reg.cfg_dcg_ctrl[12] ),
    .A1(net701),
    .S(net512),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _5263_ (.A0(\u_reg.cfg_dcg_ctrl[13] ),
    .A1(net700),
    .S(net512),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _5264_ (.A0(\u_reg.cfg_dcg_ctrl[14] ),
    .A1(net699),
    .S(net512),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _5265_ (.A0(\u_reg.cfg_dcg_ctrl[15] ),
    .A1(net697),
    .S(net512),
    .X(_0228_));
 sky130_fd_sc_hd__and3b_2 _5266_ (.A_N(net618),
    .B(net617),
    .C(net545),
    .X(_2782_));
 sky130_fd_sc_hd__mux2_1 _5267_ (.A0(\u_reg.cfg_dcg_ctrl[16] ),
    .A1(net708),
    .S(net511),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _5268_ (.A0(\u_reg.cfg_dcg_ctrl[17] ),
    .A1(net707),
    .S(net511),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _5269_ (.A0(\u_reg.cfg_dcg_ctrl[18] ),
    .A1(_2678_),
    .S(_2782_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _5270_ (.A0(\u_reg.cfg_dcg_ctrl[19] ),
    .A1(_2681_),
    .S(_2782_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _5271_ (.A0(\u_reg.cfg_dcg_ctrl[20] ),
    .A1(net706),
    .S(net511),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _5272_ (.A0(\u_reg.cfg_dcg_ctrl[21] ),
    .A1(net705),
    .S(net511),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _5273_ (.A0(\u_reg.cfg_dcg_ctrl[22] ),
    .A1(_2688_),
    .S(_2782_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _5274_ (.A0(\u_reg.cfg_dcg_ctrl[23] ),
    .A1(_2690_),
    .S(_2782_),
    .X(_0236_));
 sky130_fd_sc_hd__and3b_2 _5275_ (.A_N(net620),
    .B(net592),
    .C(net548),
    .X(_2783_));
 sky130_fd_sc_hd__mux2_1 _5276_ (.A0(\u_reg.cfg_dcg_ctrl[24] ),
    .A1(net695),
    .S(net510),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _5277_ (.A0(\u_reg.cfg_dcg_ctrl[25] ),
    .A1(net693),
    .S(net510),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _5278_ (.A0(\u_reg.cfg_dcg_ctrl[26] ),
    .A1(net692),
    .S(net510),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _5279_ (.A0(\u_reg.cfg_dcg_ctrl[27] ),
    .A1(net691),
    .S(net510),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _5280_ (.A0(\u_reg.cfg_dcg_ctrl[28] ),
    .A1(net690),
    .S(_2783_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _5281_ (.A0(\u_reg.cfg_dcg_ctrl[29] ),
    .A1(net689),
    .S(net510),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _5282_ (.A0(\u_reg.cfg_dcg_ctrl[30] ),
    .A1(net688),
    .S(net510),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _5283_ (.A0(\u_reg.cfg_dcg_ctrl[31] ),
    .A1(net687),
    .S(_2783_),
    .X(_0244_));
 sky130_fd_sc_hd__or3b_2 _5284_ (.A(_1711_),
    .B(net476),
    .C_N(net438),
    .X(_2784_));
 sky130_fd_sc_hd__or3_1 _5285_ (.A(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[0] ),
    .B(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .C(_2784_),
    .X(_2785_));
 sky130_fd_sc_hd__mux2_1 _5286_ (.A0(net1802),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][0] ),
    .S(net507),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _5287_ (.A0(net1805),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][1] ),
    .S(net507),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _5288_ (.A0(net1797),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][2] ),
    .S(net508),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _5289_ (.A0(net1795),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][3] ),
    .S(net507),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _5290_ (.A0(net1779),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][4] ),
    .S(net508),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _5291_ (.A0(net1796),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][5] ),
    .S(net508),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _5292_ (.A0(net1790),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][6] ),
    .S(net508),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _5293_ (.A0(net1493),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][7] ),
    .S(net506),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _5294_ (.A0(net1831),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][8] ),
    .S(net507),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _5295_ (.A0(net1830),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][9] ),
    .S(net507),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _5296_ (.A0(net1781),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][10] ),
    .S(net508),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _5297_ (.A0(net1813),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][11] ),
    .S(net509),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _5298_ (.A0(net1791),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][12] ),
    .S(net508),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _5299_ (.A0(net1814),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][13] ),
    .S(net509),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _5300_ (.A0(net1811),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][14] ),
    .S(net509),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _5301_ (.A0(net1801),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][15] ),
    .S(net507),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _5302_ (.A0(net1808),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][16] ),
    .S(net506),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _5303_ (.A0(net1806),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][17] ),
    .S(net508),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _5304_ (.A0(net1792),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][18] ),
    .S(net508),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _5305_ (.A0(net1809),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][19] ),
    .S(net507),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _5306_ (.A0(net1829),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][20] ),
    .S(net507),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _5307_ (.A0(net1812),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][21] ),
    .S(net506),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _5308_ (.A0(net1807),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][22] ),
    .S(net506),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _5309_ (.A0(net1828),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][23] ),
    .S(net507),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _5310_ (.A0(net1927),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][24] ),
    .S(net506),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _5311_ (.A0(net1941),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][25] ),
    .S(net506),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _5312_ (.A0(net1937),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][26] ),
    .S(net506),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _5313_ (.A0(net1810),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][27] ),
    .S(net507),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _5314_ (.A0(net1930),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][28] ),
    .S(net506),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _5315_ (.A0(net1494),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][29] ),
    .S(net506),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _5316_ (.A0(net1939),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][30] ),
    .S(net506),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _5317_ (.A0(net1943),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[0][31] ),
    .S(net509),
    .X(_0276_));
 sky130_fd_sc_hd__nor2_1 _5318_ (.A(_1674_),
    .B(_2784_),
    .Y(_2786_));
 sky130_fd_sc_hd__or3_4 _5319_ (.A(_1674_),
    .B(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .C(_2784_),
    .X(_2787_));
 sky130_fd_sc_hd__mux2_1 _5320_ (.A0(net1802),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][0] ),
    .S(net504),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _5321_ (.A0(net1805),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][1] ),
    .S(net504),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _5322_ (.A0(net1797),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][2] ),
    .S(net505),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _5323_ (.A0(net1795),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][3] ),
    .S(net504),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _5324_ (.A0(net1779),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][4] ),
    .S(net505),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _5325_ (.A0(net1796),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][5] ),
    .S(net505),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _5326_ (.A0(net1790),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][6] ),
    .S(net504),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _5327_ (.A0(net1493),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][7] ),
    .S(net503),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _5328_ (.A0(net1831),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][8] ),
    .S(net504),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _5329_ (.A0(net1830),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][9] ),
    .S(net504),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _5330_ (.A0(net1781),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][10] ),
    .S(net505),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _5331_ (.A0(net1813),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][11] ),
    .S(net502),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _5332_ (.A0(net1791),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][12] ),
    .S(net504),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _5333_ (.A0(net1814),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][13] ),
    .S(net503),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _5334_ (.A0(net1811),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][14] ),
    .S(net502),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _5335_ (.A0(net1801),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][15] ),
    .S(net502),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _5336_ (.A0(net1808),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][16] ),
    .S(net502),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _5337_ (.A0(net1806),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][17] ),
    .S(net505),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _5338_ (.A0(net1792),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][18] ),
    .S(net504),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _5339_ (.A0(net1809),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][19] ),
    .S(net502),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _5340_ (.A0(net1829),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][20] ),
    .S(net504),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _5341_ (.A0(net1812),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][21] ),
    .S(net502),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _5342_ (.A0(net1807),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][22] ),
    .S(net503),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _5343_ (.A0(net1828),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][23] ),
    .S(net504),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _5344_ (.A0(net1927),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][24] ),
    .S(net502),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _5345_ (.A0(net1941),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][25] ),
    .S(net503),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _5346_ (.A0(net1937),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][26] ),
    .S(net502),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _5347_ (.A0(net1810),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][27] ),
    .S(net502),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _5348_ (.A0(net1930),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][28] ),
    .S(net502),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _5349_ (.A0(net1494),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][29] ),
    .S(net503),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _5350_ (.A0(net1939),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][30] ),
    .S(net503),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _5351_ (.A0(net1943),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[1][31] ),
    .S(net503),
    .X(_0308_));
 sky130_fd_sc_hd__or3b_4 _5352_ (.A(_2784_),
    .B(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[0] ),
    .C_N(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .X(_2788_));
 sky130_fd_sc_hd__mux2_1 _5353_ (.A0(net1802),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][0] ),
    .S(net500),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _5354_ (.A0(net1805),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][1] ),
    .S(net501),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _5355_ (.A0(net1797),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][2] ),
    .S(net501),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _5356_ (.A0(net1795),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][3] ),
    .S(net501),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _5357_ (.A0(net1779),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][4] ),
    .S(net501),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _5358_ (.A0(net1796),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][5] ),
    .S(net501),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _5359_ (.A0(net1790),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][6] ),
    .S(net500),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _5360_ (.A0(net1493),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][7] ),
    .S(net498),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _5361_ (.A0(net1831),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][8] ),
    .S(net500),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _5362_ (.A0(net1830),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][9] ),
    .S(net500),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _5363_ (.A0(net1781),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][10] ),
    .S(net500),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _5364_ (.A0(net1813),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][11] ),
    .S(net498),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _5365_ (.A0(net1791),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][12] ),
    .S(net501),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _5366_ (.A0(net1814),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][13] ),
    .S(net498),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _5367_ (.A0(net1811),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][14] ),
    .S(net499),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _5368_ (.A0(net1801),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][15] ),
    .S(net500),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _5369_ (.A0(net1808),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][16] ),
    .S(net499),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _5370_ (.A0(net1806),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][17] ),
    .S(net501),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _5371_ (.A0(net1792),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][18] ),
    .S(net500),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _5372_ (.A0(net1809),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][19] ),
    .S(net500),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _5373_ (.A0(net1829),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][20] ),
    .S(net500),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _5374_ (.A0(net1812),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][21] ),
    .S(net498),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _5375_ (.A0(net1807),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][22] ),
    .S(net499),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _5376_ (.A0(net1828),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][23] ),
    .S(net500),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _5377_ (.A0(net1927),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][24] ),
    .S(net498),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _5378_ (.A0(net1941),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][25] ),
    .S(net498),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _5379_ (.A0(net1937),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][26] ),
    .S(net498),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _5380_ (.A0(net1810),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][27] ),
    .S(net499),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _5381_ (.A0(net1930),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][28] ),
    .S(net499),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _5382_ (.A0(net1494),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][29] ),
    .S(net498),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _5383_ (.A0(net1939),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][30] ),
    .S(net498),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _5384_ (.A0(net1943),
    .A1(\u_s2.u_sync_wbb.u_resp_if.mem[2][31] ),
    .S(net498),
    .X(_0340_));
 sky130_fd_sc_hd__and2_4 _5385_ (.A(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .B(_2786_),
    .X(_2789_));
 sky130_fd_sc_hd__mux2_1 _5386_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][0] ),
    .A1(net1802),
    .S(net483),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _5387_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][1] ),
    .A1(net1805),
    .S(net484),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _5388_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][2] ),
    .A1(net1797),
    .S(net484),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _5389_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][3] ),
    .A1(net1795),
    .S(net483),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _5390_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][4] ),
    .A1(net1779),
    .S(net483),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _5391_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][5] ),
    .A1(net1796),
    .S(net484),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _5392_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][6] ),
    .A1(net1790),
    .S(net483),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _5393_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][7] ),
    .A1(net1493),
    .S(net481),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _5394_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][8] ),
    .A1(net1831),
    .S(net483),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _5395_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][9] ),
    .A1(net1830),
    .S(net483),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _5396_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][10] ),
    .A1(net1781),
    .S(net484),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _5397_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][11] ),
    .A1(net1813),
    .S(net481),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _5398_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][12] ),
    .A1(net1791),
    .S(net484),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _5399_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][13] ),
    .A1(net1814),
    .S(net481),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _5400_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][14] ),
    .A1(net1811),
    .S(net482),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _5401_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][15] ),
    .A1(net1801),
    .S(net481),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _5402_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][16] ),
    .A1(net1808),
    .S(net482),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _5403_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][17] ),
    .A1(net1806),
    .S(net484),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _5404_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][18] ),
    .A1(net1792),
    .S(net483),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _5405_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][19] ),
    .A1(net1809),
    .S(net482),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _5406_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][20] ),
    .A1(net1829),
    .S(net483),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _5407_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][21] ),
    .A1(net1812),
    .S(net481),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _5408_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][22] ),
    .A1(net1807),
    .S(net482),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _5409_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][23] ),
    .A1(net1828),
    .S(net483),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _5410_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][24] ),
    .A1(net1927),
    .S(net482),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _5411_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][25] ),
    .A1(net1941),
    .S(net481),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _5412_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][26] ),
    .A1(net1937),
    .S(net481),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _5413_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][27] ),
    .A1(net1810),
    .S(net482),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _5414_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][28] ),
    .A1(net1930),
    .S(net482),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _5415_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][29] ),
    .A1(net1494),
    .S(net481),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _5416_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][30] ),
    .A1(net1939),
    .S(net481),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _5417_ (.A0(\u_s2.u_sync_wbb.u_resp_if.mem[3][31] ),
    .A1(net1943),
    .S(net481),
    .X(_0372_));
 sky130_fd_sc_hd__mux4_2 _5418_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][1] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][1] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][1] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][1] ),
    .S0(net1360),
    .S1(net1353),
    .X(_2790_));
 sky130_fd_sc_hd__mux2_1 _5419_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[1] ),
    .A1(_2790_),
    .S(net1510),
    .X(_0373_));
 sky130_fd_sc_hd__mux4_2 _5420_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][2] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][2] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][2] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][2] ),
    .S0(net1359),
    .S1(net1352),
    .X(_2791_));
 sky130_fd_sc_hd__mux2_1 _5421_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[2] ),
    .A1(_2791_),
    .S(net1507),
    .X(_0374_));
 sky130_fd_sc_hd__mux4_1 _5422_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][3] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][3] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][3] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][3] ),
    .S0(net1362),
    .S1(net1355),
    .X(_2792_));
 sky130_fd_sc_hd__mux2_1 _5423_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[3] ),
    .A1(_2792_),
    .S(net1509),
    .X(_0375_));
 sky130_fd_sc_hd__mux4_2 _5424_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][4] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][4] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][4] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][4] ),
    .S0(net1360),
    .S1(net1353),
    .X(_2793_));
 sky130_fd_sc_hd__mux2_1 _5425_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[4] ),
    .A1(_2793_),
    .S(net1507),
    .X(_0376_));
 sky130_fd_sc_hd__mux4_1 _5426_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][5] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][5] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][5] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][5] ),
    .S0(net1364),
    .S1(net1357),
    .X(_2794_));
 sky130_fd_sc_hd__mux2_1 _5427_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[5] ),
    .A1(_2794_),
    .S(net1507),
    .X(_0377_));
 sky130_fd_sc_hd__mux4_1 _5428_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][6] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][6] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][6] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][6] ),
    .S0(net1363),
    .S1(net1356),
    .X(_2795_));
 sky130_fd_sc_hd__mux2_1 _5429_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[6] ),
    .A1(_2795_),
    .S(net1507),
    .X(_0378_));
 sky130_fd_sc_hd__mux4_2 _5430_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][7] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][7] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][7] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][7] ),
    .S0(net1359),
    .S1(net1352),
    .X(_2796_));
 sky130_fd_sc_hd__mux2_1 _5431_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[7] ),
    .A1(_2796_),
    .S(net1507),
    .X(_0379_));
 sky130_fd_sc_hd__mux4_1 _5432_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][8] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][8] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][8] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][8] ),
    .S0(net1360),
    .S1(net1353),
    .X(_2797_));
 sky130_fd_sc_hd__mux2_1 _5433_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[8] ),
    .A1(_2797_),
    .S(net1508),
    .X(_0380_));
 sky130_fd_sc_hd__mux4_2 _5434_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[0][9] ),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[1][9] ),
    .A2(\u_s1.u_sync_wbb.u_cmd_if.mem[2][9] ),
    .A3(\u_s1.u_sync_wbb.u_cmd_if.mem[3][9] ),
    .S0(net1359),
    .S1(net1352),
    .X(_2798_));
 sky130_fd_sc_hd__mux2_1 _5435_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[9] ),
    .A1(_2798_),
    .S(net1507),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _5436_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[14] ),
    .A1(_2374_),
    .S(net1508),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _5437_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[15] ),
    .A1(_2375_),
    .S(net1504),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _5438_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[16] ),
    .A1(_2376_),
    .S(net1507),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _5439_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[17] ),
    .A1(_2377_),
    .S(net1507),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _5440_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[18] ),
    .A1(_2378_),
    .S(net1504),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _5441_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[19] ),
    .A1(_2379_),
    .S(net1506),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _5442_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[20] ),
    .A1(_2380_),
    .S(net1509),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _5443_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[21] ),
    .A1(_2381_),
    .S(net1509),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _5444_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[22] ),
    .A1(_2382_),
    .S(net1508),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _5445_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[23] ),
    .A1(_2383_),
    .S(net1505),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _5446_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[24] ),
    .A1(_2384_),
    .S(net1505),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _5447_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[25] ),
    .A1(_2385_),
    .S(net1509),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _5448_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[26] ),
    .A1(_2386_),
    .S(net1509),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _5449_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[27] ),
    .A1(_2387_),
    .S(net1508),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _5450_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[28] ),
    .A1(_2388_),
    .S(net1509),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _5451_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[29] ),
    .A1(_2389_),
    .S(net1508),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _5452_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[30] ),
    .A1(_2390_),
    .S(net1509),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_1 _5453_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[31] ),
    .A1(_2391_),
    .S(net1506),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _5454_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[32] ),
    .A1(_2392_),
    .S(net1505),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _5455_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[33] ),
    .A1(_2393_),
    .S(net1503),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _5456_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[34] ),
    .A1(_2394_),
    .S(net1505),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _5457_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[35] ),
    .A1(_2395_),
    .S(net1508),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _5458_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[36] ),
    .A1(_2396_),
    .S(net1503),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_1 _5459_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[37] ),
    .A1(_2397_),
    .S(net1503),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _5460_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[38] ),
    .A1(_2398_),
    .S(net1508),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _5461_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[39] ),
    .A1(_2399_),
    .S(net1503),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _5462_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[40] ),
    .A1(_2400_),
    .S(net1503),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _5463_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[41] ),
    .A1(_2401_),
    .S(net1509),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _5464_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[42] ),
    .A1(_2402_),
    .S(net1503),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _5465_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[43] ),
    .A1(_2403_),
    .S(net1506),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _5466_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[44] ),
    .A1(_2404_),
    .S(net1503),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _5467_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[45] ),
    .A1(_2405_),
    .S(net1509),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _5468_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[46] ),
    .A1(_2406_),
    .S(net1508),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _5469_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[47] ),
    .A1(_2407_),
    .S(net1503),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _5470_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[48] ),
    .A1(_2408_),
    .S(net1506),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _5471_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[49] ),
    .A1(_2409_),
    .S(net1503),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _5472_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[50] ),
    .A1(_2006_),
    .S(net1505),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _5473_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[53] ),
    .A1(_2410_),
    .S(net1504),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _5474_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[54] ),
    .A1(_2411_),
    .S(net1505),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _5475_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[55] ),
    .A1(_2412_),
    .S(net1505),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _5476_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[56] ),
    .A1(_2413_),
    .S(net1505),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _5477_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[57] ),
    .A1(_2414_),
    .S(net1503),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _5478_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[58] ),
    .A1(_2415_),
    .S(net1505),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _5479_ (.A0(\u_s1.u_sync_wbb.s_cmd_rd_data_l[59] ),
    .A1(_2416_),
    .S(net1504),
    .X(_0425_));
 sky130_fd_sc_hd__nand2_1 _5480_ (.A(net1952),
    .B(\u_s1.u_sync_wbb.m_cmd_wr_en ),
    .Y(_2799_));
 sky130_fd_sc_hd__and3_4 _5481_ (.A(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .B(net1952),
    .C(\u_s1.u_sync_wbb.m_cmd_wr_en ),
    .X(_2800_));
 sky130_fd_sc_hd__mux2_1 _5482_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][1] ),
    .A1(net797),
    .S(net1000),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _5483_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][2] ),
    .A1(net798),
    .S(net999),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _5484_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][3] ),
    .A1(_1860_),
    .S(net1001),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _5485_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][4] ),
    .A1(_1856_),
    .S(net998),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _5486_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][5] ),
    .A1(_1869_),
    .S(net1002),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _5487_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][6] ),
    .A1(_1868_),
    .S(net1002),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _5488_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][7] ),
    .A1(_1867_),
    .S(net999),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _5489_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][8] ),
    .A1(_1866_),
    .S(net1001),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _5490_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][9] ),
    .A1(_1873_),
    .S(net998),
    .X(_0434_));
 sky130_fd_sc_hd__a221o_1 _5491_ (.A1(net1240),
    .A2(m2_wbd_sel_i[0]),
    .B1(net1186),
    .B2(m3_wbd_sel_i[0]),
    .C1(net1192),
    .X(_2801_));
 sky130_fd_sc_hd__and2_1 _5492_ (.A(m1_wbd_sel_i[0]),
    .B(net1184),
    .X(_2802_));
 sky130_fd_sc_hd__o22a_1 _5493_ (.A1(net1565),
    .A2(_1831_),
    .B1(_2801_),
    .B2(_2802_),
    .X(_2803_));
 sky130_fd_sc_hd__mux2_1 _5494_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][14] ),
    .A1(net686),
    .S(net1003),
    .X(_0435_));
 sky130_fd_sc_hd__and3_1 _5495_ (.A(net1404),
    .B(net1405),
    .C(m3_wbd_sel_i[1]),
    .X(_2804_));
 sky130_fd_sc_hd__a221o_1 _5496_ (.A1(net1239),
    .A2(m2_wbd_sel_i[1]),
    .B1(m1_wbd_sel_i[1]),
    .B2(net1183),
    .C1(net1192),
    .X(_2805_));
 sky130_fd_sc_hd__o22a_1 _5497_ (.A1(m0_wbd_sel_i[1]),
    .A2(net1188),
    .B1(_2804_),
    .B2(_2805_),
    .X(_2806_));
 sky130_fd_sc_hd__mux2_1 _5498_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][15] ),
    .A1(net685),
    .S(net1000),
    .X(_0436_));
 sky130_fd_sc_hd__and2_1 _5499_ (.A(m1_wbd_sel_i[2]),
    .B(_1833_),
    .X(_2807_));
 sky130_fd_sc_hd__a221o_1 _5500_ (.A1(net1239),
    .A2(m2_wbd_sel_i[2]),
    .B1(net1185),
    .B2(m3_wbd_sel_i[2]),
    .C1(_1830_),
    .X(_2808_));
 sky130_fd_sc_hd__o22a_1 _5501_ (.A1(m0_wbd_sel_i[2]),
    .A2(net1187),
    .B1(_2807_),
    .B2(_2808_),
    .X(_2809_));
 sky130_fd_sc_hd__mux2_1 _5502_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][16] ),
    .A1(net684),
    .S(net1001),
    .X(_0437_));
 sky130_fd_sc_hd__and2_1 _5503_ (.A(m1_wbd_sel_i[3]),
    .B(net1183),
    .X(_2810_));
 sky130_fd_sc_hd__a221o_1 _5504_ (.A1(net1239),
    .A2(m2_wbd_sel_i[3]),
    .B1(net1185),
    .B2(m3_wbd_sel_i[3]),
    .C1(net1192),
    .X(_2811_));
 sky130_fd_sc_hd__o22a_2 _5505_ (.A1(m0_wbd_sel_i[3]),
    .A2(net1187),
    .B1(_2810_),
    .B2(_2811_),
    .X(_2812_));
 sky130_fd_sc_hd__mux2_1 _5506_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][17] ),
    .A1(net683),
    .S(net1002),
    .X(_0438_));
 sky130_fd_sc_hd__a21o_1 _5507_ (.A1(net1246),
    .A2(net1562),
    .B1(net1240),
    .X(_2813_));
 sky130_fd_sc_hd__o221a_1 _5508_ (.A1(net1246),
    .A2(m2_wbd_dat_i[0]),
    .B1(net1593),
    .B2(net1188),
    .C1(_2813_),
    .X(_2814_));
 sky130_fd_sc_hd__mux2_1 _5509_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][18] ),
    .A1(net682),
    .S(net1004),
    .X(_0439_));
 sky130_fd_sc_hd__a21o_1 _5510_ (.A1(net1246),
    .A2(net1551),
    .B1(net1240),
    .X(_2815_));
 sky130_fd_sc_hd__o221a_4 _5511_ (.A1(net1246),
    .A2(m2_wbd_dat_i[1]),
    .B1(net1582),
    .B2(net1188),
    .C1(_2815_),
    .X(_2816_));
 sky130_fd_sc_hd__mux2_1 _5512_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][19] ),
    .A1(_2816_),
    .S(net1002),
    .X(_0440_));
 sky130_fd_sc_hd__a21o_1 _5513_ (.A1(net1248),
    .A2(net1543),
    .B1(net1244),
    .X(_2817_));
 sky130_fd_sc_hd__o221a_4 _5514_ (.A1(net1248),
    .A2(m2_wbd_dat_i[2]),
    .B1(net1574),
    .B2(net1191),
    .C1(_2817_),
    .X(_2818_));
 sky130_fd_sc_hd__mux2_1 _5515_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][20] ),
    .A1(_2818_),
    .S(net1001),
    .X(_0441_));
 sky130_fd_sc_hd__a21o_1 _5516_ (.A1(net1245),
    .A2(m1_wbd_dat_i[3]),
    .B1(net1240),
    .X(_2819_));
 sky130_fd_sc_hd__o221a_1 _5517_ (.A1(net1245),
    .A2(net2088),
    .B1(m0_wbd_dat_i[3]),
    .B2(net1187),
    .C1(_2819_),
    .X(_2820_));
 sky130_fd_sc_hd__mux2_1 _5518_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][21] ),
    .A1(net681),
    .S(net1001),
    .X(_0442_));
 sky130_fd_sc_hd__or2_1 _5519_ (.A(net1571),
    .B(net1191),
    .X(_2821_));
 sky130_fd_sc_hd__a21o_1 _5520_ (.A1(net1244),
    .A2(net1518),
    .B1(net1248),
    .X(_2822_));
 sky130_fd_sc_hd__o211a_4 _5521_ (.A1(net1244),
    .A2(net1540),
    .B1(_2821_),
    .C1(_2822_),
    .X(_2823_));
 sky130_fd_sc_hd__mux2_1 _5522_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][22] ),
    .A1(_2823_),
    .S(net1003),
    .X(_0443_));
 sky130_fd_sc_hd__a21o_1 _5523_ (.A1(net1251),
    .A2(net1539),
    .B1(net1243),
    .X(_2824_));
 sky130_fd_sc_hd__o221a_4 _5524_ (.A1(net1251),
    .A2(net1517),
    .B1(net1570),
    .B2(net1190),
    .C1(_2824_),
    .X(_2825_));
 sky130_fd_sc_hd__mux2_1 _5525_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][23] ),
    .A1(_2825_),
    .S(net1003),
    .X(_0444_));
 sky130_fd_sc_hd__a21o_1 _5526_ (.A1(net1249),
    .A2(net1538),
    .B1(net1242),
    .X(_2826_));
 sky130_fd_sc_hd__o221a_1 _5527_ (.A1(net1249),
    .A2(net1516),
    .B1(net1569),
    .B2(net1189),
    .C1(_2826_),
    .X(_2827_));
 sky130_fd_sc_hd__mux2_1 _5528_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][24] ),
    .A1(_2827_),
    .S(net1000),
    .X(_0445_));
 sky130_fd_sc_hd__or2_1 _5529_ (.A(net1568),
    .B(net1189),
    .X(_2828_));
 sky130_fd_sc_hd__a21o_1 _5530_ (.A1(net1242),
    .A2(net1515),
    .B1(net1249),
    .X(_2829_));
 sky130_fd_sc_hd__o211a_2 _5531_ (.A1(net1242),
    .A2(net1537),
    .B1(_2828_),
    .C1(_2829_),
    .X(_2830_));
 sky130_fd_sc_hd__mux2_1 _5532_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][25] ),
    .A1(_2830_),
    .S(net1002),
    .X(_0446_));
 sky130_fd_sc_hd__a21o_1 _5533_ (.A1(net1249),
    .A2(net1536),
    .B1(net1241),
    .X(_2831_));
 sky130_fd_sc_hd__o221a_2 _5534_ (.A1(net1249),
    .A2(net1514),
    .B1(net1567),
    .B2(net1190),
    .C1(_2831_),
    .X(_2832_));
 sky130_fd_sc_hd__mux2_1 _5535_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][26] ),
    .A1(_2832_),
    .S(net1002),
    .X(_0447_));
 sky130_fd_sc_hd__or2_1 _5536_ (.A(net1566),
    .B(net1189),
    .X(_2833_));
 sky130_fd_sc_hd__a21o_1 _5537_ (.A1(net1241),
    .A2(net1513),
    .B1(net1249),
    .X(_2834_));
 sky130_fd_sc_hd__o211a_2 _5538_ (.A1(net1241),
    .A2(net1535),
    .B1(_2833_),
    .C1(_2834_),
    .X(_2835_));
 sky130_fd_sc_hd__mux2_1 _5539_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][27] ),
    .A1(_2835_),
    .S(net1003),
    .X(_0448_));
 sky130_fd_sc_hd__or2_1 _5540_ (.A(net1592),
    .B(net1190),
    .X(_2836_));
 sky130_fd_sc_hd__a21o_1 _5541_ (.A1(net1243),
    .A2(net1534),
    .B1(net1251),
    .X(_2837_));
 sky130_fd_sc_hd__o211a_4 _5542_ (.A1(net1243),
    .A2(net1561),
    .B1(_2836_),
    .C1(_2837_),
    .X(_2838_));
 sky130_fd_sc_hd__mux2_1 _5543_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][28] ),
    .A1(_2838_),
    .S(net1004),
    .X(_0449_));
 sky130_fd_sc_hd__or2_1 _5544_ (.A(net1591),
    .B(net1190),
    .X(_2839_));
 sky130_fd_sc_hd__a21o_1 _5545_ (.A1(net1243),
    .A2(net1533),
    .B1(net1251),
    .X(_2840_));
 sky130_fd_sc_hd__o211a_4 _5546_ (.A1(net1243),
    .A2(net1560),
    .B1(_2839_),
    .C1(_2840_),
    .X(_2841_));
 sky130_fd_sc_hd__mux2_1 _5547_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][29] ),
    .A1(_2841_),
    .S(net1004),
    .X(_0450_));
 sky130_fd_sc_hd__or2_1 _5548_ (.A(net1590),
    .B(net1189),
    .X(_2842_));
 sky130_fd_sc_hd__a21o_1 _5549_ (.A1(net1241),
    .A2(net1532),
    .B1(net1250),
    .X(_2843_));
 sky130_fd_sc_hd__o211a_2 _5550_ (.A1(net1242),
    .A2(net1559),
    .B1(_2842_),
    .C1(_2843_),
    .X(_2844_));
 sky130_fd_sc_hd__mux2_1 _5551_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][30] ),
    .A1(_2844_),
    .S(net1004),
    .X(_0451_));
 sky130_fd_sc_hd__a21o_1 _5552_ (.A1(net1247),
    .A2(net1558),
    .B1(net1244),
    .X(_2845_));
 sky130_fd_sc_hd__o221a_2 _5553_ (.A1(net1247),
    .A2(net2066),
    .B1(net1589),
    .B2(net1191),
    .C1(_2845_),
    .X(_2846_));
 sky130_fd_sc_hd__mux2_1 _5554_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][31] ),
    .A1(_2846_),
    .S(net1000),
    .X(_0452_));
 sky130_fd_sc_hd__or2_1 _5555_ (.A(net1588),
    .B(net1190),
    .X(_2847_));
 sky130_fd_sc_hd__a21o_1 _5556_ (.A1(net1243),
    .A2(net1531),
    .B1(net1251),
    .X(_2848_));
 sky130_fd_sc_hd__o211a_2 _5557_ (.A1(net1243),
    .A2(net1557),
    .B1(_2847_),
    .C1(_2848_),
    .X(_2849_));
 sky130_fd_sc_hd__mux2_1 _5558_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][32] ),
    .A1(_2849_),
    .S(net1001),
    .X(_0453_));
 sky130_fd_sc_hd__a21o_1 _5559_ (.A1(net1248),
    .A2(net1556),
    .B1(net1244),
    .X(_2850_));
 sky130_fd_sc_hd__o221a_1 _5560_ (.A1(net1248),
    .A2(net1530),
    .B1(net1587),
    .B2(net1191),
    .C1(_2850_),
    .X(_2851_));
 sky130_fd_sc_hd__mux2_1 _5561_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][33] ),
    .A1(_2851_),
    .S(net999),
    .X(_0454_));
 sky130_fd_sc_hd__or2_1 _5562_ (.A(net1586),
    .B(net1189),
    .X(_2852_));
 sky130_fd_sc_hd__a21o_1 _5563_ (.A1(net1241),
    .A2(net1529),
    .B1(net1249),
    .X(_2853_));
 sky130_fd_sc_hd__o211a_2 _5564_ (.A1(net1241),
    .A2(net1555),
    .B1(_2852_),
    .C1(_2853_),
    .X(_2854_));
 sky130_fd_sc_hd__mux2_1 _5565_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][34] ),
    .A1(_2854_),
    .S(net1002),
    .X(_0455_));
 sky130_fd_sc_hd__a21o_1 _5566_ (.A1(net1250),
    .A2(net1554),
    .B1(net1242),
    .X(_2855_));
 sky130_fd_sc_hd__o221a_2 _5567_ (.A1(net1250),
    .A2(net1528),
    .B1(net1585),
    .B2(net1189),
    .C1(_2855_),
    .X(_2856_));
 sky130_fd_sc_hd__mux2_1 _5568_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][35] ),
    .A1(_2856_),
    .S(net1003),
    .X(_0456_));
 sky130_fd_sc_hd__a21o_1 _5569_ (.A1(net1246),
    .A2(net1553),
    .B1(net1240),
    .X(_2857_));
 sky130_fd_sc_hd__o221a_2 _5570_ (.A1(net1246),
    .A2(net2056),
    .B1(net1584),
    .B2(net1188),
    .C1(_2857_),
    .X(_2858_));
 sky130_fd_sc_hd__mux2_1 _5571_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][36] ),
    .A1(_2858_),
    .S(net998),
    .X(_0457_));
 sky130_fd_sc_hd__or2_1 _5572_ (.A(net1583),
    .B(net1189),
    .X(_2859_));
 sky130_fd_sc_hd__a21o_1 _5573_ (.A1(net1241),
    .A2(net1527),
    .B1(net1250),
    .X(_2860_));
 sky130_fd_sc_hd__o211a_2 _5574_ (.A1(net1241),
    .A2(net1552),
    .B1(_2859_),
    .C1(_2860_),
    .X(_2861_));
 sky130_fd_sc_hd__mux2_1 _5575_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][37] ),
    .A1(_2861_),
    .S(net1002),
    .X(_0458_));
 sky130_fd_sc_hd__a21o_1 _5576_ (.A1(net1251),
    .A2(net1550),
    .B1(net1243),
    .X(_2862_));
 sky130_fd_sc_hd__o221a_2 _5577_ (.A1(net1249),
    .A2(net1526),
    .B1(net1581),
    .B2(net1189),
    .C1(_2862_),
    .X(_2863_));
 sky130_fd_sc_hd__mux2_1 _5578_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][38] ),
    .A1(_2863_),
    .S(net1001),
    .X(_0459_));
 sky130_fd_sc_hd__a21o_1 _5579_ (.A1(net1247),
    .A2(net1549),
    .B1(net1244),
    .X(_2864_));
 sky130_fd_sc_hd__o221a_1 _5580_ (.A1(net1247),
    .A2(net1525),
    .B1(net1580),
    .B2(net1191),
    .C1(_2864_),
    .X(_2865_));
 sky130_fd_sc_hd__mux2_1 _5581_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][39] ),
    .A1(_2865_),
    .S(net999),
    .X(_0460_));
 sky130_fd_sc_hd__a21o_1 _5582_ (.A1(net1246),
    .A2(net1548),
    .B1(net1244),
    .X(_2866_));
 sky130_fd_sc_hd__o221a_2 _5583_ (.A1(net1246),
    .A2(net2051),
    .B1(net1579),
    .B2(net1191),
    .C1(_2866_),
    .X(_2867_));
 sky130_fd_sc_hd__mux2_1 _5584_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][40] ),
    .A1(_2867_),
    .S(net998),
    .X(_0461_));
 sky130_fd_sc_hd__a21o_1 _5585_ (.A1(net1247),
    .A2(net1547),
    .B1(net1244),
    .X(_2868_));
 sky130_fd_sc_hd__o221a_2 _5586_ (.A1(net1247),
    .A2(net1524),
    .B1(net1578),
    .B2(net1191),
    .C1(_2868_),
    .X(_2869_));
 sky130_fd_sc_hd__mux2_1 _5587_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][41] ),
    .A1(_2869_),
    .S(net1000),
    .X(_0462_));
 sky130_fd_sc_hd__a21o_1 _5588_ (.A1(net1245),
    .A2(m1_wbd_dat_i[24]),
    .B1(net1239),
    .X(_2870_));
 sky130_fd_sc_hd__o221a_1 _5589_ (.A1(net1245),
    .A2(m2_wbd_dat_i[24]),
    .B1(m0_wbd_dat_i[24]),
    .B2(net1187),
    .C1(_2870_),
    .X(_2871_));
 sky130_fd_sc_hd__mux2_1 _5590_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][42] ),
    .A1(net680),
    .S(net1002),
    .X(_0463_));
 sky130_fd_sc_hd__a21o_1 _5591_ (.A1(net1245),
    .A2(m1_wbd_dat_i[25]),
    .B1(net1239),
    .X(_2872_));
 sky130_fd_sc_hd__o221a_4 _5592_ (.A1(net1245),
    .A2(net2079),
    .B1(m0_wbd_dat_i[25]),
    .B2(net1187),
    .C1(_2872_),
    .X(_2873_));
 sky130_fd_sc_hd__mux2_1 _5593_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][43] ),
    .A1(net2080),
    .S(net1000),
    .X(_0464_));
 sky130_fd_sc_hd__a21o_1 _5594_ (.A1(net1249),
    .A2(net1546),
    .B1(net1241),
    .X(_2874_));
 sky130_fd_sc_hd__o221a_2 _5595_ (.A1(net1249),
    .A2(net1523),
    .B1(net1577),
    .B2(net1189),
    .C1(_2874_),
    .X(_2875_));
 sky130_fd_sc_hd__mux2_1 _5596_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][44] ),
    .A1(_2875_),
    .S(net998),
    .X(_0465_));
 sky130_fd_sc_hd__a21o_1 _5597_ (.A1(net1250),
    .A2(net1545),
    .B1(net1241),
    .X(_2876_));
 sky130_fd_sc_hd__o221a_2 _5598_ (.A1(net1250),
    .A2(net1522),
    .B1(net1576),
    .B2(net1189),
    .C1(_2876_),
    .X(_2877_));
 sky130_fd_sc_hd__mux2_1 _5599_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][45] ),
    .A1(_2877_),
    .S(net1003),
    .X(_0466_));
 sky130_fd_sc_hd__a21o_1 _5600_ (.A1(net1246),
    .A2(m1_wbd_dat_i[28]),
    .B1(net1239),
    .X(_2878_));
 sky130_fd_sc_hd__o221a_4 _5601_ (.A1(net1245),
    .A2(m2_wbd_dat_i[28]),
    .B1(m0_wbd_dat_i[28]),
    .B2(net1187),
    .C1(_2878_),
    .X(_2879_));
 sky130_fd_sc_hd__mux2_1 _5602_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][46] ),
    .A1(net679),
    .S(net1004),
    .X(_0467_));
 sky130_fd_sc_hd__a21o_1 _5603_ (.A1(net1247),
    .A2(net1544),
    .B1(net1244),
    .X(_2880_));
 sky130_fd_sc_hd__o221a_2 _5604_ (.A1(net1247),
    .A2(net1521),
    .B1(net1575),
    .B2(net1191),
    .C1(_2880_),
    .X(_2881_));
 sky130_fd_sc_hd__mux2_1 _5605_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][47] ),
    .A1(_2881_),
    .S(net998),
    .X(_0468_));
 sky130_fd_sc_hd__a21o_1 _5606_ (.A1(net1247),
    .A2(net1542),
    .B1(net1244),
    .X(_2882_));
 sky130_fd_sc_hd__o221a_1 _5607_ (.A1(net1247),
    .A2(net1520),
    .B1(net1573),
    .B2(net1191),
    .C1(_2882_),
    .X(_2883_));
 sky130_fd_sc_hd__mux2_1 _5608_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][48] ),
    .A1(_2883_),
    .S(net999),
    .X(_0469_));
 sky130_fd_sc_hd__a21o_1 _5609_ (.A1(net1251),
    .A2(net1541),
    .B1(net1243),
    .X(_2884_));
 sky130_fd_sc_hd__o221a_2 _5610_ (.A1(net1251),
    .A2(net1519),
    .B1(net1572),
    .B2(net1190),
    .C1(_2884_),
    .X(_2885_));
 sky130_fd_sc_hd__mux2_1 _5611_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][49] ),
    .A1(_2885_),
    .S(net998),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _5612_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][50] ),
    .A1(net732),
    .S(net1002),
    .X(_0471_));
 sky130_fd_sc_hd__and3_1 _5613_ (.A(net1404),
    .B(net1406),
    .C(m3_wbd_adr_i[2]),
    .X(_2886_));
 sky130_fd_sc_hd__a221o_1 _5614_ (.A1(net1240),
    .A2(m2_wbd_adr_i[2]),
    .B1(m1_wbd_adr_i[2]),
    .B2(net1183),
    .C1(net1192),
    .X(_2887_));
 sky130_fd_sc_hd__o22a_2 _5615_ (.A1(net1598),
    .A2(net1188),
    .B1(_2886_),
    .B2(_2887_),
    .X(_2888_));
 sky130_fd_sc_hd__mux2_1 _5616_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][53] ),
    .A1(_2888_),
    .S(net998),
    .X(_0472_));
 sky130_fd_sc_hd__and3_1 _5617_ (.A(\u_s1.gnt[1] ),
    .B(net1406),
    .C(m3_wbd_adr_i[3]),
    .X(_2889_));
 sky130_fd_sc_hd__a221o_1 _5618_ (.A1(net1240),
    .A2(m2_wbd_adr_i[3]),
    .B1(m1_wbd_adr_i[3]),
    .B2(net1184),
    .C1(net1192),
    .X(_2890_));
 sky130_fd_sc_hd__o22a_4 _5619_ (.A1(net1597),
    .A2(net1188),
    .B1(_2889_),
    .B2(_2890_),
    .X(_2891_));
 sky130_fd_sc_hd__mux2_1 _5620_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][54] ),
    .A1(_2891_),
    .S(net1000),
    .X(_0473_));
 sky130_fd_sc_hd__and2_1 _5621_ (.A(m1_wbd_adr_i[4]),
    .B(net1183),
    .X(_2892_));
 sky130_fd_sc_hd__a221o_1 _5622_ (.A1(net1239),
    .A2(m2_wbd_adr_i[4]),
    .B1(net1185),
    .B2(m3_wbd_adr_i[4]),
    .C1(net1192),
    .X(_2893_));
 sky130_fd_sc_hd__o22a_4 _5623_ (.A1(net1596),
    .A2(net1188),
    .B1(_2892_),
    .B2(_2893_),
    .X(_2894_));
 sky130_fd_sc_hd__mux2_1 _5624_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][55] ),
    .A1(_2894_),
    .S(net1000),
    .X(_0474_));
 sky130_fd_sc_hd__and2_1 _5625_ (.A(m1_wbd_adr_i[5]),
    .B(net1184),
    .X(_2895_));
 sky130_fd_sc_hd__a221o_1 _5626_ (.A1(_1673_),
    .A2(net2092),
    .B1(_1832_),
    .B2(m3_wbd_adr_i[5]),
    .C1(net1192),
    .X(_2896_));
 sky130_fd_sc_hd__o22a_4 _5627_ (.A1(net1595),
    .A2(net1188),
    .B1(_2895_),
    .B2(_2896_),
    .X(_2897_));
 sky130_fd_sc_hd__mux2_1 _5628_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][56] ),
    .A1(_2897_),
    .S(net1000),
    .X(_0475_));
 sky130_fd_sc_hd__and2_1 _5629_ (.A(m1_wbd_adr_i[6]),
    .B(net1183),
    .X(_2898_));
 sky130_fd_sc_hd__a221o_1 _5630_ (.A1(net1240),
    .A2(m2_wbd_adr_i[6]),
    .B1(net1185),
    .B2(m3_wbd_adr_i[6]),
    .C1(net1192),
    .X(_2899_));
 sky130_fd_sc_hd__o22a_4 _5631_ (.A1(net2035),
    .A2(net1187),
    .B1(_2898_),
    .B2(_2899_),
    .X(_2900_));
 sky130_fd_sc_hd__mux2_1 _5632_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][57] ),
    .A1(_2900_),
    .S(net998),
    .X(_0476_));
 sky130_fd_sc_hd__and2_1 _5633_ (.A(m1_wbd_adr_i[7]),
    .B(net1184),
    .X(_2901_));
 sky130_fd_sc_hd__a221o_1 _5634_ (.A1(net1239),
    .A2(m2_wbd_adr_i[7]),
    .B1(net1185),
    .B2(m3_wbd_adr_i[7]),
    .C1(_1830_),
    .X(_2902_));
 sky130_fd_sc_hd__o22a_4 _5635_ (.A1(net1594),
    .A2(net1188),
    .B1(_2901_),
    .B2(_2902_),
    .X(_2903_));
 sky130_fd_sc_hd__mux2_1 _5636_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][58] ),
    .A1(_2903_),
    .S(net1000),
    .X(_0477_));
 sky130_fd_sc_hd__and2_1 _5637_ (.A(m1_wbd_adr_i[8]),
    .B(net1183),
    .X(_2904_));
 sky130_fd_sc_hd__a221o_1 _5638_ (.A1(net1239),
    .A2(m2_wbd_adr_i[8]),
    .B1(net1186),
    .B2(m3_wbd_adr_i[8]),
    .C1(net1192),
    .X(_2905_));
 sky130_fd_sc_hd__o22a_4 _5639_ (.A1(net2021),
    .A2(net1187),
    .B1(_2904_),
    .B2(_2905_),
    .X(_2906_));
 sky130_fd_sc_hd__mux2_1 _5640_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[3][59] ),
    .A1(_2906_),
    .S(net998),
    .X(_0478_));
 sky130_fd_sc_hd__o31a_1 _5641_ (.A1(m2_wbd_adr_i[17]),
    .A2(_1688_),
    .A3(_1775_),
    .B1(net1405),
    .X(_2907_));
 sky130_fd_sc_hd__a31o_1 _5642_ (.A1(m3_wbd_stb_i),
    .A2(net1182),
    .A3(_1853_),
    .B1(_2907_),
    .X(_2908_));
 sky130_fd_sc_hd__and2_1 _5643_ (.A(_1878_),
    .B(_2908_),
    .X(_2909_));
 sky130_fd_sc_hd__or3b_1 _5644_ (.A(_1690_),
    .B(net1183),
    .C_N(_1879_),
    .X(_2910_));
 sky130_fd_sc_hd__or2_1 _5645_ (.A(net1245),
    .B(_1878_),
    .X(_2911_));
 sky130_fd_sc_hd__a41o_1 _5646_ (.A1(m1_wbd_stb_i),
    .A2(_1834_),
    .A3(_1879_),
    .A4(_2911_),
    .B1(_2909_),
    .X(_2912_));
 sky130_fd_sc_hd__o31a_1 _5647_ (.A1(m2_wbd_adr_i[17]),
    .A2(_1688_),
    .A3(_1775_),
    .B1(net1245),
    .X(_2913_));
 sky130_fd_sc_hd__or2_1 _5648_ (.A(net1183),
    .B(_2913_),
    .X(_2914_));
 sky130_fd_sc_hd__a31o_1 _5649_ (.A1(m3_wbd_stb_i),
    .A2(_1853_),
    .A3(_2914_),
    .B1(_2912_),
    .X(_2915_));
 sky130_fd_sc_hd__nand2_2 _5650_ (.A(_1694_),
    .B(net630),
    .Y(_2916_));
 sky130_fd_sc_hd__mux2_1 _5651_ (.A0(net1405),
    .A1(_2915_),
    .S(_2916_),
    .X(_0479_));
 sky130_fd_sc_hd__o21ba_1 _5652_ (.A1(net1239),
    .A2(_1878_),
    .B1_N(_2913_),
    .X(_2917_));
 sky130_fd_sc_hd__a31o_1 _5653_ (.A1(m3_wbd_stb_i),
    .A2(_1853_),
    .A3(_2496_),
    .B1(_2917_),
    .X(_2918_));
 sky130_fd_sc_hd__and3_1 _5654_ (.A(_2910_),
    .B(_2911_),
    .C(_2918_),
    .X(_2919_));
 sky130_fd_sc_hd__mux2_1 _5655_ (.A0(\u_s1.gnt[1] ),
    .A1(_2919_),
    .S(_2916_),
    .X(_0480_));
 sky130_fd_sc_hd__nor2_4 _5656_ (.A(\u_s2.u_sync_wbb.m_state[1] ),
    .B(net1798),
    .Y(_2920_));
 sky130_fd_sc_hd__or2_4 _5657_ (.A(net1817),
    .B(net1798),
    .X(_2921_));
 sky130_fd_sc_hd__nand2_1 _5658_ (.A(_1691_),
    .B(net997),
    .Y(_2922_));
 sky130_fd_sc_hd__o21ai_2 _5659_ (.A1(_1691_),
    .A2(net583),
    .B1(_2922_),
    .Y(_2923_));
 sky130_fd_sc_hd__o21ai_1 _5660_ (.A1(_1989_),
    .A2(net996),
    .B1(_1984_),
    .Y(_2924_));
 sky130_fd_sc_hd__mux2_1 _5661_ (.A0(_2924_),
    .A1(\u_s2.u_sync_wbb.wbm_ack_o ),
    .S(_2923_),
    .X(_0481_));
 sky130_fd_sc_hd__nor2_1 _5662_ (.A(_1994_),
    .B(_2923_),
    .Y(_2925_));
 sky130_fd_sc_hd__nand2_1 _5663_ (.A(\u_s2.u_sync_wbb.m_state[1] ),
    .B(_1981_),
    .Y(_2926_));
 sky130_fd_sc_hd__o221a_1 _5664_ (.A1(\u_s2.u_sync_wbb.m_state[1] ),
    .A2(_1983_),
    .B1(_1988_),
    .B2(net1400),
    .C1(_2926_),
    .X(_2927_));
 sky130_fd_sc_hd__a31o_1 _5665_ (.A1(net726),
    .A2(_1971_),
    .A3(net997),
    .B1(_2927_),
    .X(_2928_));
 sky130_fd_sc_hd__mux2_1 _5666_ (.A0(\u_s2.u_sync_wbb.wbm_lack_o ),
    .A1(_2928_),
    .S(_2925_),
    .X(_0482_));
 sky130_fd_sc_hd__o21a_1 _5667_ (.A1(_1680_),
    .A2(_1981_),
    .B1(_2922_),
    .X(_2929_));
 sky130_fd_sc_hd__a21o_1 _5668_ (.A1(_1971_),
    .A2(net997),
    .B1(_1983_),
    .X(_2930_));
 sky130_fd_sc_hd__mux2_1 _5669_ (.A0(\u_s2.u_sync_wbb.m_cmd_wr_en ),
    .A1(_2930_),
    .S(net1818),
    .X(_0483_));
 sky130_fd_sc_hd__o21ai_2 _5670_ (.A1(_1680_),
    .A2(net1826),
    .B1(net1827),
    .Y(_2931_));
 sky130_fd_sc_hd__mux2_1 _5671_ (.A0(\u_s2.u_sync_wbb.m_resp_rd_en ),
    .A1(_1982_),
    .S(_2931_),
    .X(_0484_));
 sky130_fd_sc_hd__and2_1 _5672_ (.A(_1674_),
    .B(_2784_),
    .X(_2932_));
 sky130_fd_sc_hd__nor2_1 _5673_ (.A(_2786_),
    .B(_2932_),
    .Y(_0485_));
 sky130_fd_sc_hd__nor2_1 _5674_ (.A(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .B(_2786_),
    .Y(_2933_));
 sky130_fd_sc_hd__nor2_1 _5675_ (.A(net483),
    .B(_2933_),
    .Y(_0486_));
 sky130_fd_sc_hd__xor2_1 _5676_ (.A(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[2] ),
    .B(net484),
    .X(_0487_));
 sky130_fd_sc_hd__xor2_1 _5677_ (.A(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .B(\u_s2.u_sync_wbb.m_cmd_wr_en ),
    .X(_0488_));
 sky130_fd_sc_hd__and3_2 _5678_ (.A(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .B(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .C(\u_s2.u_sync_wbb.m_cmd_wr_en ),
    .X(_2934_));
 sky130_fd_sc_hd__a21oi_1 _5679_ (.A1(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .A2(\u_s2.u_sync_wbb.m_cmd_wr_en ),
    .B1(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .Y(_2935_));
 sky130_fd_sc_hd__nor2_1 _5680_ (.A(net993),
    .B(_2935_),
    .Y(_0489_));
 sky130_fd_sc_hd__xor2_1 _5681_ (.A(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[2] ),
    .B(net995),
    .X(_0490_));
 sky130_fd_sc_hd__or4_1 _5682_ (.A(_2570_),
    .B(_2571_),
    .C(net1816),
    .D(_2573_),
    .X(_2936_));
 sky130_fd_sc_hd__or4b_1 _5683_ (.A(_2568_),
    .B(_2936_),
    .C(_2569_),
    .D_N(net717),
    .X(_2937_));
 sky130_fd_sc_hd__or4_1 _5684_ (.A(net1804),
    .B(_2575_),
    .C(_2576_),
    .D(_2937_),
    .X(_2938_));
 sky130_fd_sc_hd__or4_1 _5685_ (.A(\u_s2.u_sync_wbb.s_cmd_rd_data_l[7] ),
    .B(\u_s2.u_sync_wbb.s_cmd_rd_data_l[6] ),
    .C(\u_s2.u_sync_wbb.s_cmd_rd_data_l[5] ),
    .D(\u_s2.u_sync_wbb.s_cmd_rd_data_l[4] ),
    .X(_2939_));
 sky130_fd_sc_hd__or4_1 _5686_ (.A(\u_s2.u_sync_wbb.s_cmd_rd_data_l[9] ),
    .B(\u_s2.u_sync_wbb.s_cmd_rd_data_l[8] ),
    .C(net717),
    .D(_2939_),
    .X(_2940_));
 sky130_fd_sc_hd__o41a_1 _5687_ (.A1(\u_s2.u_sync_wbb.s_cmd_rd_data_l[3] ),
    .A2(\u_s2.u_sync_wbb.s_cmd_rd_data_l[2] ),
    .A3(\u_s2.u_sync_wbb.s_cmd_rd_data_l[1] ),
    .A4(_2940_),
    .B1(_1710_),
    .X(_2941_));
 sky130_fd_sc_hd__a32o_1 _5688_ (.A1(net438),
    .A2(_2938_),
    .A3(_2941_),
    .B1(_1711_),
    .B2(\u_s2.u_sync_wbb.wbs_burst ),
    .X(_0491_));
 sky130_fd_sc_hd__xor2_1 _5689_ (.A(net1397),
    .B(net1501),
    .X(_0492_));
 sky130_fd_sc_hd__a21oi_1 _5690_ (.A1(net1397),
    .A2(net1501),
    .B1(net1391),
    .Y(_2942_));
 sky130_fd_sc_hd__and3_1 _5691_ (.A(net1390),
    .B(net1398),
    .C(net1501),
    .X(_2943_));
 sky130_fd_sc_hd__nor2_1 _5692_ (.A(_2942_),
    .B(_2943_),
    .Y(_0493_));
 sky130_fd_sc_hd__xor2_1 _5693_ (.A(\u_s2.u_sync_wbb.u_cmd_if.rd_ptr[2] ),
    .B(_2943_),
    .X(_0494_));
 sky130_fd_sc_hd__nor2_4 _5694_ (.A(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .B(_2799_),
    .Y(_2944_));
 sky130_fd_sc_hd__mux2_1 _5695_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][1] ),
    .A1(net797),
    .S(net751),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _5696_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][2] ),
    .A1(net798),
    .S(net749),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _5697_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][3] ),
    .A1(_1860_),
    .S(net751),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _5698_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][4] ),
    .A1(_1856_),
    .S(net750),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _5699_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][5] ),
    .A1(_1869_),
    .S(net754),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _5700_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][6] ),
    .A1(_1868_),
    .S(net752),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _5701_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][7] ),
    .A1(_1867_),
    .S(net749),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _5702_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][8] ),
    .A1(_1866_),
    .S(net751),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _5703_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][9] ),
    .A1(_1873_),
    .S(net749),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_1 _5704_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][14] ),
    .A1(net686),
    .S(net754),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _5705_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][15] ),
    .A1(net685),
    .S(net751),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _5706_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][16] ),
    .A1(net684),
    .S(net752),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _5707_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][17] ),
    .A1(net683),
    .S(net753),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _5708_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][18] ),
    .A1(net682),
    .S(net755),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _5709_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][19] ),
    .A1(_2816_),
    .S(net752),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _5710_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][20] ),
    .A1(_2818_),
    .S(net752),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _5711_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][21] ),
    .A1(net681),
    .S(net752),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _5712_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][22] ),
    .A1(_2823_),
    .S(net754),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _5713_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][23] ),
    .A1(_2825_),
    .S(net753),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _5714_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][24] ),
    .A1(_2827_),
    .S(net751),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _5715_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][25] ),
    .A1(_2830_),
    .S(net754),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _5716_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][26] ),
    .A1(_2832_),
    .S(net753),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _5717_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][27] ),
    .A1(_2835_),
    .S(net754),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _5718_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][28] ),
    .A1(_2838_),
    .S(net754),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _5719_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][29] ),
    .A1(_2841_),
    .S(net754),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_1 _5720_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][30] ),
    .A1(_2844_),
    .S(net754),
    .X(_0520_));
 sky130_fd_sc_hd__mux2_1 _5721_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][31] ),
    .A1(_2846_),
    .S(net751),
    .X(_0521_));
 sky130_fd_sc_hd__mux2_1 _5722_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][32] ),
    .A1(_2849_),
    .S(net752),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_1 _5723_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][33] ),
    .A1(_2851_),
    .S(net750),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_1 _5724_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][34] ),
    .A1(_2854_),
    .S(net752),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _5725_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][35] ),
    .A1(_2856_),
    .S(net754),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_1 _5726_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][36] ),
    .A1(_2858_),
    .S(net750),
    .X(_0526_));
 sky130_fd_sc_hd__mux2_1 _5727_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][37] ),
    .A1(_2861_),
    .S(net753),
    .X(_0527_));
 sky130_fd_sc_hd__mux2_1 _5728_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][38] ),
    .A1(_2863_),
    .S(net752),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_1 _5729_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][39] ),
    .A1(_2865_),
    .S(net749),
    .X(_0529_));
 sky130_fd_sc_hd__mux2_1 _5730_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][40] ),
    .A1(_2867_),
    .S(net750),
    .X(_0530_));
 sky130_fd_sc_hd__mux2_1 _5731_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][41] ),
    .A1(_2869_),
    .S(net751),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _5732_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][42] ),
    .A1(net680),
    .S(net752),
    .X(_0532_));
 sky130_fd_sc_hd__mux2_1 _5733_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][43] ),
    .A1(net2080),
    .S(net751),
    .X(_0533_));
 sky130_fd_sc_hd__mux2_1 _5734_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][44] ),
    .A1(_2875_),
    .S(net750),
    .X(_0534_));
 sky130_fd_sc_hd__mux2_1 _5735_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][45] ),
    .A1(_2877_),
    .S(net754),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_1 _5736_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][46] ),
    .A1(net679),
    .S(net755),
    .X(_0536_));
 sky130_fd_sc_hd__mux2_1 _5737_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][47] ),
    .A1(_2881_),
    .S(net749),
    .X(_0537_));
 sky130_fd_sc_hd__mux2_1 _5738_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][48] ),
    .A1(_2883_),
    .S(net749),
    .X(_0538_));
 sky130_fd_sc_hd__mux2_1 _5739_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][49] ),
    .A1(_2885_),
    .S(net750),
    .X(_0539_));
 sky130_fd_sc_hd__mux2_1 _5740_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][50] ),
    .A1(net732),
    .S(net753),
    .X(_0540_));
 sky130_fd_sc_hd__mux2_1 _5741_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][53] ),
    .A1(_2888_),
    .S(net749),
    .X(_0541_));
 sky130_fd_sc_hd__mux2_1 _5742_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][54] ),
    .A1(_2891_),
    .S(net750),
    .X(_0542_));
 sky130_fd_sc_hd__mux2_1 _5743_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][55] ),
    .A1(_2894_),
    .S(net749),
    .X(_0543_));
 sky130_fd_sc_hd__mux2_1 _5744_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][56] ),
    .A1(_2897_),
    .S(net751),
    .X(_0544_));
 sky130_fd_sc_hd__mux2_1 _5745_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][57] ),
    .A1(_2900_),
    .S(net749),
    .X(_0545_));
 sky130_fd_sc_hd__mux2_1 _5746_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][58] ),
    .A1(_2903_),
    .S(_2944_),
    .X(_0546_));
 sky130_fd_sc_hd__mux2_1 _5747_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[1][59] ),
    .A1(_2906_),
    .S(net749),
    .X(_0547_));
 sky130_fd_sc_hd__or3b_1 _5748_ (.A(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .B(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .C_N(\u_s0.u_sync_wbb.m_cmd_wr_en ),
    .X(_2945_));
 sky130_fd_sc_hd__mux2_1 _5749_ (.A0(_1786_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][0] ),
    .S(net985),
    .X(_0548_));
 sky130_fd_sc_hd__mux2_1 _5750_ (.A0(_1789_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][1] ),
    .S(net981),
    .X(_0549_));
 sky130_fd_sc_hd__mux2_1 _5751_ (.A0(_1792_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][2] ),
    .S(net987),
    .X(_0550_));
 sky130_fd_sc_hd__mux2_1 _5752_ (.A0(_1794_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][3] ),
    .S(net986),
    .X(_0551_));
 sky130_fd_sc_hd__mux2_1 _5753_ (.A0(_1793_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][4] ),
    .S(net986),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_1 _5754_ (.A0(net808),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][5] ),
    .S(net987),
    .X(_0553_));
 sky130_fd_sc_hd__mux2_1 _5755_ (.A0(_1797_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][6] ),
    .S(net987),
    .X(_0554_));
 sky130_fd_sc_hd__mux2_1 _5756_ (.A0(_1796_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][7] ),
    .S(net987),
    .X(_0555_));
 sky130_fd_sc_hd__mux2_1 _5757_ (.A0(_1799_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][8] ),
    .S(net987),
    .X(_0556_));
 sky130_fd_sc_hd__mux2_1 _5758_ (.A0(_1787_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][9] ),
    .S(net985),
    .X(_0557_));
 sky130_fd_sc_hd__and3_1 _5759_ (.A(net1371),
    .B(net1375),
    .C(m3_wbd_sel_i[0]),
    .X(_2946_));
 sky130_fd_sc_hd__a221o_1 _5760_ (.A1(net1259),
    .A2(net2082),
    .B1(net2085),
    .B2(net823),
    .C1(net1205),
    .X(_2947_));
 sky130_fd_sc_hd__o22a_2 _5761_ (.A1(net1565),
    .A2(net1199),
    .B1(_2946_),
    .B2(_2947_),
    .X(_2948_));
 sky130_fd_sc_hd__mux2_1 _5762_ (.A0(_2948_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][14] ),
    .S(net983),
    .X(_0558_));
 sky130_fd_sc_hd__a221o_2 _5763_ (.A1(net1259),
    .A2(m2_wbd_sel_i[1]),
    .B1(net1208),
    .B2(m3_wbd_sel_i[1]),
    .C1(net1204),
    .X(_2949_));
 sky130_fd_sc_hd__a21o_1 _5764_ (.A1(m1_wbd_sel_i[1]),
    .A2(net823),
    .B1(_2949_),
    .X(_2950_));
 sky130_fd_sc_hd__o21a_1 _5765_ (.A1(net2030),
    .A2(net1196),
    .B1(_2950_),
    .X(_2951_));
 sky130_fd_sc_hd__mux2_1 _5766_ (.A0(_2951_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][15] ),
    .S(net988),
    .X(_0559_));
 sky130_fd_sc_hd__a221o_2 _5767_ (.A1(net1259),
    .A2(m2_wbd_sel_i[2]),
    .B1(net1206),
    .B2(m3_wbd_sel_i[2]),
    .C1(net1205),
    .X(_2952_));
 sky130_fd_sc_hd__a21o_1 _5768_ (.A1(m1_wbd_sel_i[2]),
    .A2(net823),
    .B1(_2952_),
    .X(_2953_));
 sky130_fd_sc_hd__o21a_2 _5769_ (.A1(net2046),
    .A2(net1195),
    .B1(_2953_),
    .X(_2954_));
 sky130_fd_sc_hd__mux2_1 _5770_ (.A0(_2954_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][16] ),
    .S(net980),
    .X(_0560_));
 sky130_fd_sc_hd__a221o_2 _5771_ (.A1(net1259),
    .A2(m2_wbd_sel_i[3]),
    .B1(net1206),
    .B2(m3_wbd_sel_i[3]),
    .C1(net1205),
    .X(_2955_));
 sky130_fd_sc_hd__a21o_1 _5772_ (.A1(m1_wbd_sel_i[3]),
    .A2(net823),
    .B1(_2955_),
    .X(_2956_));
 sky130_fd_sc_hd__o21a_2 _5773_ (.A1(net2027),
    .A2(net1196),
    .B1(_2956_),
    .X(_2957_));
 sky130_fd_sc_hd__mux2_1 _5774_ (.A0(_2957_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][17] ),
    .S(net980),
    .X(_0561_));
 sky130_fd_sc_hd__or2_1 _5775_ (.A(net1593),
    .B(net1201),
    .X(_2958_));
 sky130_fd_sc_hd__a21o_1 _5776_ (.A1(net1262),
    .A2(m2_wbd_dat_i[0]),
    .B1(net1272),
    .X(_2959_));
 sky130_fd_sc_hd__o211a_1 _5777_ (.A1(net1262),
    .A2(net1562),
    .B1(_2958_),
    .C1(_2959_),
    .X(_2960_));
 sky130_fd_sc_hd__mux2_1 _5778_ (.A0(_2960_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][18] ),
    .S(net987),
    .X(_0562_));
 sky130_fd_sc_hd__a21o_1 _5779_ (.A1(net1273),
    .A2(net1551),
    .B1(net1263),
    .X(_2961_));
 sky130_fd_sc_hd__o221a_1 _5780_ (.A1(net1273),
    .A2(m2_wbd_dat_i[1]),
    .B1(net1582),
    .B2(net1201),
    .C1(_2961_),
    .X(_2962_));
 sky130_fd_sc_hd__mux2_1 _5781_ (.A0(_2962_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][19] ),
    .S(net986),
    .X(_0563_));
 sky130_fd_sc_hd__a21o_1 _5782_ (.A1(net1272),
    .A2(net1543),
    .B1(net1262),
    .X(_2963_));
 sky130_fd_sc_hd__o221a_2 _5783_ (.A1(net1273),
    .A2(m2_wbd_dat_i[2]),
    .B1(net1574),
    .B2(net1201),
    .C1(_2963_),
    .X(_2964_));
 sky130_fd_sc_hd__mux2_1 _5784_ (.A0(_2964_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][20] ),
    .S(net987),
    .X(_0564_));
 sky130_fd_sc_hd__a21o_1 _5785_ (.A1(net1270),
    .A2(m1_wbd_dat_i[3]),
    .B1(net1261),
    .X(_2965_));
 sky130_fd_sc_hd__o221a_2 _5786_ (.A1(net1270),
    .A2(net2088),
    .B1(m0_wbd_dat_i[3]),
    .B2(net1200),
    .C1(_2965_),
    .X(_2966_));
 sky130_fd_sc_hd__mux2_1 _5787_ (.A0(_2966_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][21] ),
    .S(net986),
    .X(_0565_));
 sky130_fd_sc_hd__or2_1 _5788_ (.A(m0_wbd_dat_i[4]),
    .B(net1199),
    .X(_2967_));
 sky130_fd_sc_hd__a21o_1 _5789_ (.A1(net1260),
    .A2(m2_wbd_dat_i[4]),
    .B1(net1269),
    .X(_2968_));
 sky130_fd_sc_hd__o211a_1 _5790_ (.A1(net1260),
    .A2(net2006),
    .B1(_2967_),
    .C1(_2968_),
    .X(_2969_));
 sky130_fd_sc_hd__mux2_1 _5791_ (.A0(_2969_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][22] ),
    .S(net984),
    .X(_0566_));
 sky130_fd_sc_hd__a21o_1 _5792_ (.A1(net1273),
    .A2(net1539),
    .B1(net1262),
    .X(_2970_));
 sky130_fd_sc_hd__o221a_1 _5793_ (.A1(net1273),
    .A2(net1517),
    .B1(net1570),
    .B2(net1201),
    .C1(_2970_),
    .X(_2971_));
 sky130_fd_sc_hd__mux2_1 _5794_ (.A0(_2971_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][23] ),
    .S(net984),
    .X(_0567_));
 sky130_fd_sc_hd__a21o_1 _5795_ (.A1(net1270),
    .A2(net1538),
    .B1(net1261),
    .X(_2972_));
 sky130_fd_sc_hd__o221a_1 _5796_ (.A1(net1270),
    .A2(net1516),
    .B1(net1569),
    .B2(_1730_),
    .C1(_2972_),
    .X(_2973_));
 sky130_fd_sc_hd__mux2_1 _5797_ (.A0(_2973_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][24] ),
    .S(net986),
    .X(_0568_));
 sky130_fd_sc_hd__or2_1 _5798_ (.A(m0_wbd_dat_i[7]),
    .B(net1197),
    .X(_2974_));
 sky130_fd_sc_hd__a21o_1 _5799_ (.A1(net1255),
    .A2(m2_wbd_dat_i[7]),
    .B1(net1265),
    .X(_2975_));
 sky130_fd_sc_hd__o211a_1 _5800_ (.A1(net1255),
    .A2(net2084),
    .B1(_2974_),
    .C1(_2975_),
    .X(_2976_));
 sky130_fd_sc_hd__mux2_1 _5801_ (.A0(_2976_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][25] ),
    .S(net984),
    .X(_0569_));
 sky130_fd_sc_hd__or2_1 _5802_ (.A(m0_wbd_dat_i[8]),
    .B(net1200),
    .X(_2977_));
 sky130_fd_sc_hd__a21o_1 _5803_ (.A1(net1261),
    .A2(m2_wbd_dat_i[8]),
    .B1(net1270),
    .X(_2978_));
 sky130_fd_sc_hd__o211a_1 _5804_ (.A1(net1261),
    .A2(net2077),
    .B1(_2977_),
    .C1(_2978_),
    .X(_2979_));
 sky130_fd_sc_hd__mux2_1 _5805_ (.A0(_2979_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][26] ),
    .S(net984),
    .X(_0570_));
 sky130_fd_sc_hd__a21o_1 _5806_ (.A1(net1272),
    .A2(net1535),
    .B1(net1262),
    .X(_2980_));
 sky130_fd_sc_hd__o221a_1 _5807_ (.A1(net1272),
    .A2(net1513),
    .B1(net1566),
    .B2(net1201),
    .C1(_2980_),
    .X(_2981_));
 sky130_fd_sc_hd__mux2_1 _5808_ (.A0(_2981_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][27] ),
    .S(net986),
    .X(_0571_));
 sky130_fd_sc_hd__a21o_1 _5809_ (.A1(net1272),
    .A2(net1561),
    .B1(net1262),
    .X(_2982_));
 sky130_fd_sc_hd__o221a_1 _5810_ (.A1(net1272),
    .A2(net1534),
    .B1(net1592),
    .B2(net1201),
    .C1(_2982_),
    .X(_2983_));
 sky130_fd_sc_hd__mux2_1 _5811_ (.A0(_2983_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][28] ),
    .S(net986),
    .X(_0572_));
 sky130_fd_sc_hd__a21o_1 _5812_ (.A1(net1272),
    .A2(net1560),
    .B1(net1262),
    .X(_2984_));
 sky130_fd_sc_hd__o221a_1 _5813_ (.A1(net1272),
    .A2(net1533),
    .B1(net1591),
    .B2(net1201),
    .C1(_2984_),
    .X(_2985_));
 sky130_fd_sc_hd__mux2_1 _5814_ (.A0(_2985_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][29] ),
    .S(net986),
    .X(_0573_));
 sky130_fd_sc_hd__or2_1 _5815_ (.A(m0_wbd_dat_i[12]),
    .B(net1197),
    .X(_2986_));
 sky130_fd_sc_hd__a21o_1 _5816_ (.A1(net1257),
    .A2(m2_wbd_dat_i[12]),
    .B1(net1267),
    .X(_2987_));
 sky130_fd_sc_hd__o211a_1 _5817_ (.A1(net1257),
    .A2(net2055),
    .B1(_2986_),
    .C1(_2987_),
    .X(_2988_));
 sky130_fd_sc_hd__mux2_1 _5818_ (.A0(_2988_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][30] ),
    .S(net980),
    .X(_0574_));
 sky130_fd_sc_hd__or2_1 _5819_ (.A(net1589),
    .B(net1198),
    .X(_2989_));
 sky130_fd_sc_hd__a21o_1 _5820_ (.A1(net1256),
    .A2(m2_wbd_dat_i[13]),
    .B1(net1266),
    .X(_2990_));
 sky130_fd_sc_hd__o211a_1 _5821_ (.A1(net1255),
    .A2(net1558),
    .B1(_2989_),
    .C1(_2990_),
    .X(_2991_));
 sky130_fd_sc_hd__mux2_1 _5822_ (.A0(_2991_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][31] ),
    .S(net983),
    .X(_0575_));
 sky130_fd_sc_hd__a21o_1 _5823_ (.A1(net1272),
    .A2(net1557),
    .B1(net1262),
    .X(_2992_));
 sky130_fd_sc_hd__o221a_1 _5824_ (.A1(net1272),
    .A2(net1531),
    .B1(net1588),
    .B2(net1201),
    .C1(_2992_),
    .X(_2993_));
 sky130_fd_sc_hd__mux2_1 _5825_ (.A0(_2993_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][32] ),
    .S(net986),
    .X(_0576_));
 sky130_fd_sc_hd__a21o_1 _5826_ (.A1(net1265),
    .A2(net1556),
    .B1(net1260),
    .X(_2994_));
 sky130_fd_sc_hd__o221a_1 _5827_ (.A1(net1266),
    .A2(net2036),
    .B1(net1587),
    .B2(net1199),
    .C1(_2994_),
    .X(_2995_));
 sky130_fd_sc_hd__mux2_1 _5828_ (.A0(_2995_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][33] ),
    .S(net984),
    .X(_0577_));
 sky130_fd_sc_hd__or2_1 _5829_ (.A(m0_wbd_dat_i[16]),
    .B(net1199),
    .X(_2996_));
 sky130_fd_sc_hd__a21o_1 _5830_ (.A1(net1255),
    .A2(m2_wbd_dat_i[16]),
    .B1(net1265),
    .X(_2997_));
 sky130_fd_sc_hd__o211a_2 _5831_ (.A1(net1255),
    .A2(net2039),
    .B1(_2996_),
    .C1(_2997_),
    .X(_2998_));
 sky130_fd_sc_hd__mux2_1 _5832_ (.A0(_2998_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][34] ),
    .S(net983),
    .X(_0578_));
 sky130_fd_sc_hd__or2_1 _5833_ (.A(net1585),
    .B(net1200),
    .X(_2999_));
 sky130_fd_sc_hd__a21o_1 _5834_ (.A1(net1261),
    .A2(net1528),
    .B1(net1270),
    .X(_3000_));
 sky130_fd_sc_hd__o211a_1 _5835_ (.A1(net1261),
    .A2(net1554),
    .B1(_2999_),
    .C1(_3000_),
    .X(_3001_));
 sky130_fd_sc_hd__mux2_1 _5836_ (.A0(_3001_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][35] ),
    .S(net986),
    .X(_0579_));
 sky130_fd_sc_hd__or2_1 _5837_ (.A(net1584),
    .B(net1197),
    .X(_3002_));
 sky130_fd_sc_hd__a21o_1 _5838_ (.A1(net1255),
    .A2(m2_wbd_dat_i[18]),
    .B1(net1265),
    .X(_3003_));
 sky130_fd_sc_hd__o211a_1 _5839_ (.A1(net1257),
    .A2(net1553),
    .B1(_3002_),
    .C1(_3003_),
    .X(_3004_));
 sky130_fd_sc_hd__mux2_1 _5840_ (.A0(_3004_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][36] ),
    .S(net980),
    .X(_0580_));
 sky130_fd_sc_hd__or2_1 _5841_ (.A(net1583),
    .B(net1200),
    .X(_3005_));
 sky130_fd_sc_hd__a21o_1 _5842_ (.A1(net1260),
    .A2(m2_wbd_dat_i[19]),
    .B1(net1269),
    .X(_3006_));
 sky130_fd_sc_hd__o211a_1 _5843_ (.A1(net1260),
    .A2(net2008),
    .B1(_3005_),
    .C1(_3006_),
    .X(_3007_));
 sky130_fd_sc_hd__mux2_1 _5844_ (.A0(net2009),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][37] ),
    .S(net984),
    .X(_0581_));
 sky130_fd_sc_hd__or2_1 _5845_ (.A(m0_wbd_dat_i[20]),
    .B(net1197),
    .X(_3008_));
 sky130_fd_sc_hd__a21o_1 _5846_ (.A1(net1255),
    .A2(m2_wbd_dat_i[20]),
    .B1(net1265),
    .X(_3009_));
 sky130_fd_sc_hd__o211a_2 _5847_ (.A1(net1255),
    .A2(net2064),
    .B1(_3008_),
    .C1(_3009_),
    .X(_3010_));
 sky130_fd_sc_hd__mux2_1 _5848_ (.A0(_3010_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][38] ),
    .S(net980),
    .X(_0582_));
 sky130_fd_sc_hd__a21o_1 _5849_ (.A1(net1269),
    .A2(net1549),
    .B1(net1260),
    .X(_3011_));
 sky130_fd_sc_hd__o221a_1 _5850_ (.A1(net1269),
    .A2(net1525),
    .B1(net1580),
    .B2(net1200),
    .C1(_3011_),
    .X(_3012_));
 sky130_fd_sc_hd__mux2_1 _5851_ (.A0(_3012_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][39] ),
    .S(net984),
    .X(_0583_));
 sky130_fd_sc_hd__a21o_1 _5852_ (.A1(net1265),
    .A2(net1548),
    .B1(net1256),
    .X(_3013_));
 sky130_fd_sc_hd__o221a_2 _5853_ (.A1(net1266),
    .A2(net2051),
    .B1(net1579),
    .B2(net1198),
    .C1(_3013_),
    .X(_3014_));
 sky130_fd_sc_hd__mux2_1 _5854_ (.A0(_3014_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][40] ),
    .S(net983),
    .X(_0584_));
 sky130_fd_sc_hd__a21o_1 _5855_ (.A1(net1269),
    .A2(net1547),
    .B1(net1260),
    .X(_3015_));
 sky130_fd_sc_hd__o221a_2 _5856_ (.A1(net1269),
    .A2(net1524),
    .B1(net1578),
    .B2(net1199),
    .C1(_3015_),
    .X(_3016_));
 sky130_fd_sc_hd__mux2_1 _5857_ (.A0(_3016_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][41] ),
    .S(net985),
    .X(_0585_));
 sky130_fd_sc_hd__or2_1 _5858_ (.A(m0_wbd_dat_i[24]),
    .B(net1197),
    .X(_3017_));
 sky130_fd_sc_hd__a21o_1 _5859_ (.A1(net1256),
    .A2(m2_wbd_dat_i[24]),
    .B1(net1266),
    .X(_3018_));
 sky130_fd_sc_hd__o211a_1 _5860_ (.A1(net1256),
    .A2(net2016),
    .B1(_3017_),
    .C1(_3018_),
    .X(_3019_));
 sky130_fd_sc_hd__mux2_1 _5861_ (.A0(net2017),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][42] ),
    .S(net983),
    .X(_0586_));
 sky130_fd_sc_hd__or2_1 _5862_ (.A(m0_wbd_dat_i[25]),
    .B(net1200),
    .X(_3020_));
 sky130_fd_sc_hd__a21o_1 _5863_ (.A1(net1260),
    .A2(m2_wbd_dat_i[25]),
    .B1(net1269),
    .X(_3021_));
 sky130_fd_sc_hd__o211a_1 _5864_ (.A1(net1260),
    .A2(net2037),
    .B1(_3020_),
    .C1(_3021_),
    .X(_3022_));
 sky130_fd_sc_hd__mux2_1 _5865_ (.A0(net2038),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][43] ),
    .S(net984),
    .X(_0587_));
 sky130_fd_sc_hd__a21o_1 _5866_ (.A1(net1265),
    .A2(m1_wbd_dat_i[26]),
    .B1(net1255),
    .X(_3023_));
 sky130_fd_sc_hd__o221a_1 _5867_ (.A1(net1265),
    .A2(net2067),
    .B1(net2018),
    .B2(net1198),
    .C1(_3023_),
    .X(_3024_));
 sky130_fd_sc_hd__mux2_1 _5868_ (.A0(_3024_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][44] ),
    .S(net983),
    .X(_0588_));
 sky130_fd_sc_hd__a21o_1 _5869_ (.A1(net1267),
    .A2(net2043),
    .B1(net1257),
    .X(_3025_));
 sky130_fd_sc_hd__o221a_1 _5870_ (.A1(net1267),
    .A2(net2041),
    .B1(net2010),
    .B2(net1197),
    .C1(_3025_),
    .X(_3026_));
 sky130_fd_sc_hd__mux2_1 _5871_ (.A0(_3026_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][45] ),
    .S(net988),
    .X(_0589_));
 sky130_fd_sc_hd__or2_1 _5872_ (.A(m0_wbd_dat_i[28]),
    .B(net1197),
    .X(_3027_));
 sky130_fd_sc_hd__a21o_1 _5873_ (.A1(net1257),
    .A2(m2_wbd_dat_i[28]),
    .B1(net1267),
    .X(_3028_));
 sky130_fd_sc_hd__o211a_2 _5874_ (.A1(net1257),
    .A2(net2091),
    .B1(_3027_),
    .C1(_3028_),
    .X(_3029_));
 sky130_fd_sc_hd__mux2_1 _5875_ (.A0(_3029_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][46] ),
    .S(net980),
    .X(_0590_));
 sky130_fd_sc_hd__a21o_1 _5876_ (.A1(net1265),
    .A2(m1_wbd_dat_i[29]),
    .B1(net1255),
    .X(_3030_));
 sky130_fd_sc_hd__o221a_1 _5877_ (.A1(net1265),
    .A2(net2061),
    .B1(net1575),
    .B2(net1199),
    .C1(_3030_),
    .X(_3031_));
 sky130_fd_sc_hd__mux2_1 _5878_ (.A0(_3031_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][47] ),
    .S(net983),
    .X(_0591_));
 sky130_fd_sc_hd__a21o_1 _5879_ (.A1(net1269),
    .A2(net1542),
    .B1(net1260),
    .X(_3032_));
 sky130_fd_sc_hd__o221a_1 _5880_ (.A1(net1269),
    .A2(net1520),
    .B1(net1573),
    .B2(net1199),
    .C1(_3032_),
    .X(_3033_));
 sky130_fd_sc_hd__mux2_1 _5881_ (.A0(_3033_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][48] ),
    .S(net984),
    .X(_0592_));
 sky130_fd_sc_hd__a21o_1 _5882_ (.A1(net1268),
    .A2(m1_wbd_dat_i[31]),
    .B1(_1670_),
    .X(_3034_));
 sky130_fd_sc_hd__o221a_1 _5883_ (.A1(net1268),
    .A2(m2_wbd_dat_i[31]),
    .B1(net2057),
    .B2(net1196),
    .C1(_3034_),
    .X(_3035_));
 sky130_fd_sc_hd__mux2_1 _5884_ (.A0(net2058),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][49] ),
    .S(net981),
    .X(_0593_));
 sky130_fd_sc_hd__mux2_1 _5885_ (.A0(_1806_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][50] ),
    .S(net984),
    .X(_0594_));
 sky130_fd_sc_hd__and3_1 _5886_ (.A(net1371),
    .B(net1375),
    .C(m3_wbd_adr_i[2]),
    .X(_3036_));
 sky130_fd_sc_hd__a221o_1 _5887_ (.A1(net1258),
    .A2(m2_wbd_adr_i[2]),
    .B1(m1_wbd_adr_i[2]),
    .B2(net823),
    .C1(net1204),
    .X(_3037_));
 sky130_fd_sc_hd__o22a_1 _5888_ (.A1(net1598),
    .A2(net1197),
    .B1(_3036_),
    .B2(_3037_),
    .X(_3038_));
 sky130_fd_sc_hd__mux2_1 _5889_ (.A0(_3038_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][53] ),
    .S(net985),
    .X(_0595_));
 sky130_fd_sc_hd__and3_1 _5890_ (.A(net1271),
    .B(net1375),
    .C(m1_wbd_adr_i[3]),
    .X(_3039_));
 sky130_fd_sc_hd__a221o_1 _5891_ (.A1(net1263),
    .A2(m2_wbd_adr_i[3]),
    .B1(net1208),
    .B2(m3_wbd_adr_i[3]),
    .C1(net1205),
    .X(_3040_));
 sky130_fd_sc_hd__o22a_2 _5892_ (.A1(net1597),
    .A2(net1199),
    .B1(_3039_),
    .B2(_3040_),
    .X(_3041_));
 sky130_fd_sc_hd__mux2_1 _5893_ (.A0(_3041_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][54] ),
    .S(net983),
    .X(_0596_));
 sky130_fd_sc_hd__and3_1 _5894_ (.A(net1271),
    .B(net1375),
    .C(m1_wbd_adr_i[4]),
    .X(_3042_));
 sky130_fd_sc_hd__a221o_1 _5895_ (.A1(net1259),
    .A2(m2_wbd_adr_i[4]),
    .B1(net1208),
    .B2(m3_wbd_adr_i[4]),
    .C1(net1204),
    .X(_3043_));
 sky130_fd_sc_hd__o22a_1 _5896_ (.A1(net1596),
    .A2(net1199),
    .B1(_3042_),
    .B2(_3043_),
    .X(_3044_));
 sky130_fd_sc_hd__mux2_1 _5897_ (.A0(_3044_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][55] ),
    .S(net982),
    .X(_0597_));
 sky130_fd_sc_hd__and3_1 _5898_ (.A(net1270),
    .B(net1375),
    .C(m1_wbd_adr_i[5]),
    .X(_3045_));
 sky130_fd_sc_hd__a221o_1 _5899_ (.A1(net1262),
    .A2(m2_wbd_adr_i[5]),
    .B1(net1207),
    .B2(m3_wbd_adr_i[5]),
    .C1(net1205),
    .X(_3046_));
 sky130_fd_sc_hd__o22a_2 _5900_ (.A1(net1595),
    .A2(net1201),
    .B1(_3045_),
    .B2(_3046_),
    .X(_3047_));
 sky130_fd_sc_hd__mux2_1 _5901_ (.A0(_3047_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][56] ),
    .S(net982),
    .X(_0598_));
 sky130_fd_sc_hd__a221o_1 _5902_ (.A1(net1259),
    .A2(m2_wbd_adr_i[6]),
    .B1(net1208),
    .B2(m3_wbd_adr_i[6]),
    .C1(_1729_),
    .X(_3048_));
 sky130_fd_sc_hd__a21o_1 _5903_ (.A1(net1983),
    .A2(_1724_),
    .B1(_3048_),
    .X(_3049_));
 sky130_fd_sc_hd__o21a_2 _5904_ (.A1(net1832),
    .A2(net1198),
    .B1(_3049_),
    .X(_3050_));
 sky130_fd_sc_hd__mux2_1 _5905_ (.A0(_3050_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][57] ),
    .S(net980),
    .X(_0599_));
 sky130_fd_sc_hd__a221o_4 _5906_ (.A1(net1261),
    .A2(m2_wbd_adr_i[7]),
    .B1(net1208),
    .B2(m3_wbd_adr_i[7]),
    .C1(net1205),
    .X(_3051_));
 sky130_fd_sc_hd__a21o_1 _5907_ (.A1(m1_wbd_adr_i[7]),
    .A2(net822),
    .B1(_3051_),
    .X(_3052_));
 sky130_fd_sc_hd__o21a_1 _5908_ (.A1(net1594),
    .A2(net1194),
    .B1(_3052_),
    .X(_3053_));
 sky130_fd_sc_hd__mux2_1 _5909_ (.A0(_3053_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][58] ),
    .S(net980),
    .X(_0600_));
 sky130_fd_sc_hd__and3_1 _5910_ (.A(net1269),
    .B(net1375),
    .C(m1_wbd_adr_i[8]),
    .X(_3054_));
 sky130_fd_sc_hd__a221o_1 _5911_ (.A1(net1261),
    .A2(m2_wbd_adr_i[8]),
    .B1(net1208),
    .B2(m3_wbd_adr_i[8]),
    .C1(net1205),
    .X(_3055_));
 sky130_fd_sc_hd__o22a_2 _5912_ (.A1(net2021),
    .A2(net1200),
    .B1(_3054_),
    .B2(_3055_),
    .X(_3056_));
 sky130_fd_sc_hd__mux2_1 _5913_ (.A0(net2022),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][59] ),
    .S(net982),
    .X(_0601_));
 sky130_fd_sc_hd__and3_1 _5914_ (.A(net1268),
    .B(net1374),
    .C(m1_wbd_adr_i[9]),
    .X(_3057_));
 sky130_fd_sc_hd__a221o_1 _5915_ (.A1(net1258),
    .A2(m2_wbd_adr_i[9]),
    .B1(net1206),
    .B2(m3_wbd_adr_i[9]),
    .C1(net1204),
    .X(_3058_));
 sky130_fd_sc_hd__o22a_1 _5916_ (.A1(net2031),
    .A2(net1197),
    .B1(_3057_),
    .B2(_3058_),
    .X(_3059_));
 sky130_fd_sc_hd__mux2_1 _5917_ (.A0(_3059_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][60] ),
    .S(net982),
    .X(_0602_));
 sky130_fd_sc_hd__and3_1 _5918_ (.A(net1370),
    .B(net1374),
    .C(m3_wbd_adr_i[10]),
    .X(_3060_));
 sky130_fd_sc_hd__a221o_1 _5919_ (.A1(net1258),
    .A2(m2_wbd_adr_i[10]),
    .B1(m1_wbd_adr_i[10]),
    .B2(net823),
    .C1(net1204),
    .X(_3061_));
 sky130_fd_sc_hd__o22a_1 _5920_ (.A1(m0_wbd_adr_i[10]),
    .A2(net1197),
    .B1(_3060_),
    .B2(_3061_),
    .X(_3062_));
 sky130_fd_sc_hd__mux2_1 _5921_ (.A0(_3062_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][61] ),
    .S(net983),
    .X(_0603_));
 sky130_fd_sc_hd__o21a_1 _5922_ (.A1(net1264),
    .A2(m2_wbd_adr_i[11]),
    .B1(net1254),
    .X(_3063_));
 sky130_fd_sc_hd__a22o_1 _5923_ (.A1(net1264),
    .A2(m1_wbd_adr_i[11]),
    .B1(net1206),
    .B2(m3_wbd_adr_i[11]),
    .X(_3064_));
 sky130_fd_sc_hd__o22a_1 _5924_ (.A1(m0_wbd_adr_i[11]),
    .A2(net1196),
    .B1(_3063_),
    .B2(_3064_),
    .X(_3065_));
 sky130_fd_sc_hd__mux2_1 _5925_ (.A0(_3065_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][62] ),
    .S(net979),
    .X(_0604_));
 sky130_fd_sc_hd__o21a_1 _5926_ (.A1(net1264),
    .A2(m2_wbd_adr_i[12]),
    .B1(net1254),
    .X(_3066_));
 sky130_fd_sc_hd__a22o_1 _5927_ (.A1(net1264),
    .A2(m1_wbd_adr_i[12]),
    .B1(net1206),
    .B2(m3_wbd_adr_i[12]),
    .X(_3067_));
 sky130_fd_sc_hd__o22a_1 _5928_ (.A1(m0_wbd_adr_i[12]),
    .A2(net1196),
    .B1(_3066_),
    .B2(_3067_),
    .X(_3068_));
 sky130_fd_sc_hd__mux2_1 _5929_ (.A0(_3068_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][63] ),
    .S(net982),
    .X(_0605_));
 sky130_fd_sc_hd__o21a_1 _5930_ (.A1(net1264),
    .A2(m2_wbd_adr_i[13]),
    .B1(net1258),
    .X(_3069_));
 sky130_fd_sc_hd__a22o_1 _5931_ (.A1(net1268),
    .A2(m1_wbd_adr_i[13]),
    .B1(net1206),
    .B2(m3_wbd_adr_i[13]),
    .X(_3070_));
 sky130_fd_sc_hd__o22a_1 _5932_ (.A1(net1908),
    .A2(net1196),
    .B1(_3069_),
    .B2(_3070_),
    .X(_3071_));
 sky130_fd_sc_hd__mux2_1 _5933_ (.A0(_3071_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][64] ),
    .S(net982),
    .X(_0606_));
 sky130_fd_sc_hd__o21a_1 _5934_ (.A1(net1264),
    .A2(net1997),
    .B1(net1253),
    .X(_3072_));
 sky130_fd_sc_hd__a22o_1 _5935_ (.A1(net1264),
    .A2(m1_wbd_adr_i[14]),
    .B1(net1206),
    .B2(m3_wbd_adr_i[14]),
    .X(_3073_));
 sky130_fd_sc_hd__o22a_1 _5936_ (.A1(net1858),
    .A2(net1194),
    .B1(_3072_),
    .B2(_3073_),
    .X(_3074_));
 sky130_fd_sc_hd__mux2_1 _5937_ (.A0(net1998),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][65] ),
    .S(net979),
    .X(_0607_));
 sky130_fd_sc_hd__o21a_1 _5938_ (.A1(net1264),
    .A2(m2_wbd_adr_i[15]),
    .B1(net1254),
    .X(_3075_));
 sky130_fd_sc_hd__a22o_1 _5939_ (.A1(net1264),
    .A2(m1_wbd_adr_i[15]),
    .B1(net1206),
    .B2(m3_wbd_adr_i[15]),
    .X(_3076_));
 sky130_fd_sc_hd__o22a_1 _5940_ (.A1(net1868),
    .A2(net1195),
    .B1(_3075_),
    .B2(_3076_),
    .X(_3077_));
 sky130_fd_sc_hd__mux2_1 _5941_ (.A0(_3077_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][66] ),
    .S(net979),
    .X(_0608_));
 sky130_fd_sc_hd__a221o_2 _5942_ (.A1(net1258),
    .A2(m2_wbd_adr_i[16]),
    .B1(net1209),
    .B2(m3_wbd_adr_i[16]),
    .C1(net1204),
    .X(_3078_));
 sky130_fd_sc_hd__a21oi_2 _5943_ (.A1(m1_wbd_adr_i[16]),
    .A2(net822),
    .B1(_3078_),
    .Y(_3079_));
 sky130_fd_sc_hd__a21oi_2 _5944_ (.A1(_1685_),
    .A2(net1203),
    .B1(_3079_),
    .Y(_3080_));
 sky130_fd_sc_hd__mux2_1 _5945_ (.A0(_3080_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][67] ),
    .S(net982),
    .X(_0609_));
 sky130_fd_sc_hd__a221o_2 _5946_ (.A1(net1259),
    .A2(m2_wbd_adr_i[17]),
    .B1(net1209),
    .B2(m3_wbd_adr_i[17]),
    .C1(net1204),
    .X(_3081_));
 sky130_fd_sc_hd__a21oi_2 _5947_ (.A1(m1_wbd_adr_i[17]),
    .A2(net822),
    .B1(_3081_),
    .Y(_3082_));
 sky130_fd_sc_hd__a21oi_2 _5948_ (.A1(_1684_),
    .A2(net1203),
    .B1(_3082_),
    .Y(_3083_));
 sky130_fd_sc_hd__mux2_1 _5949_ (.A0(_3083_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][68] ),
    .S(net982),
    .X(_0610_));
 sky130_fd_sc_hd__and3_1 _5950_ (.A(net1368),
    .B(net1372),
    .C(m3_wbd_adr_i[18]),
    .X(_3084_));
 sky130_fd_sc_hd__a221o_1 _5951_ (.A1(net1253),
    .A2(m2_wbd_adr_i[18]),
    .B1(net2004),
    .B2(net821),
    .C1(net1202),
    .X(_3085_));
 sky130_fd_sc_hd__o22a_1 _5952_ (.A1(net1854),
    .A2(net1194),
    .B1(_3084_),
    .B2(net2005),
    .X(_3086_));
 sky130_fd_sc_hd__mux2_1 _5953_ (.A0(_3086_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][69] ),
    .S(net979),
    .X(_0611_));
 sky130_fd_sc_hd__a221o_2 _5954_ (.A1(net1259),
    .A2(m2_wbd_adr_i[19]),
    .B1(net1206),
    .B2(m3_wbd_adr_i[19]),
    .C1(net1205),
    .X(_3087_));
 sky130_fd_sc_hd__a21o_1 _5955_ (.A1(net1995),
    .A2(net821),
    .B1(_3087_),
    .X(_3088_));
 sky130_fd_sc_hd__o21a_1 _5956_ (.A1(net1843),
    .A2(net1194),
    .B1(_3088_),
    .X(_3089_));
 sky130_fd_sc_hd__mux2_1 _5957_ (.A0(_3089_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][70] ),
    .S(net980),
    .X(_0612_));
 sky130_fd_sc_hd__and3_1 _5958_ (.A(net1368),
    .B(net1372),
    .C(m3_wbd_adr_i[20]),
    .X(_3090_));
 sky130_fd_sc_hd__a221o_1 _5959_ (.A1(net1253),
    .A2(m2_wbd_adr_i[20]),
    .B1(m1_wbd_adr_i[20]),
    .B2(net821),
    .C1(net1202),
    .X(_3091_));
 sky130_fd_sc_hd__o22a_2 _5960_ (.A1(net2015),
    .A2(net1194),
    .B1(_3090_),
    .B2(_3091_),
    .X(_3092_));
 sky130_fd_sc_hd__mux2_1 _5961_ (.A0(_3092_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][71] ),
    .S(net982),
    .X(_0613_));
 sky130_fd_sc_hd__and3_1 _5962_ (.A(net1369),
    .B(net1373),
    .C(m3_wbd_adr_i[21]),
    .X(_3093_));
 sky130_fd_sc_hd__a221o_1 _5963_ (.A1(net1253),
    .A2(m2_wbd_adr_i[21]),
    .B1(net2000),
    .B2(net822),
    .C1(net1202),
    .X(_3094_));
 sky130_fd_sc_hd__o22a_1 _5964_ (.A1(net1894),
    .A2(net1195),
    .B1(_3093_),
    .B2(net2001),
    .X(_3095_));
 sky130_fd_sc_hd__mux2_1 _5965_ (.A0(_3095_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][72] ),
    .S(net981),
    .X(_0614_));
 sky130_fd_sc_hd__and3_1 _5966_ (.A(net1368),
    .B(net1372),
    .C(m3_wbd_adr_i[22]),
    .X(_3096_));
 sky130_fd_sc_hd__a221o_1 _5967_ (.A1(net1254),
    .A2(m2_wbd_adr_i[22]),
    .B1(m1_wbd_adr_i[22]),
    .B2(net822),
    .C1(net1203),
    .X(_3097_));
 sky130_fd_sc_hd__o22a_1 _5968_ (.A1(net2034),
    .A2(net1196),
    .B1(_3096_),
    .B2(_3097_),
    .X(_3098_));
 sky130_fd_sc_hd__mux2_1 _5969_ (.A0(_3098_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][73] ),
    .S(net982),
    .X(_0615_));
 sky130_fd_sc_hd__and3_1 _5970_ (.A(net1368),
    .B(net1372),
    .C(m3_wbd_adr_i[23]),
    .X(_3099_));
 sky130_fd_sc_hd__a221o_1 _5971_ (.A1(net1253),
    .A2(m2_wbd_adr_i[23]),
    .B1(net1991),
    .B2(net821),
    .C1(net1202),
    .X(_3100_));
 sky130_fd_sc_hd__o22a_1 _5972_ (.A1(net1842),
    .A2(net1194),
    .B1(_3099_),
    .B2(net1992),
    .X(_3101_));
 sky130_fd_sc_hd__mux2_1 _5973_ (.A0(_3101_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][74] ),
    .S(net979),
    .X(_0616_));
 sky130_fd_sc_hd__and3_1 _5974_ (.A(net1368),
    .B(net1372),
    .C(m3_wbd_adr_i[24]),
    .X(_3102_));
 sky130_fd_sc_hd__a221o_1 _5975_ (.A1(net1253),
    .A2(m2_wbd_adr_i[24]),
    .B1(m1_wbd_adr_i[24]),
    .B2(net822),
    .C1(net1202),
    .X(_3103_));
 sky130_fd_sc_hd__o22a_1 _5976_ (.A1(net1990),
    .A2(net1195),
    .B1(_3102_),
    .B2(_3103_),
    .X(_3104_));
 sky130_fd_sc_hd__mux2_1 _5977_ (.A0(_3104_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][75] ),
    .S(net979),
    .X(_0617_));
 sky130_fd_sc_hd__and3_1 _5978_ (.A(net1369),
    .B(net1373),
    .C(m3_wbd_adr_i[25]),
    .X(_3105_));
 sky130_fd_sc_hd__a221o_1 _5979_ (.A1(net1254),
    .A2(m2_wbd_adr_i[25]),
    .B1(m1_wbd_adr_i[25]),
    .B2(net822),
    .C1(net1202),
    .X(_3106_));
 sky130_fd_sc_hd__o22a_1 _5980_ (.A1(net2012),
    .A2(net1196),
    .B1(_3105_),
    .B2(_3106_),
    .X(_3107_));
 sky130_fd_sc_hd__mux2_1 _5981_ (.A0(_3107_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][76] ),
    .S(net981),
    .X(_0618_));
 sky130_fd_sc_hd__and3_1 _5982_ (.A(net1370),
    .B(net1373),
    .C(m3_wbd_adr_i[26]),
    .X(_3108_));
 sky130_fd_sc_hd__a221o_1 _5983_ (.A1(net1253),
    .A2(m2_wbd_adr_i[26]),
    .B1(net2090),
    .B2(net822),
    .C1(net1202),
    .X(_3109_));
 sky130_fd_sc_hd__o22a_1 _5984_ (.A1(net1847),
    .A2(net1195),
    .B1(_3108_),
    .B2(_3109_),
    .X(_3110_));
 sky130_fd_sc_hd__mux2_1 _5985_ (.A0(net1848),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][77] ),
    .S(net979),
    .X(_0619_));
 sky130_fd_sc_hd__and3_1 _5986_ (.A(net1368),
    .B(net1372),
    .C(m3_wbd_adr_i[27]),
    .X(_3111_));
 sky130_fd_sc_hd__a221o_1 _5987_ (.A1(net1253),
    .A2(m2_wbd_adr_i[27]),
    .B1(m1_wbd_adr_i[27]),
    .B2(net821),
    .C1(net1202),
    .X(_3112_));
 sky130_fd_sc_hd__o22a_1 _5988_ (.A1(net1981),
    .A2(net1194),
    .B1(_3111_),
    .B2(_3112_),
    .X(_3113_));
 sky130_fd_sc_hd__mux2_1 _5989_ (.A0(_3113_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][78] ),
    .S(net979),
    .X(_0620_));
 sky130_fd_sc_hd__a221o_2 _5990_ (.A1(net1258),
    .A2(m2_wbd_adr_i[28]),
    .B1(net1209),
    .B2(m3_wbd_adr_i[28]),
    .C1(net1204),
    .X(_3114_));
 sky130_fd_sc_hd__a21oi_2 _5991_ (.A1(m1_wbd_adr_i[28]),
    .A2(net821),
    .B1(_3114_),
    .Y(_3115_));
 sky130_fd_sc_hd__a21oi_2 _5992_ (.A1(_1683_),
    .A2(net1203),
    .B1(_3115_),
    .Y(_3116_));
 sky130_fd_sc_hd__mux2_1 _5993_ (.A0(net1901),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][79] ),
    .S(net981),
    .X(_0621_));
 sky130_fd_sc_hd__and3_2 _5994_ (.A(net1370),
    .B(net1374),
    .C(m3_wbd_adr_i[29]),
    .X(_3117_));
 sky130_fd_sc_hd__a221o_1 _5995_ (.A1(net1253),
    .A2(m2_wbd_adr_i[29]),
    .B1(m1_wbd_adr_i[29]),
    .B2(net821),
    .C1(net1202),
    .X(_3118_));
 sky130_fd_sc_hd__o22a_1 _5996_ (.A1(net1994),
    .A2(net1194),
    .B1(_3117_),
    .B2(_3118_),
    .X(_3119_));
 sky130_fd_sc_hd__mux2_1 _5997_ (.A0(_3119_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][80] ),
    .S(net979),
    .X(_0622_));
 sky130_fd_sc_hd__and3_2 _5998_ (.A(net1370),
    .B(net1374),
    .C(m3_wbd_adr_i[30]),
    .X(_3120_));
 sky130_fd_sc_hd__a221o_1 _5999_ (.A1(net1253),
    .A2(m2_wbd_adr_i[30]),
    .B1(net2086),
    .B2(net821),
    .C1(net1202),
    .X(_3121_));
 sky130_fd_sc_hd__o22a_1 _6000_ (.A1(net1866),
    .A2(net1194),
    .B1(_3120_),
    .B2(_3121_),
    .X(_3122_));
 sky130_fd_sc_hd__mux2_1 _6001_ (.A0(_3122_),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][81] ),
    .S(net979),
    .X(_0623_));
 sky130_fd_sc_hd__a221o_2 _6002_ (.A1(net1258),
    .A2(m2_wbd_adr_i[31]),
    .B1(net1206),
    .B2(m3_wbd_adr_i[31]),
    .C1(net1204),
    .X(_3123_));
 sky130_fd_sc_hd__a21o_1 _6003_ (.A1(m1_wbd_adr_i[31]),
    .A2(net821),
    .B1(_3123_),
    .X(_3124_));
 sky130_fd_sc_hd__o21a_1 _6004_ (.A1(net1852),
    .A2(net1194),
    .B1(_3124_),
    .X(_3125_));
 sky130_fd_sc_hd__mux2_1 _6005_ (.A0(net1853),
    .A1(\u_s0.u_sync_wbb.u_cmd_if.mem[0][82] ),
    .S(net980),
    .X(_0624_));
 sky130_fd_sc_hd__xor2_1 _6006_ (.A(net1382),
    .B(\u_s2.u_sync_wbb.m_resp_rd_en ),
    .X(_0625_));
 sky130_fd_sc_hd__a21oi_1 _6007_ (.A1(net1384),
    .A2(\u_s2.u_sync_wbb.m_resp_rd_en ),
    .B1(\u_s2.u_sync_wbb.u_resp_if.rd_ptr[1] ),
    .Y(_3126_));
 sky130_fd_sc_hd__and3_1 _6008_ (.A(net1379),
    .B(net1384),
    .C(\u_s2.u_sync_wbb.m_resp_rd_en ),
    .X(_3127_));
 sky130_fd_sc_hd__nor2_1 _6009_ (.A(_3126_),
    .B(_3127_),
    .Y(_0626_));
 sky130_fd_sc_hd__xor2_1 _6010_ (.A(\u_s2.u_sync_wbb.u_resp_if.rd_ptr[2] ),
    .B(_3127_),
    .X(_0627_));
 sky130_fd_sc_hd__or3_4 _6011_ (.A(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[0] ),
    .B(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .C(_2423_),
    .X(_3128_));
 sky130_fd_sc_hd__mux2_1 _6012_ (.A0(net1984),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][0] ),
    .S(net541),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _6013_ (.A0(net1902),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][1] ),
    .S(net543),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _6014_ (.A0(net2060),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][2] ),
    .S(net543),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _6015_ (.A0(net1903),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][3] ),
    .S(net543),
    .X(_0631_));
 sky130_fd_sc_hd__mux2_1 _6016_ (.A0(net2063),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][4] ),
    .S(net543),
    .X(_0632_));
 sky130_fd_sc_hd__mux2_1 _6017_ (.A0(net2065),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][5] ),
    .S(net544),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_1 _6018_ (.A0(net1880),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][6] ),
    .S(net544),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_1 _6019_ (.A0(net1886),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][7] ),
    .S(net544),
    .X(_0635_));
 sky130_fd_sc_hd__mux2_1 _6020_ (.A0(net1904),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][8] ),
    .S(net543),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _6021_ (.A0(net1892),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][9] ),
    .S(net543),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_1 _6022_ (.A0(net1898),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][10] ),
    .S(net543),
    .X(_0638_));
 sky130_fd_sc_hd__mux2_1 _6023_ (.A0(net1996),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][11] ),
    .S(net542),
    .X(_0639_));
 sky130_fd_sc_hd__mux2_1 _6024_ (.A0(net1980),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][12] ),
    .S(net541),
    .X(_0640_));
 sky130_fd_sc_hd__mux2_1 _6025_ (.A0(net1897),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][13] ),
    .S(net543),
    .X(_0641_));
 sky130_fd_sc_hd__mux2_1 _6026_ (.A0(net1841),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][14] ),
    .S(net541),
    .X(_0642_));
 sky130_fd_sc_hd__mux2_1 _6027_ (.A0(net1881),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][15] ),
    .S(net544),
    .X(_0643_));
 sky130_fd_sc_hd__mux2_1 _6028_ (.A0(net1851),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][16] ),
    .S(net541),
    .X(_0644_));
 sky130_fd_sc_hd__mux2_1 _6029_ (.A0(net1879),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][17] ),
    .S(net544),
    .X(_0645_));
 sky130_fd_sc_hd__mux2_1 _6030_ (.A0(net1889),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][18] ),
    .S(net544),
    .X(_0646_));
 sky130_fd_sc_hd__mux2_1 _6031_ (.A0(net1993),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][19] ),
    .S(net541),
    .X(_0647_));
 sky130_fd_sc_hd__mux2_1 _6032_ (.A0(net1835),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][20] ),
    .S(net541),
    .X(_0648_));
 sky130_fd_sc_hd__mux2_1 _6033_ (.A0(net1912),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][21] ),
    .S(net544),
    .X(_0649_));
 sky130_fd_sc_hd__mux2_1 _6034_ (.A0(net1844),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][22] ),
    .S(net541),
    .X(_0650_));
 sky130_fd_sc_hd__mux2_1 _6035_ (.A0(net1989),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][23] ),
    .S(net542),
    .X(_0651_));
 sky130_fd_sc_hd__mux2_1 _6036_ (.A0(net1893),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][24] ),
    .S(net543),
    .X(_0652_));
 sky130_fd_sc_hd__mux2_1 _6037_ (.A0(net2002),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][25] ),
    .S(net542),
    .X(_0653_));
 sky130_fd_sc_hd__mux2_1 _6038_ (.A0(net1988),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][26] ),
    .S(net541),
    .X(_0654_));
 sky130_fd_sc_hd__mux2_1 _6039_ (.A0(net1836),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][27] ),
    .S(net542),
    .X(_0655_));
 sky130_fd_sc_hd__mux2_1 _6040_ (.A0(net1979),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][28] ),
    .S(net542),
    .X(_0656_));
 sky130_fd_sc_hd__mux2_1 _6041_ (.A0(net1845),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][29] ),
    .S(net541),
    .X(_0657_));
 sky130_fd_sc_hd__mux2_1 _6042_ (.A0(net1838),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][30] ),
    .S(net541),
    .X(_0658_));
 sky130_fd_sc_hd__mux2_1 _6043_ (.A0(net1899),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[0][31] ),
    .S(net543),
    .X(_0659_));
 sky130_fd_sc_hd__or3b_1 _6044_ (.A(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .B(_2423_),
    .C_N(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[0] ),
    .X(_3129_));
 sky130_fd_sc_hd__mux2_1 _6045_ (.A0(net1984),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][0] ),
    .S(net537),
    .X(_0660_));
 sky130_fd_sc_hd__mux2_1 _6046_ (.A0(net1902),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][1] ),
    .S(net538),
    .X(_0661_));
 sky130_fd_sc_hd__mux2_1 _6047_ (.A0(net1882),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][2] ),
    .S(net539),
    .X(_0662_));
 sky130_fd_sc_hd__mux2_1 _6048_ (.A0(net1903),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][3] ),
    .S(net538),
    .X(_0663_));
 sky130_fd_sc_hd__mux2_1 _6049_ (.A0(net2063),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][4] ),
    .S(net539),
    .X(_0664_));
 sky130_fd_sc_hd__mux2_1 _6050_ (.A0(net2065),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][5] ),
    .S(net539),
    .X(_0665_));
 sky130_fd_sc_hd__mux2_1 _6051_ (.A0(net1880),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][6] ),
    .S(net539),
    .X(_0666_));
 sky130_fd_sc_hd__mux2_1 _6052_ (.A0(net1886),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][7] ),
    .S(net539),
    .X(_0667_));
 sky130_fd_sc_hd__mux2_1 _6053_ (.A0(net1904),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][8] ),
    .S(net538),
    .X(_0668_));
 sky130_fd_sc_hd__mux2_1 _6054_ (.A0(net1892),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][9] ),
    .S(net539),
    .X(_0669_));
 sky130_fd_sc_hd__mux2_1 _6055_ (.A0(net1898),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][10] ),
    .S(net538),
    .X(_0670_));
 sky130_fd_sc_hd__mux2_1 _6056_ (.A0(net1996),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][11] ),
    .S(net540),
    .X(_0671_));
 sky130_fd_sc_hd__mux2_1 _6057_ (.A0(net1834),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][12] ),
    .S(net540),
    .X(_0672_));
 sky130_fd_sc_hd__mux2_1 _6058_ (.A0(net2003),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][13] ),
    .S(net540),
    .X(_0673_));
 sky130_fd_sc_hd__mux2_1 _6059_ (.A0(net1841),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][14] ),
    .S(net537),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_1 _6060_ (.A0(net1881),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][15] ),
    .S(net538),
    .X(_0675_));
 sky130_fd_sc_hd__mux2_1 _6061_ (.A0(net1851),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][16] ),
    .S(net537),
    .X(_0676_));
 sky130_fd_sc_hd__mux2_1 _6062_ (.A0(net1879),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][17] ),
    .S(net539),
    .X(_0677_));
 sky130_fd_sc_hd__mux2_1 _6063_ (.A0(net1889),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][18] ),
    .S(net539),
    .X(_0678_));
 sky130_fd_sc_hd__mux2_1 _6064_ (.A0(net1993),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][19] ),
    .S(net538),
    .X(_0679_));
 sky130_fd_sc_hd__mux2_1 _6065_ (.A0(net1835),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][20] ),
    .S(net537),
    .X(_0680_));
 sky130_fd_sc_hd__mux2_1 _6066_ (.A0(net1912),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][21] ),
    .S(net539),
    .X(_0681_));
 sky130_fd_sc_hd__mux2_1 _6067_ (.A0(net1844),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][22] ),
    .S(net537),
    .X(_0682_));
 sky130_fd_sc_hd__mux2_1 _6068_ (.A0(net1989),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][23] ),
    .S(net537),
    .X(_0683_));
 sky130_fd_sc_hd__mux2_1 _6069_ (.A0(net1893),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][24] ),
    .S(net538),
    .X(_0684_));
 sky130_fd_sc_hd__mux2_1 _6070_ (.A0(net1907),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][25] ),
    .S(net538),
    .X(_0685_));
 sky130_fd_sc_hd__mux2_1 _6071_ (.A0(net1891),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][26] ),
    .S(net538),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_1 _6072_ (.A0(net1836),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][27] ),
    .S(net537),
    .X(_0687_));
 sky130_fd_sc_hd__mux2_1 _6073_ (.A0(net1979),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][28] ),
    .S(net537),
    .X(_0688_));
 sky130_fd_sc_hd__mux2_1 _6074_ (.A0(net1845),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][29] ),
    .S(net537),
    .X(_0689_));
 sky130_fd_sc_hd__mux2_1 _6075_ (.A0(net1838),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][30] ),
    .S(net537),
    .X(_0690_));
 sky130_fd_sc_hd__mux2_1 _6076_ (.A0(net1899),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[1][31] ),
    .S(net538),
    .X(_0691_));
 sky130_fd_sc_hd__or3b_1 _6077_ (.A(_2423_),
    .B(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[0] ),
    .C_N(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .X(_3130_));
 sky130_fd_sc_hd__mux2_1 _6078_ (.A0(net1984),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][0] ),
    .S(net533),
    .X(_0692_));
 sky130_fd_sc_hd__mux2_1 _6079_ (.A0(net1902),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][1] ),
    .S(net534),
    .X(_0693_));
 sky130_fd_sc_hd__mux2_1 _6080_ (.A0(net1882),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][2] ),
    .S(net535),
    .X(_0694_));
 sky130_fd_sc_hd__mux2_1 _6081_ (.A0(net1903),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][3] ),
    .S(net534),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_1 _6082_ (.A0(net1890),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][4] ),
    .S(net535),
    .X(_0696_));
 sky130_fd_sc_hd__mux2_1 _6083_ (.A0(net2065),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][5] ),
    .S(net535),
    .X(_0697_));
 sky130_fd_sc_hd__mux2_1 _6084_ (.A0(net1880),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][6] ),
    .S(net535),
    .X(_0698_));
 sky130_fd_sc_hd__mux2_1 _6085_ (.A0(net1886),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][7] ),
    .S(net535),
    .X(_0699_));
 sky130_fd_sc_hd__mux2_1 _6086_ (.A0(net1904),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][8] ),
    .S(net534),
    .X(_0700_));
 sky130_fd_sc_hd__mux2_1 _6087_ (.A0(net1892),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][9] ),
    .S(net535),
    .X(_0701_));
 sky130_fd_sc_hd__mux2_1 _6088_ (.A0(net1898),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][10] ),
    .S(net534),
    .X(_0702_));
 sky130_fd_sc_hd__mux2_1 _6089_ (.A0(net1996),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][11] ),
    .S(net536),
    .X(_0703_));
 sky130_fd_sc_hd__mux2_1 _6090_ (.A0(net1834),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][12] ),
    .S(net536),
    .X(_0704_));
 sky130_fd_sc_hd__mux2_1 _6091_ (.A0(net2003),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][13] ),
    .S(net536),
    .X(_0705_));
 sky130_fd_sc_hd__mux2_1 _6092_ (.A0(net1987),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][14] ),
    .S(net533),
    .X(_0706_));
 sky130_fd_sc_hd__mux2_1 _6093_ (.A0(net1881),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][15] ),
    .S(net534),
    .X(_0707_));
 sky130_fd_sc_hd__mux2_1 _6094_ (.A0(net1851),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][16] ),
    .S(net533),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_1 _6095_ (.A0(net1879),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][17] ),
    .S(net534),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_1 _6096_ (.A0(net1889),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][18] ),
    .S(net535),
    .X(_0710_));
 sky130_fd_sc_hd__mux2_1 _6097_ (.A0(net1993),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][19] ),
    .S(net534),
    .X(_0711_));
 sky130_fd_sc_hd__mux2_1 _6098_ (.A0(net1835),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][20] ),
    .S(net533),
    .X(_0712_));
 sky130_fd_sc_hd__mux2_1 _6099_ (.A0(net1912),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][21] ),
    .S(net535),
    .X(_0713_));
 sky130_fd_sc_hd__mux2_1 _6100_ (.A0(net1844),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][22] ),
    .S(net533),
    .X(_0714_));
 sky130_fd_sc_hd__mux2_1 _6101_ (.A0(net1846),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][23] ),
    .S(net533),
    .X(_0715_));
 sky130_fd_sc_hd__mux2_1 _6102_ (.A0(net1893),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][24] ),
    .S(net534),
    .X(_0716_));
 sky130_fd_sc_hd__mux2_1 _6103_ (.A0(net1907),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][25] ),
    .S(net534),
    .X(_0717_));
 sky130_fd_sc_hd__mux2_1 _6104_ (.A0(net1891),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][26] ),
    .S(net534),
    .X(_0718_));
 sky130_fd_sc_hd__mux2_1 _6105_ (.A0(net1982),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][27] ),
    .S(net536),
    .X(_0719_));
 sky130_fd_sc_hd__mux2_1 _6106_ (.A0(net1837),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][28] ),
    .S(net533),
    .X(_0720_));
 sky130_fd_sc_hd__mux2_1 _6107_ (.A0(net1845),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][29] ),
    .S(net533),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_1 _6108_ (.A0(net1838),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][30] ),
    .S(net533),
    .X(_0722_));
 sky130_fd_sc_hd__mux2_1 _6109_ (.A0(net1899),
    .A1(\u_s0.u_sync_wbb.u_resp_if.mem[2][31] ),
    .S(net533),
    .X(_0723_));
 sky130_fd_sc_hd__and3_2 _6110_ (.A(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[0] ),
    .B(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .C(_2424_),
    .X(_3131_));
 sky130_fd_sc_hd__mux2_1 _6111_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][0] ),
    .A1(net1984),
    .S(net495),
    .X(_0724_));
 sky130_fd_sc_hd__mux2_1 _6112_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][1] ),
    .A1(net1902),
    .S(net497),
    .X(_0725_));
 sky130_fd_sc_hd__mux2_1 _6113_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][2] ),
    .A1(net1882),
    .S(net496),
    .X(_0726_));
 sky130_fd_sc_hd__mux2_1 _6114_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][3] ),
    .A1(net1903),
    .S(net497),
    .X(_0727_));
 sky130_fd_sc_hd__mux2_1 _6115_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][4] ),
    .A1(net2063),
    .S(net496),
    .X(_0728_));
 sky130_fd_sc_hd__mux2_1 _6116_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][5] ),
    .A1(net2065),
    .S(net496),
    .X(_0729_));
 sky130_fd_sc_hd__mux2_1 _6117_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][6] ),
    .A1(net1880),
    .S(net496),
    .X(_0730_));
 sky130_fd_sc_hd__mux2_1 _6118_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][7] ),
    .A1(net1886),
    .S(net496),
    .X(_0731_));
 sky130_fd_sc_hd__mux2_1 _6119_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][8] ),
    .A1(net1904),
    .S(net497),
    .X(_0732_));
 sky130_fd_sc_hd__mux2_1 _6120_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][9] ),
    .A1(net1892),
    .S(net496),
    .X(_0733_));
 sky130_fd_sc_hd__mux2_1 _6121_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][10] ),
    .A1(net1999),
    .S(net497),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_1 _6122_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][11] ),
    .A1(net1996),
    .S(net495),
    .X(_0735_));
 sky130_fd_sc_hd__mux2_1 _6123_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][12] ),
    .A1(net1980),
    .S(net494),
    .X(_0736_));
 sky130_fd_sc_hd__mux2_1 _6124_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][13] ),
    .A1(net2003),
    .S(net495),
    .X(_0737_));
 sky130_fd_sc_hd__mux2_1 _6125_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][14] ),
    .A1(net1987),
    .S(net494),
    .X(_0738_));
 sky130_fd_sc_hd__mux2_1 _6126_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][15] ),
    .A1(net1881),
    .S(net496),
    .X(_0739_));
 sky130_fd_sc_hd__mux2_1 _6127_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][16] ),
    .A1(net1851),
    .S(net494),
    .X(_0740_));
 sky130_fd_sc_hd__mux2_1 _6128_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][17] ),
    .A1(net1879),
    .S(net496),
    .X(_0741_));
 sky130_fd_sc_hd__mux2_1 _6129_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][18] ),
    .A1(net1889),
    .S(net497),
    .X(_0742_));
 sky130_fd_sc_hd__mux2_1 _6130_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][19] ),
    .A1(net1993),
    .S(net494),
    .X(_0743_));
 sky130_fd_sc_hd__mux2_1 _6131_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][20] ),
    .A1(net1978),
    .S(net494),
    .X(_0744_));
 sky130_fd_sc_hd__mux2_1 _6132_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][21] ),
    .A1(net1912),
    .S(net496),
    .X(_0745_));
 sky130_fd_sc_hd__mux2_1 _6133_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][22] ),
    .A1(net1844),
    .S(net494),
    .X(_0746_));
 sky130_fd_sc_hd__mux2_1 _6134_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][23] ),
    .A1(net1846),
    .S(net495),
    .X(_0747_));
 sky130_fd_sc_hd__mux2_1 _6135_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][24] ),
    .A1(net1893),
    .S(net497),
    .X(_0748_));
 sky130_fd_sc_hd__mux2_1 _6136_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][25] ),
    .A1(net1907),
    .S(net497),
    .X(_0749_));
 sky130_fd_sc_hd__mux2_1 _6137_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][26] ),
    .A1(net1891),
    .S(net494),
    .X(_0750_));
 sky130_fd_sc_hd__mux2_1 _6138_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][27] ),
    .A1(net1836),
    .S(net495),
    .X(_0751_));
 sky130_fd_sc_hd__mux2_1 _6139_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][28] ),
    .A1(net1837),
    .S(net494),
    .X(_0752_));
 sky130_fd_sc_hd__mux2_1 _6140_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][29] ),
    .A1(net1845),
    .S(net494),
    .X(_0753_));
 sky130_fd_sc_hd__mux2_1 _6141_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][30] ),
    .A1(net1838),
    .S(net494),
    .X(_0754_));
 sky130_fd_sc_hd__mux2_1 _6142_ (.A0(\u_s0.u_sync_wbb.u_resp_if.mem[3][31] ),
    .A1(net1899),
    .S(net497),
    .X(_0755_));
 sky130_fd_sc_hd__mux2_1 _6143_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][1] ),
    .A1(net791),
    .S(net995),
    .X(_0756_));
 sky130_fd_sc_hd__mux2_1 _6144_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][2] ),
    .A1(net794),
    .S(net993),
    .X(_0757_));
 sky130_fd_sc_hd__mux2_1 _6145_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][3] ),
    .A1(net792),
    .S(net995),
    .X(_0758_));
 sky130_fd_sc_hd__mux2_1 _6146_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][4] ),
    .A1(net795),
    .S(net995),
    .X(_0759_));
 sky130_fd_sc_hd__mux2_1 _6147_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][5] ),
    .A1(net786),
    .S(net989),
    .X(_0760_));
 sky130_fd_sc_hd__mux2_1 _6148_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][6] ),
    .A1(net788),
    .S(net993),
    .X(_0761_));
 sky130_fd_sc_hd__mux2_1 _6149_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][7] ),
    .A1(net789),
    .S(net990),
    .X(_0762_));
 sky130_fd_sc_hd__mux2_1 _6150_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][8] ),
    .A1(net790),
    .S(net990),
    .X(_0763_));
 sky130_fd_sc_hd__mux2_1 _6151_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][9] ),
    .A1(net785),
    .S(net994),
    .X(_0764_));
 sky130_fd_sc_hd__and2_1 _6152_ (.A(m1_wbd_sel_i[0]),
    .B(net1175),
    .X(_3132_));
 sky130_fd_sc_hd__a221o_1 _6153_ (.A1(net1238),
    .A2(net2082),
    .B1(net1179),
    .B2(m3_wbd_sel_i[0]),
    .C1(net1172),
    .X(_3133_));
 sky130_fd_sc_hd__o22a_2 _6154_ (.A1(net1565),
    .A2(net1171),
    .B1(_3132_),
    .B2(_3133_),
    .X(_3134_));
 sky130_fd_sc_hd__mux2_1 _6155_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][14] ),
    .A1(net677),
    .S(net995),
    .X(_0765_));
 sky130_fd_sc_hd__and3_1 _6156_ (.A(net1410),
    .B(net1408),
    .C(m3_wbd_sel_i[1]),
    .X(_3135_));
 sky130_fd_sc_hd__a221o_1 _6157_ (.A1(net1233),
    .A2(m2_wbd_sel_i[1]),
    .B1(m1_wbd_sel_i[1]),
    .B2(net1174),
    .C1(net1172),
    .X(_3136_));
 sky130_fd_sc_hd__o22a_4 _6158_ (.A1(net1915),
    .A2(net1167),
    .B1(_3135_),
    .B2(_3136_),
    .X(_3137_));
 sky130_fd_sc_hd__mux2_1 _6159_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][15] ),
    .A1(net675),
    .S(net995),
    .X(_0766_));
 sky130_fd_sc_hd__and3_1 _6160_ (.A(net1410),
    .B(net1408),
    .C(m3_wbd_sel_i[2]),
    .X(_3138_));
 sky130_fd_sc_hd__a221o_1 _6161_ (.A1(net1232),
    .A2(m2_wbd_sel_i[2]),
    .B1(m1_wbd_sel_i[2]),
    .B2(net1174),
    .C1(net1173),
    .X(_3139_));
 sky130_fd_sc_hd__o22a_1 _6162_ (.A1(net1974),
    .A2(net1166),
    .B1(_3138_),
    .B2(_3139_),
    .X(_3140_));
 sky130_fd_sc_hd__mux2_1 _6163_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][16] ),
    .A1(net673),
    .S(net994),
    .X(_0767_));
 sky130_fd_sc_hd__and3_1 _6164_ (.A(net1410),
    .B(net1407),
    .C(m3_wbd_sel_i[3]),
    .X(_3141_));
 sky130_fd_sc_hd__a221o_1 _6165_ (.A1(net1232),
    .A2(net2087),
    .B1(net2059),
    .B2(net1174),
    .C1(net1172),
    .X(_3142_));
 sky130_fd_sc_hd__o22a_4 _6166_ (.A1(net1970),
    .A2(net1166),
    .B1(_3141_),
    .B2(_3142_),
    .X(_3143_));
 sky130_fd_sc_hd__mux2_1 _6167_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][17] ),
    .A1(net672),
    .S(net990),
    .X(_0768_));
 sky130_fd_sc_hd__a21o_1 _6168_ (.A1(net1225),
    .A2(net1562),
    .B1(net1233),
    .X(_3144_));
 sky130_fd_sc_hd__o221a_4 _6169_ (.A1(net1225),
    .A2(net2050),
    .B1(net1593),
    .B2(net1167),
    .C1(_3144_),
    .X(_3145_));
 sky130_fd_sc_hd__mux2_1 _6170_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][18] ),
    .A1(net671),
    .S(net991),
    .X(_0769_));
 sky130_fd_sc_hd__a21o_1 _6171_ (.A1(net1225),
    .A2(net1551),
    .B1(net1233),
    .X(_3146_));
 sky130_fd_sc_hd__o221a_2 _6172_ (.A1(net1225),
    .A2(net2078),
    .B1(net1582),
    .B2(net1167),
    .C1(_3146_),
    .X(_3147_));
 sky130_fd_sc_hd__mux2_1 _6173_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][19] ),
    .A1(net670),
    .S(net990),
    .X(_0770_));
 sky130_fd_sc_hd__or2_1 _6174_ (.A(net1574),
    .B(net1170),
    .X(_3148_));
 sky130_fd_sc_hd__a21o_1 _6175_ (.A1(net1227),
    .A2(net1543),
    .B1(net1237),
    .X(_3149_));
 sky130_fd_sc_hd__o211a_4 _6176_ (.A1(net1227),
    .A2(net1855),
    .B1(_3148_),
    .C1(_3149_),
    .X(_3150_));
 sky130_fd_sc_hd__mux2_1 _6177_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][20] ),
    .A1(net669),
    .S(net995),
    .X(_0771_));
 sky130_fd_sc_hd__or2_1 _6178_ (.A(m0_wbd_dat_i[3]),
    .B(net1166),
    .X(_3151_));
 sky130_fd_sc_hd__a21o_1 _6179_ (.A1(net1224),
    .A2(m1_wbd_dat_i[3]),
    .B1(net1232),
    .X(_3152_));
 sky130_fd_sc_hd__o211a_1 _6180_ (.A1(net1224),
    .A2(net2088),
    .B1(_3151_),
    .C1(_3152_),
    .X(_3153_));
 sky130_fd_sc_hd__mux2_1 _6181_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][21] ),
    .A1(net667),
    .S(net994),
    .X(_0772_));
 sky130_fd_sc_hd__a21o_1 _6182_ (.A1(net1226),
    .A2(net1540),
    .B1(net1237),
    .X(_3154_));
 sky130_fd_sc_hd__o221a_4 _6183_ (.A1(net1226),
    .A2(net1518),
    .B1(net1571),
    .B2(net1170),
    .C1(_3154_),
    .X(_3155_));
 sky130_fd_sc_hd__mux2_1 _6184_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][22] ),
    .A1(net666),
    .S(net994),
    .X(_0773_));
 sky130_fd_sc_hd__a21o_1 _6185_ (.A1(net1228),
    .A2(net1539),
    .B1(net1236),
    .X(_3156_));
 sky130_fd_sc_hd__o221a_1 _6186_ (.A1(net1228),
    .A2(net1517),
    .B1(net1570),
    .B2(net1169),
    .C1(_3156_),
    .X(_3157_));
 sky130_fd_sc_hd__mux2_1 _6187_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][23] ),
    .A1(net665),
    .S(net990),
    .X(_0774_));
 sky130_fd_sc_hd__or2_1 _6188_ (.A(net1569),
    .B(net1168),
    .X(_3158_));
 sky130_fd_sc_hd__a21o_1 _6189_ (.A1(net1235),
    .A2(net1516),
    .B1(net1230),
    .X(_3159_));
 sky130_fd_sc_hd__o211a_1 _6190_ (.A1(net1235),
    .A2(net1538),
    .B1(_3158_),
    .C1(_3159_),
    .X(_3160_));
 sky130_fd_sc_hd__mux2_1 _6191_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][24] ),
    .A1(net664),
    .S(net991),
    .X(_0775_));
 sky130_fd_sc_hd__a21o_1 _6192_ (.A1(net1230),
    .A2(net1537),
    .B1(net1235),
    .X(_3161_));
 sky130_fd_sc_hd__o221a_4 _6193_ (.A1(net1230),
    .A2(net1515),
    .B1(net1568),
    .B2(net1168),
    .C1(_3161_),
    .X(_3162_));
 sky130_fd_sc_hd__mux2_1 _6194_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][25] ),
    .A1(net663),
    .S(net995),
    .X(_0776_));
 sky130_fd_sc_hd__a21o_1 _6195_ (.A1(net1229),
    .A2(net1536),
    .B1(net1234),
    .X(_3163_));
 sky130_fd_sc_hd__o221a_4 _6196_ (.A1(net1229),
    .A2(net1514),
    .B1(net1567),
    .B2(net1168),
    .C1(_3163_),
    .X(_3164_));
 sky130_fd_sc_hd__mux2_1 _6197_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][26] ),
    .A1(_3164_),
    .S(net992),
    .X(_0777_));
 sky130_fd_sc_hd__or2_1 _6198_ (.A(net1566),
    .B(net1168),
    .X(_3165_));
 sky130_fd_sc_hd__a21o_1 _6199_ (.A1(net1229),
    .A2(net1535),
    .B1(net1234),
    .X(_3166_));
 sky130_fd_sc_hd__o211a_1 _6200_ (.A1(net1229),
    .A2(net1513),
    .B1(_3165_),
    .C1(_3166_),
    .X(_3167_));
 sky130_fd_sc_hd__mux2_1 _6201_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][27] ),
    .A1(net662),
    .S(net994),
    .X(_0778_));
 sky130_fd_sc_hd__or2_1 _6202_ (.A(net1592),
    .B(net1169),
    .X(_3168_));
 sky130_fd_sc_hd__a21o_1 _6203_ (.A1(net1236),
    .A2(net1534),
    .B1(net1228),
    .X(_3169_));
 sky130_fd_sc_hd__o211a_2 _6204_ (.A1(net1236),
    .A2(net1561),
    .B1(_3168_),
    .C1(_3169_),
    .X(_3170_));
 sky130_fd_sc_hd__mux2_1 _6205_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][28] ),
    .A1(net661),
    .S(net993),
    .X(_0779_));
 sky130_fd_sc_hd__a21o_1 _6206_ (.A1(net1228),
    .A2(net1560),
    .B1(net1236),
    .X(_3171_));
 sky130_fd_sc_hd__o221a_1 _6207_ (.A1(net1228),
    .A2(net1533),
    .B1(net1591),
    .B2(net1169),
    .C1(_3171_),
    .X(_3172_));
 sky130_fd_sc_hd__mux2_1 _6208_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][29] ),
    .A1(net660),
    .S(net989),
    .X(_0780_));
 sky130_fd_sc_hd__a21o_1 _6209_ (.A1(net1230),
    .A2(net1559),
    .B1(net1234),
    .X(_3173_));
 sky130_fd_sc_hd__o221a_1 _6210_ (.A1(net1230),
    .A2(net1532),
    .B1(net1590),
    .B2(net1168),
    .C1(_3173_),
    .X(_3174_));
 sky130_fd_sc_hd__mux2_1 _6211_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][30] ),
    .A1(net659),
    .S(net994),
    .X(_0781_));
 sky130_fd_sc_hd__a21o_1 _6212_ (.A1(net1226),
    .A2(net1558),
    .B1(net1237),
    .X(_3175_));
 sky130_fd_sc_hd__o221a_1 _6213_ (.A1(net1226),
    .A2(net2066),
    .B1(net1589),
    .B2(net1170),
    .C1(_3175_),
    .X(_3176_));
 sky130_fd_sc_hd__mux2_1 _6214_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][31] ),
    .A1(net658),
    .S(net989),
    .X(_0782_));
 sky130_fd_sc_hd__or2_1 _6215_ (.A(net1588),
    .B(net1169),
    .X(_3177_));
 sky130_fd_sc_hd__a21o_1 _6216_ (.A1(net1228),
    .A2(net1557),
    .B1(net1236),
    .X(_3178_));
 sky130_fd_sc_hd__o211a_2 _6217_ (.A1(net1228),
    .A2(net1531),
    .B1(_3177_),
    .C1(_3178_),
    .X(_3179_));
 sky130_fd_sc_hd__mux2_1 _6218_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][32] ),
    .A1(net657),
    .S(net993),
    .X(_0783_));
 sky130_fd_sc_hd__or2_1 _6219_ (.A(net1587),
    .B(net1170),
    .X(_3180_));
 sky130_fd_sc_hd__a21o_1 _6220_ (.A1(net1227),
    .A2(net1556),
    .B1(net1237),
    .X(_3181_));
 sky130_fd_sc_hd__o211a_2 _6221_ (.A1(net1227),
    .A2(net1530),
    .B1(_3180_),
    .C1(_3181_),
    .X(_3182_));
 sky130_fd_sc_hd__mux2_1 _6222_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][33] ),
    .A1(net656),
    .S(net991),
    .X(_0784_));
 sky130_fd_sc_hd__or2_1 _6223_ (.A(net1586),
    .B(net1168),
    .X(_3183_));
 sky130_fd_sc_hd__a21o_1 _6224_ (.A1(net1234),
    .A2(net1529),
    .B1(net1229),
    .X(_3184_));
 sky130_fd_sc_hd__o211a_2 _6225_ (.A1(net1234),
    .A2(net1555),
    .B1(_3183_),
    .C1(_3184_),
    .X(_3185_));
 sky130_fd_sc_hd__mux2_1 _6226_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][34] ),
    .A1(net655),
    .S(net993),
    .X(_0785_));
 sky130_fd_sc_hd__or2_1 _6227_ (.A(net1585),
    .B(net1168),
    .X(_3186_));
 sky130_fd_sc_hd__a21o_1 _6228_ (.A1(net1234),
    .A2(net1528),
    .B1(net1229),
    .X(_3187_));
 sky130_fd_sc_hd__o211a_2 _6229_ (.A1(net1234),
    .A2(net1554),
    .B1(_3186_),
    .C1(_3187_),
    .X(_3188_));
 sky130_fd_sc_hd__mux2_1 _6230_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][35] ),
    .A1(net654),
    .S(net993),
    .X(_0786_));
 sky130_fd_sc_hd__or2_1 _6231_ (.A(net1584),
    .B(net1167),
    .X(_3189_));
 sky130_fd_sc_hd__a21o_1 _6232_ (.A1(net1225),
    .A2(net1553),
    .B1(net1233),
    .X(_3190_));
 sky130_fd_sc_hd__o211a_1 _6233_ (.A1(net1225),
    .A2(net1928),
    .B1(_3189_),
    .C1(_3190_),
    .X(_3191_));
 sky130_fd_sc_hd__mux2_1 _6234_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][36] ),
    .A1(net652),
    .S(net993),
    .X(_0787_));
 sky130_fd_sc_hd__a21o_1 _6235_ (.A1(net1229),
    .A2(net1552),
    .B1(net1234),
    .X(_3192_));
 sky130_fd_sc_hd__o221a_2 _6236_ (.A1(net1229),
    .A2(net1527),
    .B1(net1583),
    .B2(net1169),
    .C1(_3192_),
    .X(_3193_));
 sky130_fd_sc_hd__mux2_1 _6237_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][37] ),
    .A1(net651),
    .S(_2934_),
    .X(_0788_));
 sky130_fd_sc_hd__a21o_1 _6238_ (.A1(net1230),
    .A2(net1550),
    .B1(net1235),
    .X(_3194_));
 sky130_fd_sc_hd__o221a_4 _6239_ (.A1(net1230),
    .A2(net1526),
    .B1(net1581),
    .B2(net1168),
    .C1(_3194_),
    .X(_3195_));
 sky130_fd_sc_hd__mux2_1 _6240_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][38] ),
    .A1(_3195_),
    .S(net989),
    .X(_0789_));
 sky130_fd_sc_hd__a21o_1 _6241_ (.A1(net1226),
    .A2(net1549),
    .B1(net1237),
    .X(_3196_));
 sky130_fd_sc_hd__o221a_1 _6242_ (.A1(net1226),
    .A2(net1525),
    .B1(net1580),
    .B2(net1170),
    .C1(_3196_),
    .X(_3197_));
 sky130_fd_sc_hd__mux2_1 _6243_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][39] ),
    .A1(net650),
    .S(net989),
    .X(_0790_));
 sky130_fd_sc_hd__or2_1 _6244_ (.A(net1579),
    .B(net1170),
    .X(_3198_));
 sky130_fd_sc_hd__a21o_1 _6245_ (.A1(net1226),
    .A2(net1548),
    .B1(net1237),
    .X(_3199_));
 sky130_fd_sc_hd__o211a_1 _6246_ (.A1(net1226),
    .A2(net2051),
    .B1(_3198_),
    .C1(_3199_),
    .X(_3200_));
 sky130_fd_sc_hd__mux2_1 _6247_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][40] ),
    .A1(net649),
    .S(net990),
    .X(_0791_));
 sky130_fd_sc_hd__a21o_1 _6248_ (.A1(net1226),
    .A2(net1547),
    .B1(net1237),
    .X(_3201_));
 sky130_fd_sc_hd__o221a_1 _6249_ (.A1(net1226),
    .A2(net1524),
    .B1(net1578),
    .B2(net1170),
    .C1(_3201_),
    .X(_3202_));
 sky130_fd_sc_hd__mux2_1 _6250_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][41] ),
    .A1(net648),
    .S(net989),
    .X(_0792_));
 sky130_fd_sc_hd__a21o_1 _6251_ (.A1(net1224),
    .A2(m1_wbd_dat_i[24]),
    .B1(net1232),
    .X(_3203_));
 sky130_fd_sc_hd__o221a_4 _6252_ (.A1(net1224),
    .A2(net1839),
    .B1(m0_wbd_dat_i[24]),
    .B2(net1166),
    .C1(_3203_),
    .X(_3204_));
 sky130_fd_sc_hd__mux2_1 _6253_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][42] ),
    .A1(net647),
    .S(net990),
    .X(_0793_));
 sky130_fd_sc_hd__a21o_1 _6254_ (.A1(net1224),
    .A2(m1_wbd_dat_i[25]),
    .B1(net1232),
    .X(_3205_));
 sky130_fd_sc_hd__o221a_1 _6255_ (.A1(net1224),
    .A2(net1934),
    .B1(m0_wbd_dat_i[25]),
    .B2(net1166),
    .C1(_3205_),
    .X(_3206_));
 sky130_fd_sc_hd__mux2_1 _6256_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][43] ),
    .A1(net645),
    .S(net990),
    .X(_0794_));
 sky130_fd_sc_hd__or2_1 _6257_ (.A(net1577),
    .B(net1168),
    .X(_3207_));
 sky130_fd_sc_hd__a21o_1 _6258_ (.A1(net1229),
    .A2(net1546),
    .B1(net1235),
    .X(_3208_));
 sky130_fd_sc_hd__o211a_4 _6259_ (.A1(net1230),
    .A2(net1523),
    .B1(_3207_),
    .C1(_3208_),
    .X(_3209_));
 sky130_fd_sc_hd__mux2_1 _6260_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][44] ),
    .A1(net644),
    .S(net995),
    .X(_0795_));
 sky130_fd_sc_hd__or2_1 _6261_ (.A(net1576),
    .B(net1168),
    .X(_3210_));
 sky130_fd_sc_hd__a21o_1 _6262_ (.A1(net1234),
    .A2(net1522),
    .B1(net1229),
    .X(_3211_));
 sky130_fd_sc_hd__o211a_1 _6263_ (.A1(net1234),
    .A2(net1545),
    .B1(_3210_),
    .C1(_3211_),
    .X(_3212_));
 sky130_fd_sc_hd__mux2_1 _6264_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][45] ),
    .A1(net643),
    .S(net993),
    .X(_0796_));
 sky130_fd_sc_hd__a21o_1 _6265_ (.A1(net1224),
    .A2(m1_wbd_dat_i[28]),
    .B1(net1232),
    .X(_3213_));
 sky130_fd_sc_hd__o221a_4 _6266_ (.A1(net1224),
    .A2(net2013),
    .B1(m0_wbd_dat_i[28]),
    .B2(net1166),
    .C1(_3213_),
    .X(_3214_));
 sky130_fd_sc_hd__mux2_1 _6267_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][46] ),
    .A1(net642),
    .S(net992),
    .X(_0797_));
 sky130_fd_sc_hd__a21o_1 _6268_ (.A1(net1228),
    .A2(net1544),
    .B1(net1236),
    .X(_3215_));
 sky130_fd_sc_hd__o221a_4 _6269_ (.A1(net1228),
    .A2(net1521),
    .B1(net1575),
    .B2(net1169),
    .C1(_3215_),
    .X(_3216_));
 sky130_fd_sc_hd__mux2_1 _6270_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][47] ),
    .A1(net2029),
    .S(net989),
    .X(_0798_));
 sky130_fd_sc_hd__or2_1 _6271_ (.A(net1573),
    .B(net1170),
    .X(_3217_));
 sky130_fd_sc_hd__a21o_1 _6272_ (.A1(net1227),
    .A2(net1542),
    .B1(net1237),
    .X(_3218_));
 sky130_fd_sc_hd__o211a_2 _6273_ (.A1(net1227),
    .A2(net1520),
    .B1(_3217_),
    .C1(_3218_),
    .X(_3219_));
 sky130_fd_sc_hd__mux2_1 _6274_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][48] ),
    .A1(net641),
    .S(net991),
    .X(_0799_));
 sky130_fd_sc_hd__a21o_1 _6275_ (.A1(net1228),
    .A2(net1541),
    .B1(net1236),
    .X(_3220_));
 sky130_fd_sc_hd__o221a_1 _6276_ (.A1(net1231),
    .A2(net1519),
    .B1(net1572),
    .B2(net1169),
    .C1(_3220_),
    .X(_3221_));
 sky130_fd_sc_hd__mux2_1 _6277_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][49] ),
    .A1(net640),
    .S(net992),
    .X(_0800_));
 sky130_fd_sc_hd__mux2_1 _6278_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][50] ),
    .A1(net726),
    .S(net993),
    .X(_0801_));
 sky130_fd_sc_hd__a221o_1 _6279_ (.A1(net1238),
    .A2(m2_wbd_adr_i[2]),
    .B1(net1178),
    .B2(m3_wbd_adr_i[2]),
    .C1(net1172),
    .X(_3222_));
 sky130_fd_sc_hd__a21o_1 _6280_ (.A1(net1883),
    .A2(net1175),
    .B1(_3222_),
    .X(_3223_));
 sky130_fd_sc_hd__o21a_4 _6281_ (.A1(net1598),
    .A2(net1171),
    .B1(net1884),
    .X(_3224_));
 sky130_fd_sc_hd__mux2_1 _6282_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][53] ),
    .A1(net585),
    .S(net991),
    .X(_0802_));
 sky130_fd_sc_hd__and3_1 _6283_ (.A(net1410),
    .B(net1408),
    .C(m3_wbd_adr_i[3]),
    .X(_3225_));
 sky130_fd_sc_hd__a221o_1 _6284_ (.A1(net1233),
    .A2(net1931),
    .B1(m1_wbd_adr_i[3]),
    .B2(net1174),
    .C1(net1172),
    .X(_3226_));
 sky130_fd_sc_hd__o22a_4 _6285_ (.A1(net1597),
    .A2(net1167),
    .B1(_3225_),
    .B2(net1932),
    .X(_3227_));
 sky130_fd_sc_hd__mux2_1 _6286_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][54] ),
    .A1(net639),
    .S(net991),
    .X(_0803_));
 sky130_fd_sc_hd__and3_1 _6287_ (.A(\u_s2.gnt[0] ),
    .B(net1408),
    .C(m3_wbd_adr_i[4]),
    .X(_3228_));
 sky130_fd_sc_hd__a221o_1 _6288_ (.A1(net1238),
    .A2(net1917),
    .B1(m1_wbd_adr_i[4]),
    .B2(net1175),
    .C1(net1172),
    .X(_3229_));
 sky130_fd_sc_hd__o22a_4 _6289_ (.A1(net1596),
    .A2(net1171),
    .B1(_3228_),
    .B2(net1918),
    .X(_3230_));
 sky130_fd_sc_hd__mux2_1 _6290_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][55] ),
    .A1(net638),
    .S(net991),
    .X(_0804_));
 sky130_fd_sc_hd__and2_1 _6291_ (.A(m1_wbd_adr_i[5]),
    .B(net1175),
    .X(_3231_));
 sky130_fd_sc_hd__a221o_1 _6292_ (.A1(net1233),
    .A2(net1887),
    .B1(net1178),
    .B2(m3_wbd_adr_i[5]),
    .C1(net1172),
    .X(_3232_));
 sky130_fd_sc_hd__o22a_4 _6293_ (.A1(net1595),
    .A2(net1167),
    .B1(_3231_),
    .B2(_3232_),
    .X(_3233_));
 sky130_fd_sc_hd__mux2_1 _6294_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][56] ),
    .A1(net637),
    .S(net990),
    .X(_0805_));
 sky130_fd_sc_hd__and3_1 _6295_ (.A(net1409),
    .B(\u_s2.gnt[1] ),
    .C(m3_wbd_adr_i[6]),
    .X(_3234_));
 sky130_fd_sc_hd__a221o_1 _6296_ (.A1(net1233),
    .A2(m2_wbd_adr_i[6]),
    .B1(m1_wbd_adr_i[6]),
    .B2(net1174),
    .C1(net1172),
    .X(_3235_));
 sky130_fd_sc_hd__o22a_4 _6297_ (.A1(net1832),
    .A2(net1167),
    .B1(_3234_),
    .B2(_3235_),
    .X(_3236_));
 sky130_fd_sc_hd__mux2_1 _6298_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][57] ),
    .A1(net636),
    .S(net990),
    .X(_0806_));
 sky130_fd_sc_hd__and2_1 _6299_ (.A(m1_wbd_adr_i[7]),
    .B(net1175),
    .X(_3237_));
 sky130_fd_sc_hd__a221o_1 _6300_ (.A1(net1238),
    .A2(m2_wbd_adr_i[7]),
    .B1(net1178),
    .B2(m3_wbd_adr_i[7]),
    .C1(net1173),
    .X(_3238_));
 sky130_fd_sc_hd__o22a_2 _6301_ (.A1(net1594),
    .A2(net1171),
    .B1(_3237_),
    .B2(_3238_),
    .X(_3239_));
 sky130_fd_sc_hd__mux2_1 _6302_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][58] ),
    .A1(net635),
    .S(net989),
    .X(_0807_));
 sky130_fd_sc_hd__and2_1 _6303_ (.A(m1_wbd_adr_i[8]),
    .B(net1174),
    .X(_3240_));
 sky130_fd_sc_hd__a221o_1 _6304_ (.A1(net1233),
    .A2(net2025),
    .B1(net1179),
    .B2(m3_wbd_adr_i[8]),
    .C1(net1172),
    .X(_3241_));
 sky130_fd_sc_hd__o22a_1 _6305_ (.A1(net1946),
    .A2(net1167),
    .B1(_3240_),
    .B2(_3241_),
    .X(_3242_));
 sky130_fd_sc_hd__mux2_1 _6306_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][59] ),
    .A1(net633),
    .S(net991),
    .X(_0808_));
 sky130_fd_sc_hd__and3_1 _6307_ (.A(net1409),
    .B(net1407),
    .C(m3_wbd_adr_i[9]),
    .X(_3243_));
 sky130_fd_sc_hd__a221o_1 _6308_ (.A1(net1232),
    .A2(net2074),
    .B1(net2032),
    .B2(net1176),
    .C1(net1173),
    .X(_3244_));
 sky130_fd_sc_hd__o22a_4 _6309_ (.A1(net1954),
    .A2(net1166),
    .B1(_3243_),
    .B2(_3244_),
    .X(_3245_));
 sky130_fd_sc_hd__mux2_1 _6310_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][60] ),
    .A1(net632),
    .S(net989),
    .X(_0809_));
 sky130_fd_sc_hd__and3_1 _6311_ (.A(net1409),
    .B(net1407),
    .C(m3_wbd_adr_i[10]),
    .X(_3246_));
 sky130_fd_sc_hd__a221o_1 _6312_ (.A1(net1232),
    .A2(m2_wbd_adr_i[10]),
    .B1(m1_wbd_adr_i[10]),
    .B2(net1176),
    .C1(net1173),
    .X(_3247_));
 sky130_fd_sc_hd__o22a_4 _6313_ (.A1(m0_wbd_adr_i[10]),
    .A2(net1166),
    .B1(_3246_),
    .B2(_3247_),
    .X(_3248_));
 sky130_fd_sc_hd__mux2_1 _6314_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[3][61] ),
    .A1(net631),
    .S(net989),
    .X(_0810_));
 sky130_fd_sc_hd__mux2_1 _6315_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[0] ),
    .A1(_2426_),
    .S(net567),
    .X(_0811_));
 sky130_fd_sc_hd__mux2_1 _6316_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[1] ),
    .A1(_1912_),
    .S(net565),
    .X(_0812_));
 sky130_fd_sc_hd__mux2_1 _6317_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[2] ),
    .A1(net1181),
    .S(net565),
    .X(_0813_));
 sky130_fd_sc_hd__mux2_1 _6318_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[3] ),
    .A1(_1910_),
    .S(net569),
    .X(_0814_));
 sky130_fd_sc_hd__mux2_1 _6319_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[4] ),
    .A1(_1909_),
    .S(net568),
    .X(_0815_));
 sky130_fd_sc_hd__mux2_1 _6320_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[5] ),
    .A1(_1908_),
    .S(net569),
    .X(_0816_));
 sky130_fd_sc_hd__mux2_1 _6321_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[6] ),
    .A1(_1907_),
    .S(net569),
    .X(_0817_));
 sky130_fd_sc_hd__mux2_1 _6322_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[7] ),
    .A1(_1906_),
    .S(net569),
    .X(_0818_));
 sky130_fd_sc_hd__mux2_1 _6323_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[8] ),
    .A1(_1905_),
    .S(net571),
    .X(_0819_));
 sky130_fd_sc_hd__mux2_1 _6324_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[9] ),
    .A1(_1904_),
    .S(net570),
    .X(_0820_));
 sky130_fd_sc_hd__mux2_1 _6325_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[14] ),
    .A1(_2427_),
    .S(net567),
    .X(_0821_));
 sky130_fd_sc_hd__mux2_1 _6326_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[15] ),
    .A1(_2428_),
    .S(net564),
    .X(_0822_));
 sky130_fd_sc_hd__mux2_1 _6327_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[16] ),
    .A1(_2429_),
    .S(net563),
    .X(_0823_));
 sky130_fd_sc_hd__mux2_1 _6328_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[17] ),
    .A1(_2430_),
    .S(net562),
    .X(_0824_));
 sky130_fd_sc_hd__mux2_1 _6329_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[18] ),
    .A1(_2431_),
    .S(net569),
    .X(_0825_));
 sky130_fd_sc_hd__mux2_1 _6330_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[19] ),
    .A1(_2432_),
    .S(net570),
    .X(_0826_));
 sky130_fd_sc_hd__mux2_1 _6331_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[20] ),
    .A1(_2433_),
    .S(net571),
    .X(_0827_));
 sky130_fd_sc_hd__mux2_1 _6332_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[21] ),
    .A1(_2434_),
    .S(net570),
    .X(_0828_));
 sky130_fd_sc_hd__mux2_1 _6333_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[22] ),
    .A1(_2435_),
    .S(net570),
    .X(_0829_));
 sky130_fd_sc_hd__mux2_1 _6334_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[23] ),
    .A1(_2436_),
    .S(net571),
    .X(_0830_));
 sky130_fd_sc_hd__mux2_1 _6335_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[24] ),
    .A1(_2437_),
    .S(net570),
    .X(_0831_));
 sky130_fd_sc_hd__mux2_1 _6336_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[25] ),
    .A1(_2438_),
    .S(net563),
    .X(_0832_));
 sky130_fd_sc_hd__mux2_1 _6337_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[26] ),
    .A1(_2439_),
    .S(net567),
    .X(_0833_));
 sky130_fd_sc_hd__mux2_1 _6338_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[27] ),
    .A1(_2440_),
    .S(net569),
    .X(_0834_));
 sky130_fd_sc_hd__mux2_1 _6339_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[28] ),
    .A1(_2441_),
    .S(net567),
    .X(_0835_));
 sky130_fd_sc_hd__mux2_1 _6340_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[29] ),
    .A1(net1958),
    .S(net569),
    .X(_0836_));
 sky130_fd_sc_hd__mux2_1 _6341_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[30] ),
    .A1(_2443_),
    .S(net565),
    .X(_0837_));
 sky130_fd_sc_hd__mux2_1 _6342_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[31] ),
    .A1(_2444_),
    .S(net568),
    .X(_0838_));
 sky130_fd_sc_hd__mux2_1 _6343_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[32] ),
    .A1(_2445_),
    .S(net569),
    .X(_0839_));
 sky130_fd_sc_hd__mux2_1 _6344_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[33] ),
    .A1(_2446_),
    .S(net567),
    .X(_0840_));
 sky130_fd_sc_hd__mux2_1 _6345_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[34] ),
    .A1(_2447_),
    .S(net565),
    .X(_0841_));
 sky130_fd_sc_hd__mux2_1 _6346_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[35] ),
    .A1(_2448_),
    .S(net568),
    .X(_0842_));
 sky130_fd_sc_hd__mux2_1 _6347_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[36] ),
    .A1(_2449_),
    .S(net565),
    .X(_0843_));
 sky130_fd_sc_hd__mux2_1 _6348_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[37] ),
    .A1(_2450_),
    .S(net570),
    .X(_0844_));
 sky130_fd_sc_hd__mux2_1 _6349_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[38] ),
    .A1(_2451_),
    .S(net565),
    .X(_0845_));
 sky130_fd_sc_hd__mux2_1 _6350_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[39] ),
    .A1(_2452_),
    .S(net570),
    .X(_0846_));
 sky130_fd_sc_hd__mux2_1 _6351_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[40] ),
    .A1(_2453_),
    .S(net565),
    .X(_0847_));
 sky130_fd_sc_hd__mux2_1 _6352_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[41] ),
    .A1(_2454_),
    .S(net565),
    .X(_0848_));
 sky130_fd_sc_hd__mux2_1 _6353_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[42] ),
    .A1(_2455_),
    .S(net568),
    .X(_0849_));
 sky130_fd_sc_hd__mux2_1 _6354_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[43] ),
    .A1(_2456_),
    .S(net567),
    .X(_0850_));
 sky130_fd_sc_hd__mux2_1 _6355_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[44] ),
    .A1(_2457_),
    .S(net568),
    .X(_0851_));
 sky130_fd_sc_hd__mux2_1 _6356_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[45] ),
    .A1(_2458_),
    .S(net568),
    .X(_0852_));
 sky130_fd_sc_hd__mux2_1 _6357_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[46] ),
    .A1(_2459_),
    .S(net564),
    .X(_0853_));
 sky130_fd_sc_hd__mux2_1 _6358_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[47] ),
    .A1(_2460_),
    .S(net568),
    .X(_0854_));
 sky130_fd_sc_hd__mux2_1 _6359_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[48] ),
    .A1(_2461_),
    .S(net570),
    .X(_0855_));
 sky130_fd_sc_hd__mux2_1 _6360_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[49] ),
    .A1(_2462_),
    .S(net565),
    .X(_0856_));
 sky130_fd_sc_hd__mux2_1 _6361_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[50] ),
    .A1(_2007_),
    .S(net569),
    .X(_0857_));
 sky130_fd_sc_hd__mux2_1 _6362_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[53] ),
    .A1(_2463_),
    .S(net566),
    .X(_0858_));
 sky130_fd_sc_hd__mux2_1 _6363_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[54] ),
    .A1(_2464_),
    .S(net568),
    .X(_0859_));
 sky130_fd_sc_hd__mux2_1 _6364_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[55] ),
    .A1(_2465_),
    .S(net567),
    .X(_0860_));
 sky130_fd_sc_hd__mux2_1 _6365_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[56] ),
    .A1(_2466_),
    .S(net567),
    .X(_0861_));
 sky130_fd_sc_hd__mux2_1 _6366_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[57] ),
    .A1(_2467_),
    .S(net566),
    .X(_0862_));
 sky130_fd_sc_hd__mux2_1 _6367_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[58] ),
    .A1(_2468_),
    .S(net562),
    .X(_0863_));
 sky130_fd_sc_hd__mux2_1 _6368_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[59] ),
    .A1(_2469_),
    .S(net567),
    .X(_0864_));
 sky130_fd_sc_hd__mux2_1 _6369_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[60] ),
    .A1(_2470_),
    .S(net563),
    .X(_0865_));
 sky130_fd_sc_hd__mux2_1 _6370_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[61] ),
    .A1(_2471_),
    .S(net563),
    .X(_0866_));
 sky130_fd_sc_hd__mux2_1 _6371_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[62] ),
    .A1(_2472_),
    .S(net563),
    .X(_0867_));
 sky130_fd_sc_hd__mux2_1 _6372_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[63] ),
    .A1(_2473_),
    .S(net565),
    .X(_0868_));
 sky130_fd_sc_hd__mux2_1 _6373_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[64] ),
    .A1(_2474_),
    .S(net571),
    .X(_0869_));
 sky130_fd_sc_hd__mux2_1 _6374_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[65] ),
    .A1(_2475_),
    .S(net564),
    .X(_0870_));
 sky130_fd_sc_hd__mux2_1 _6375_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[66] ),
    .A1(_2476_),
    .S(net562),
    .X(_0871_));
 sky130_fd_sc_hd__mux2_1 _6376_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[67] ),
    .A1(_2477_),
    .S(net564),
    .X(_0872_));
 sky130_fd_sc_hd__mux2_1 _6377_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[68] ),
    .A1(_2478_),
    .S(net564),
    .X(_0873_));
 sky130_fd_sc_hd__mux2_1 _6378_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[69] ),
    .A1(_2479_),
    .S(net564),
    .X(_0874_));
 sky130_fd_sc_hd__mux2_1 _6379_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[70] ),
    .A1(_2480_),
    .S(net562),
    .X(_0875_));
 sky130_fd_sc_hd__mux2_1 _6380_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[71] ),
    .A1(_2481_),
    .S(net563),
    .X(_0876_));
 sky130_fd_sc_hd__mux2_1 _6381_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[72] ),
    .A1(_2482_),
    .S(net566),
    .X(_0877_));
 sky130_fd_sc_hd__mux2_1 _6382_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[73] ),
    .A1(_2483_),
    .S(net568),
    .X(_0878_));
 sky130_fd_sc_hd__mux2_1 _6383_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[74] ),
    .A1(_2484_),
    .S(net562),
    .X(_0879_));
 sky130_fd_sc_hd__mux2_1 _6384_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[75] ),
    .A1(_2485_),
    .S(net563),
    .X(_0880_));
 sky130_fd_sc_hd__mux2_1 _6385_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[76] ),
    .A1(_2486_),
    .S(net562),
    .X(_0881_));
 sky130_fd_sc_hd__mux2_1 _6386_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[77] ),
    .A1(_2487_),
    .S(net562),
    .X(_0882_));
 sky130_fd_sc_hd__mux2_1 _6387_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[78] ),
    .A1(_2488_),
    .S(net563),
    .X(_0883_));
 sky130_fd_sc_hd__mux2_1 _6388_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[79] ),
    .A1(_2489_),
    .S(net563),
    .X(_0884_));
 sky130_fd_sc_hd__mux2_1 _6389_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[80] ),
    .A1(_2490_),
    .S(net562),
    .X(_0885_));
 sky130_fd_sc_hd__mux2_1 _6390_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[81] ),
    .A1(_2491_),
    .S(net562),
    .X(_0886_));
 sky130_fd_sc_hd__mux2_1 _6391_ (.A0(\u_s0.u_sync_wbb.s_cmd_rd_data_l[82] ),
    .A1(_2492_),
    .S(net562),
    .X(_0887_));
 sky130_fd_sc_hd__or3b_2 _6392_ (.A(_1704_),
    .B(net427),
    .C_N(net389),
    .X(_3249_));
 sky130_fd_sc_hd__inv_2 _6393_ (.A(_3249_),
    .Y(_3250_));
 sky130_fd_sc_hd__and3_1 _6394_ (.A(\u_s1.u_sync_wbb.u_resp_if.wr_ptr[0] ),
    .B(\u_s1.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .C(_3250_),
    .X(_3251_));
 sky130_fd_sc_hd__mux2_1 _6395_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][0] ),
    .A1(net1913),
    .S(net492),
    .X(_0888_));
 sky130_fd_sc_hd__mux2_1 _6396_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][1] ),
    .A1(net1924),
    .S(net493),
    .X(_0889_));
 sky130_fd_sc_hd__mux2_1 _6397_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][2] ),
    .A1(net1929),
    .S(net493),
    .X(_0890_));
 sky130_fd_sc_hd__mux2_1 _6398_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][3] ),
    .A1(net1850),
    .S(net491),
    .X(_0891_));
 sky130_fd_sc_hd__mux2_1 _6399_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][4] ),
    .A1(net1911),
    .S(net492),
    .X(_0892_));
 sky130_fd_sc_hd__mux2_1 _6400_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][5] ),
    .A1(net1936),
    .S(net492),
    .X(_0893_));
 sky130_fd_sc_hd__mux2_1 _6401_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][6] ),
    .A1(net1942),
    .S(net492),
    .X(_0894_));
 sky130_fd_sc_hd__mux2_1 _6402_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][7] ),
    .A1(net1906),
    .S(net492),
    .X(_0895_));
 sky130_fd_sc_hd__mux2_1 _6403_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][8] ),
    .A1(net1938),
    .S(net493),
    .X(_0896_));
 sky130_fd_sc_hd__mux2_1 _6404_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][9] ),
    .A1(net1910),
    .S(net492),
    .X(_0897_));
 sky130_fd_sc_hd__mux2_1 _6405_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][10] ),
    .A1(net2044),
    .S(net490),
    .X(_0898_));
 sky130_fd_sc_hd__mux2_1 _6406_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][11] ),
    .A1(net1864),
    .S(net491),
    .X(_0899_));
 sky130_fd_sc_hd__mux2_1 _6407_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][12] ),
    .A1(net1905),
    .S(net491),
    .X(_0900_));
 sky130_fd_sc_hd__mux2_1 _6408_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][13] ),
    .A1(net1856),
    .S(net491),
    .X(_0901_));
 sky130_fd_sc_hd__mux2_1 _6409_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][14] ),
    .A1(net1914),
    .S(net492),
    .X(_0902_));
 sky130_fd_sc_hd__mux2_1 _6410_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][15] ),
    .A1(net1920),
    .S(net492),
    .X(_0903_));
 sky130_fd_sc_hd__mux2_1 _6411_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][16] ),
    .A1(net1921),
    .S(net492),
    .X(_0904_));
 sky130_fd_sc_hd__mux2_1 _6412_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][17] ),
    .A1(net1860),
    .S(net491),
    .X(_0905_));
 sky130_fd_sc_hd__mux2_1 _6413_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][18] ),
    .A1(net1923),
    .S(net493),
    .X(_0906_));
 sky130_fd_sc_hd__mux2_1 _6414_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][19] ),
    .A1(net1877),
    .S(net490),
    .X(_0907_));
 sky130_fd_sc_hd__mux2_1 _6415_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][20] ),
    .A1(net1857),
    .S(net491),
    .X(_0908_));
 sky130_fd_sc_hd__mux2_1 _6416_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][21] ),
    .A1(net1862),
    .S(net491),
    .X(_0909_));
 sky130_fd_sc_hd__mux2_1 _6417_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][22] ),
    .A1(net1871),
    .S(net490),
    .X(_0910_));
 sky130_fd_sc_hd__mux2_1 _6418_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][23] ),
    .A1(net1870),
    .S(net490),
    .X(_0911_));
 sky130_fd_sc_hd__mux2_1 _6419_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][24] ),
    .A1(net1875),
    .S(net490),
    .X(_0912_));
 sky130_fd_sc_hd__mux2_1 _6420_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][25] ),
    .A1(net1865),
    .S(net491),
    .X(_0913_));
 sky130_fd_sc_hd__mux2_1 _6421_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][26] ),
    .A1(net2048),
    .S(net490),
    .X(_0914_));
 sky130_fd_sc_hd__mux2_1 _6422_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][27] ),
    .A1(net1873),
    .S(net490),
    .X(_0915_));
 sky130_fd_sc_hd__mux2_1 _6423_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][28] ),
    .A1(net1861),
    .S(net490),
    .X(_0916_));
 sky130_fd_sc_hd__mux2_1 _6424_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][29] ),
    .A1(net1859),
    .S(net491),
    .X(_0917_));
 sky130_fd_sc_hd__mux2_1 _6425_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][30] ),
    .A1(net1872),
    .S(net490),
    .X(_0918_));
 sky130_fd_sc_hd__mux2_1 _6426_ (.A0(\u_s1.u_sync_wbb.u_resp_if.mem[3][31] ),
    .A1(net1863),
    .S(net490),
    .X(_0919_));
 sky130_fd_sc_hd__or3b_1 _6427_ (.A(_3249_),
    .B(\u_s1.u_sync_wbb.u_resp_if.wr_ptr[0] ),
    .C_N(\u_s1.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .X(_3252_));
 sky130_fd_sc_hd__mux2_1 _6428_ (.A0(net1913),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][0] ),
    .S(net531),
    .X(_0920_));
 sky130_fd_sc_hd__mux2_1 _6429_ (.A0(net1924),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][1] ),
    .S(net532),
    .X(_0921_));
 sky130_fd_sc_hd__mux2_1 _6430_ (.A0(net1929),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][2] ),
    .S(net531),
    .X(_0922_));
 sky130_fd_sc_hd__mux2_1 _6431_ (.A0(net1850),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][3] ),
    .S(net530),
    .X(_0923_));
 sky130_fd_sc_hd__mux2_1 _6432_ (.A0(net1911),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][4] ),
    .S(net531),
    .X(_0924_));
 sky130_fd_sc_hd__mux2_1 _6433_ (.A0(net1936),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][5] ),
    .S(net531),
    .X(_0925_));
 sky130_fd_sc_hd__mux2_1 _6434_ (.A0(net1942),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][6] ),
    .S(net531),
    .X(_0926_));
 sky130_fd_sc_hd__mux2_1 _6435_ (.A0(net1906),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][7] ),
    .S(net530),
    .X(_0927_));
 sky130_fd_sc_hd__mux2_1 _6436_ (.A0(net1938),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][8] ),
    .S(net532),
    .X(_0928_));
 sky130_fd_sc_hd__mux2_1 _6437_ (.A0(net1910),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][9] ),
    .S(net531),
    .X(_0929_));
 sky130_fd_sc_hd__mux2_1 _6438_ (.A0(net1876),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][10] ),
    .S(net529),
    .X(_0930_));
 sky130_fd_sc_hd__mux2_1 _6439_ (.A0(net1864),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][11] ),
    .S(net532),
    .X(_0931_));
 sky130_fd_sc_hd__mux2_1 _6440_ (.A0(net1905),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][12] ),
    .S(net530),
    .X(_0932_));
 sky130_fd_sc_hd__mux2_1 _6441_ (.A0(net1856),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][13] ),
    .S(net530),
    .X(_0933_));
 sky130_fd_sc_hd__mux2_1 _6442_ (.A0(net1914),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][14] ),
    .S(net531),
    .X(_0934_));
 sky130_fd_sc_hd__mux2_1 _6443_ (.A0(net1920),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][15] ),
    .S(net531),
    .X(_0935_));
 sky130_fd_sc_hd__mux2_1 _6444_ (.A0(net1921),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][16] ),
    .S(net531),
    .X(_0936_));
 sky130_fd_sc_hd__mux2_1 _6445_ (.A0(net1860),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][17] ),
    .S(net530),
    .X(_0937_));
 sky130_fd_sc_hd__mux2_1 _6446_ (.A0(net1923),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][18] ),
    .S(net531),
    .X(_0938_));
 sky130_fd_sc_hd__mux2_1 _6447_ (.A0(net1877),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][19] ),
    .S(net529),
    .X(_0939_));
 sky130_fd_sc_hd__mux2_1 _6448_ (.A0(net1857),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][20] ),
    .S(net530),
    .X(_0940_));
 sky130_fd_sc_hd__mux2_1 _6449_ (.A0(net1862),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][21] ),
    .S(net530),
    .X(_0941_));
 sky130_fd_sc_hd__mux2_1 _6450_ (.A0(net2033),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][22] ),
    .S(net529),
    .X(_0942_));
 sky130_fd_sc_hd__mux2_1 _6451_ (.A0(net1870),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][23] ),
    .S(net529),
    .X(_0943_));
 sky130_fd_sc_hd__mux2_1 _6452_ (.A0(net2045),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][24] ),
    .S(net529),
    .X(_0944_));
 sky130_fd_sc_hd__mux2_1 _6453_ (.A0(net1865),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][25] ),
    .S(net529),
    .X(_0945_));
 sky130_fd_sc_hd__mux2_1 _6454_ (.A0(net2048),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][26] ),
    .S(net529),
    .X(_0946_));
 sky130_fd_sc_hd__mux2_1 _6455_ (.A0(net1873),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][27] ),
    .S(net529),
    .X(_0947_));
 sky130_fd_sc_hd__mux2_1 _6456_ (.A0(net1861),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][28] ),
    .S(net530),
    .X(_0948_));
 sky130_fd_sc_hd__mux2_1 _6457_ (.A0(net1859),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][29] ),
    .S(net530),
    .X(_0949_));
 sky130_fd_sc_hd__mux2_1 _6458_ (.A0(net1872),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][30] ),
    .S(net529),
    .X(_0950_));
 sky130_fd_sc_hd__mux2_1 _6459_ (.A0(net1863),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[2][31] ),
    .S(net529),
    .X(_0951_));
 sky130_fd_sc_hd__or3_1 _6460_ (.A(_1675_),
    .B(\u_s1.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .C(_3249_),
    .X(_3253_));
 sky130_fd_sc_hd__mux2_1 _6461_ (.A0(net1913),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][0] ),
    .S(net527),
    .X(_0952_));
 sky130_fd_sc_hd__mux2_1 _6462_ (.A0(net1924),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][1] ),
    .S(net527),
    .X(_0953_));
 sky130_fd_sc_hd__mux2_1 _6463_ (.A0(net1929),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][2] ),
    .S(net527),
    .X(_0954_));
 sky130_fd_sc_hd__mux2_1 _6464_ (.A0(net1850),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][3] ),
    .S(net525),
    .X(_0955_));
 sky130_fd_sc_hd__mux2_1 _6465_ (.A0(net1911),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][4] ),
    .S(net527),
    .X(_0956_));
 sky130_fd_sc_hd__mux2_1 _6466_ (.A0(net1936),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][5] ),
    .S(net528),
    .X(_0957_));
 sky130_fd_sc_hd__mux2_1 _6467_ (.A0(net1942),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][6] ),
    .S(net527),
    .X(_0958_));
 sky130_fd_sc_hd__mux2_1 _6468_ (.A0(net1906),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][7] ),
    .S(net525),
    .X(_0959_));
 sky130_fd_sc_hd__mux2_1 _6469_ (.A0(net1938),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][8] ),
    .S(net527),
    .X(_0960_));
 sky130_fd_sc_hd__mux2_1 _6470_ (.A0(net1910),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][9] ),
    .S(net525),
    .X(_0961_));
 sky130_fd_sc_hd__mux2_1 _6471_ (.A0(net2044),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][10] ),
    .S(net526),
    .X(_0962_));
 sky130_fd_sc_hd__mux2_1 _6472_ (.A0(net1864),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][11] ),
    .S(net526),
    .X(_0963_));
 sky130_fd_sc_hd__mux2_1 _6473_ (.A0(net1905),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][12] ),
    .S(net528),
    .X(_0964_));
 sky130_fd_sc_hd__mux2_1 _6474_ (.A0(net1856),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][13] ),
    .S(net525),
    .X(_0965_));
 sky130_fd_sc_hd__mux2_1 _6475_ (.A0(net1914),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][14] ),
    .S(net527),
    .X(_0966_));
 sky130_fd_sc_hd__mux2_1 _6476_ (.A0(net1920),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][15] ),
    .S(net527),
    .X(_0967_));
 sky130_fd_sc_hd__mux2_1 _6477_ (.A0(net1921),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][16] ),
    .S(net527),
    .X(_0968_));
 sky130_fd_sc_hd__mux2_1 _6478_ (.A0(net1860),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][17] ),
    .S(net525),
    .X(_0969_));
 sky130_fd_sc_hd__mux2_1 _6479_ (.A0(net1923),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][18] ),
    .S(net527),
    .X(_0970_));
 sky130_fd_sc_hd__mux2_1 _6480_ (.A0(net2042),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][19] ),
    .S(net526),
    .X(_0971_));
 sky130_fd_sc_hd__mux2_1 _6481_ (.A0(net1857),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][20] ),
    .S(net525),
    .X(_0972_));
 sky130_fd_sc_hd__mux2_1 _6482_ (.A0(net1862),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][21] ),
    .S(net525),
    .X(_0973_));
 sky130_fd_sc_hd__mux2_1 _6483_ (.A0(net1871),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][22] ),
    .S(net526),
    .X(_0974_));
 sky130_fd_sc_hd__mux2_1 _6484_ (.A0(net1870),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][23] ),
    .S(net526),
    .X(_0975_));
 sky130_fd_sc_hd__mux2_1 _6485_ (.A0(net1875),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][24] ),
    .S(net526),
    .X(_0976_));
 sky130_fd_sc_hd__mux2_1 _6486_ (.A0(net1865),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][25] ),
    .S(net525),
    .X(_0977_));
 sky130_fd_sc_hd__mux2_1 _6487_ (.A0(net2048),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][26] ),
    .S(net526),
    .X(_0978_));
 sky130_fd_sc_hd__mux2_1 _6488_ (.A0(net1873),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][27] ),
    .S(net526),
    .X(_0979_));
 sky130_fd_sc_hd__mux2_1 _6489_ (.A0(net1861),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][28] ),
    .S(net526),
    .X(_0980_));
 sky130_fd_sc_hd__mux2_1 _6490_ (.A0(net1859),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][29] ),
    .S(net525),
    .X(_0981_));
 sky130_fd_sc_hd__mux2_1 _6491_ (.A0(net1872),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][30] ),
    .S(net526),
    .X(_0982_));
 sky130_fd_sc_hd__mux2_1 _6492_ (.A0(net1863),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[1][31] ),
    .S(net525),
    .X(_0983_));
 sky130_fd_sc_hd__or3_1 _6493_ (.A(\u_s1.u_sync_wbb.u_resp_if.wr_ptr[0] ),
    .B(\u_s1.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .C(_3249_),
    .X(_3254_));
 sky130_fd_sc_hd__mux2_1 _6494_ (.A0(net1913),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][0] ),
    .S(net523),
    .X(_0984_));
 sky130_fd_sc_hd__mux2_1 _6495_ (.A0(net1924),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][1] ),
    .S(net523),
    .X(_0985_));
 sky130_fd_sc_hd__mux2_1 _6496_ (.A0(net1929),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][2] ),
    .S(net524),
    .X(_0986_));
 sky130_fd_sc_hd__mux2_1 _6497_ (.A0(net1850),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][3] ),
    .S(net522),
    .X(_0987_));
 sky130_fd_sc_hd__mux2_1 _6498_ (.A0(net1911),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][4] ),
    .S(net523),
    .X(_0988_));
 sky130_fd_sc_hd__mux2_1 _6499_ (.A0(net1936),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][5] ),
    .S(net524),
    .X(_0989_));
 sky130_fd_sc_hd__mux2_1 _6500_ (.A0(net1942),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][6] ),
    .S(net523),
    .X(_0990_));
 sky130_fd_sc_hd__mux2_1 _6501_ (.A0(net1906),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][7] ),
    .S(net523),
    .X(_0991_));
 sky130_fd_sc_hd__mux2_1 _6502_ (.A0(net1938),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][8] ),
    .S(net524),
    .X(_0992_));
 sky130_fd_sc_hd__mux2_1 _6503_ (.A0(net1910),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][9] ),
    .S(net523),
    .X(_0993_));
 sky130_fd_sc_hd__mux2_1 _6504_ (.A0(net2044),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][10] ),
    .S(net521),
    .X(_0994_));
 sky130_fd_sc_hd__mux2_1 _6505_ (.A0(net1864),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][11] ),
    .S(net521),
    .X(_0995_));
 sky130_fd_sc_hd__mux2_1 _6506_ (.A0(net1905),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][12] ),
    .S(net522),
    .X(_0996_));
 sky130_fd_sc_hd__mux2_1 _6507_ (.A0(net1856),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][13] ),
    .S(net522),
    .X(_0997_));
 sky130_fd_sc_hd__mux2_1 _6508_ (.A0(net1914),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][14] ),
    .S(net523),
    .X(_0998_));
 sky130_fd_sc_hd__mux2_1 _6509_ (.A0(net1920),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][15] ),
    .S(net523),
    .X(_0999_));
 sky130_fd_sc_hd__mux2_1 _6510_ (.A0(net1921),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][16] ),
    .S(net523),
    .X(_1000_));
 sky130_fd_sc_hd__mux2_1 _6511_ (.A0(net1860),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][17] ),
    .S(net522),
    .X(_1001_));
 sky130_fd_sc_hd__mux2_1 _6512_ (.A0(net1923),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][18] ),
    .S(net523),
    .X(_1002_));
 sky130_fd_sc_hd__mux2_1 _6513_ (.A0(net1877),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][19] ),
    .S(net521),
    .X(_1003_));
 sky130_fd_sc_hd__mux2_1 _6514_ (.A0(net1857),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][20] ),
    .S(net522),
    .X(_1004_));
 sky130_fd_sc_hd__mux2_1 _6515_ (.A0(net1862),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][21] ),
    .S(net522),
    .X(_1005_));
 sky130_fd_sc_hd__mux2_1 _6516_ (.A0(net1871),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][22] ),
    .S(net521),
    .X(_1006_));
 sky130_fd_sc_hd__mux2_1 _6517_ (.A0(net1870),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][23] ),
    .S(net521),
    .X(_1007_));
 sky130_fd_sc_hd__mux2_1 _6518_ (.A0(net2045),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][24] ),
    .S(net521),
    .X(_1008_));
 sky130_fd_sc_hd__mux2_1 _6519_ (.A0(net1865),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][25] ),
    .S(net522),
    .X(_1009_));
 sky130_fd_sc_hd__mux2_1 _6520_ (.A0(net2048),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][26] ),
    .S(net521),
    .X(_1010_));
 sky130_fd_sc_hd__mux2_1 _6521_ (.A0(net1873),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][27] ),
    .S(net521),
    .X(_1011_));
 sky130_fd_sc_hd__mux2_1 _6522_ (.A0(net1861),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][28] ),
    .S(net522),
    .X(_1012_));
 sky130_fd_sc_hd__mux2_1 _6523_ (.A0(net1859),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][29] ),
    .S(net522),
    .X(_1013_));
 sky130_fd_sc_hd__mux2_1 _6524_ (.A0(net1872),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][30] ),
    .S(net521),
    .X(_1014_));
 sky130_fd_sc_hd__mux2_1 _6525_ (.A0(net1863),
    .A1(\u_s1.u_sync_wbb.u_resp_if.mem[0][31] ),
    .S(net521),
    .X(_1015_));
 sky130_fd_sc_hd__o21ai_1 _6526_ (.A1(_1758_),
    .A2(_1781_),
    .B1(_1783_),
    .Y(_3255_));
 sky130_fd_sc_hd__and3_1 _6527_ (.A(m1_wbd_stb_i),
    .B(_1767_),
    .C(_1768_),
    .X(_3256_));
 sky130_fd_sc_hd__nand2_1 _6528_ (.A(net1368),
    .B(_1758_),
    .Y(_3257_));
 sky130_fd_sc_hd__nand2_2 _6529_ (.A(m3_wbd_stb_i),
    .B(_2494_),
    .Y(_3258_));
 sky130_fd_sc_hd__o221a_1 _6530_ (.A1(_1732_),
    .A2(_1758_),
    .B1(_1781_),
    .B2(net1369),
    .C1(_1725_),
    .X(_3259_));
 sky130_fd_sc_hd__nor2_1 _6531_ (.A(_3258_),
    .B(_3259_),
    .Y(_3260_));
 sky130_fd_sc_hd__a31o_1 _6532_ (.A1(_1725_),
    .A2(_3256_),
    .A3(_3257_),
    .B1(_3260_),
    .X(_3261_));
 sky130_fd_sc_hd__a22o_1 _6533_ (.A1(net1372),
    .A2(_3255_),
    .B1(_3261_),
    .B2(_1783_),
    .X(_1016_));
 sky130_fd_sc_hd__a2bb2o_1 _6534_ (.A1_N(net1369),
    .A2_N(_1781_),
    .B1(_1758_),
    .B2(net1373),
    .X(_3262_));
 sky130_fd_sc_hd__a22o_1 _6535_ (.A1(net1369),
    .A2(_1758_),
    .B1(_3258_),
    .B2(_3262_),
    .X(_3263_));
 sky130_fd_sc_hd__a21oi_1 _6536_ (.A1(_1725_),
    .A2(_3256_),
    .B1(_3263_),
    .Y(_3264_));
 sky130_fd_sc_hd__mux2_1 _6537_ (.A0(net1368),
    .A1(_3264_),
    .S(_1783_),
    .X(_1017_));
 sky130_fd_sc_hd__nor2_2 _6538_ (.A(\u_s1.u_sync_wbb.m_state[1] ),
    .B(\u_s1.u_sync_wbb.m_state[2] ),
    .Y(_3265_));
 sky130_fd_sc_hd__or2_1 _6539_ (.A(\u_s1.u_sync_wbb.m_state[1] ),
    .B(\u_s1.u_sync_wbb.m_state[2] ),
    .X(_3266_));
 sky130_fd_sc_hd__nor2_1 _6540_ (.A(\u_s1.u_sync_wbb.m_state[0] ),
    .B(net976),
    .Y(_3267_));
 sky130_fd_sc_hd__mux2_1 _6541_ (.A0(net976),
    .A1(_2002_),
    .S(\u_s1.u_sync_wbb.m_state[0] ),
    .X(_3268_));
 sky130_fd_sc_hd__a31o_1 _6542_ (.A1(net732),
    .A2(_1883_),
    .A3(net978),
    .B1(_1895_),
    .X(_3269_));
 sky130_fd_sc_hd__mux2_1 _6543_ (.A0(\u_s1.u_sync_wbb.wbm_ack_o ),
    .A1(_3269_),
    .S(_3268_),
    .X(_1018_));
 sky130_fd_sc_hd__and2b_1 _6544_ (.A_N(_1995_),
    .B(_3268_),
    .X(_3270_));
 sky130_fd_sc_hd__nand2_1 _6545_ (.A(\u_s1.u_sync_wbb.m_state[1] ),
    .B(_1892_),
    .Y(_3271_));
 sky130_fd_sc_hd__o221a_1 _6546_ (.A1(\u_s1.u_sync_wbb.m_state[1] ),
    .A2(_1894_),
    .B1(_1902_),
    .B2(\u_s1.u_sync_wbb.wbm_lack_o ),
    .C1(_3271_),
    .X(_3272_));
 sky130_fd_sc_hd__a31o_1 _6547_ (.A1(net732),
    .A2(_1883_),
    .A3(_3265_),
    .B1(_3272_),
    .X(_3273_));
 sky130_fd_sc_hd__mux2_1 _6548_ (.A0(\u_s1.u_sync_wbb.wbm_lack_o ),
    .A1(_3273_),
    .S(_3270_),
    .X(_1019_));
 sky130_fd_sc_hd__nor2_1 _6549_ (.A(_1903_),
    .B(net976),
    .Y(_3274_));
 sky130_fd_sc_hd__nor2_1 _6550_ (.A(_1893_),
    .B(_3267_),
    .Y(_3275_));
 sky130_fd_sc_hd__o22a_1 _6551_ (.A1(_1895_),
    .A2(_3274_),
    .B1(_3275_),
    .B2(\u_s1.u_sync_wbb.m_cmd_wr_en ),
    .X(_1020_));
 sky130_fd_sc_hd__o21ba_1 _6552_ (.A1(_1692_),
    .A2(\u_s1.u_sync_wbb.m_state[0] ),
    .B1_N(_1903_),
    .X(_3276_));
 sky130_fd_sc_hd__mux2_1 _6553_ (.A0(_1893_),
    .A1(\u_s1.u_sync_wbb.m_resp_rd_en ),
    .S(_3276_),
    .X(_1021_));
 sky130_fd_sc_hd__a221oi_2 _6554_ (.A1(net1798),
    .A2(_1955_),
    .B1(_1981_),
    .B2(net1817),
    .C1(_1988_),
    .Y(_3277_));
 sky130_fd_sc_hd__o211ai_1 _6555_ (.A1(net997),
    .A2(_3277_),
    .B1(_2922_),
    .C1(net1827),
    .Y(_3278_));
 sky130_fd_sc_hd__xnor2_2 _6556_ (.A(net784),
    .B(net582),
    .Y(_3279_));
 sky130_fd_sc_hd__mux2_1 _6557_ (.A0(_1679_),
    .A1(_3279_),
    .S(net1799),
    .X(_3280_));
 sky130_fd_sc_hd__mux2_1 _6558_ (.A0(_3280_),
    .A1(\u_s2.u_sync_wbb.m_bl_cnt[0] ),
    .S(net488),
    .X(_1022_));
 sky130_fd_sc_hd__a21boi_1 _6559_ (.A1(net784),
    .A2(net583),
    .B1_N(net791),
    .Y(_3281_));
 sky130_fd_sc_hd__or3b_1 _6560_ (.A(net791),
    .B(net783),
    .C_N(net582),
    .X(_3282_));
 sky130_fd_sc_hd__and3b_1 _6561_ (.A_N(_3281_),
    .B(_3282_),
    .C(net997),
    .X(_3283_));
 sky130_fd_sc_hd__nand2_1 _6562_ (.A(\u_s2.u_sync_wbb.m_bl_cnt[0] ),
    .B(\u_s2.u_sync_wbb.m_bl_cnt[1] ),
    .Y(_3284_));
 sky130_fd_sc_hd__or2_1 _6563_ (.A(\u_s2.u_sync_wbb.m_bl_cnt[0] ),
    .B(\u_s2.u_sync_wbb.m_bl_cnt[1] ),
    .X(_3285_));
 sky130_fd_sc_hd__a31o_1 _6564_ (.A1(net996),
    .A2(_3284_),
    .A3(_3285_),
    .B1(net488),
    .X(_3286_));
 sky130_fd_sc_hd__a2bb2o_1 _6565_ (.A1_N(_3283_),
    .A2_N(_3286_),
    .B1(\u_s2.u_sync_wbb.m_bl_cnt[1] ),
    .B2(net489),
    .X(_1023_));
 sky130_fd_sc_hd__nor3_1 _6566_ (.A(net794),
    .B(net791),
    .C(net783),
    .Y(_3287_));
 sky130_fd_sc_hd__a21o_1 _6567_ (.A1(net582),
    .A2(_3287_),
    .B1(net996),
    .X(_3288_));
 sky130_fd_sc_hd__a21oi_1 _6568_ (.A1(net794),
    .A2(_3282_),
    .B1(_3288_),
    .Y(_3289_));
 sky130_fd_sc_hd__nand2_1 _6569_ (.A(\u_s2.u_sync_wbb.m_bl_cnt[2] ),
    .B(_3285_),
    .Y(_3290_));
 sky130_fd_sc_hd__or2_1 _6570_ (.A(\u_s2.u_sync_wbb.m_bl_cnt[2] ),
    .B(_3285_),
    .X(_3291_));
 sky130_fd_sc_hd__a31o_1 _6571_ (.A1(net996),
    .A2(_3290_),
    .A3(_3291_),
    .B1(net488),
    .X(_3292_));
 sky130_fd_sc_hd__a2bb2o_1 _6572_ (.A1_N(_3289_),
    .A2_N(_3292_),
    .B1(\u_s2.u_sync_wbb.m_bl_cnt[2] ),
    .B2(net488),
    .X(_1024_));
 sky130_fd_sc_hd__a21bo_1 _6573_ (.A1(net582),
    .A2(_3287_),
    .B1_N(net792),
    .X(_3293_));
 sky130_fd_sc_hd__nand3b_1 _6574_ (.A_N(net792),
    .B(net583),
    .C(_3287_),
    .Y(_3294_));
 sky130_fd_sc_hd__nand2_1 _6575_ (.A(\u_s2.u_sync_wbb.m_bl_cnt[3] ),
    .B(_3291_),
    .Y(_3295_));
 sky130_fd_sc_hd__or4_2 _6576_ (.A(\u_s2.u_sync_wbb.m_bl_cnt[0] ),
    .B(\u_s2.u_sync_wbb.m_bl_cnt[1] ),
    .C(\u_s2.u_sync_wbb.m_bl_cnt[3] ),
    .D(\u_s2.u_sync_wbb.m_bl_cnt[2] ),
    .X(_3296_));
 sky130_fd_sc_hd__and3_1 _6577_ (.A(net996),
    .B(_3295_),
    .C(_3296_),
    .X(_3297_));
 sky130_fd_sc_hd__a311o_1 _6578_ (.A1(net997),
    .A2(_3293_),
    .A3(_3294_),
    .B1(_3297_),
    .C1(net488),
    .X(_3298_));
 sky130_fd_sc_hd__a21bo_1 _6579_ (.A1(\u_s2.u_sync_wbb.m_bl_cnt[3] ),
    .A2(net488),
    .B1_N(_3298_),
    .X(_1025_));
 sky130_fd_sc_hd__nor2_4 _6580_ (.A(_1925_),
    .B(net783),
    .Y(_3299_));
 sky130_fd_sc_hd__a221o_1 _6581_ (.A1(net795),
    .A2(_3294_),
    .B1(_3299_),
    .B2(net582),
    .C1(net996),
    .X(_3300_));
 sky130_fd_sc_hd__a21oi_1 _6582_ (.A1(\u_s2.u_sync_wbb.m_bl_cnt[4] ),
    .A2(_3296_),
    .B1(net997),
    .Y(_3301_));
 sky130_fd_sc_hd__o21a_1 _6583_ (.A1(\u_s2.u_sync_wbb.m_bl_cnt[4] ),
    .A2(_3296_),
    .B1(_3301_),
    .X(_3302_));
 sky130_fd_sc_hd__nor2_1 _6584_ (.A(net488),
    .B(_3302_),
    .Y(_3303_));
 sky130_fd_sc_hd__a22o_1 _6585_ (.A1(\u_s2.u_sync_wbb.m_bl_cnt[4] ),
    .A2(net488),
    .B1(_3300_),
    .B2(_3303_),
    .X(_1026_));
 sky130_fd_sc_hd__a21oi_1 _6586_ (.A1(net584),
    .A2(_3299_),
    .B1(net787),
    .Y(_3304_));
 sky130_fd_sc_hd__a31o_1 _6587_ (.A1(net787),
    .A2(net584),
    .A3(_3299_),
    .B1(net996),
    .X(_3305_));
 sky130_fd_sc_hd__nor2_2 _6588_ (.A(_3304_),
    .B(_3305_),
    .Y(_3306_));
 sky130_fd_sc_hd__or3_1 _6589_ (.A(\u_s2.u_sync_wbb.m_bl_cnt[5] ),
    .B(\u_s2.u_sync_wbb.m_bl_cnt[4] ),
    .C(_3296_),
    .X(_3307_));
 sky130_fd_sc_hd__o21ai_1 _6590_ (.A1(\u_s2.u_sync_wbb.m_bl_cnt[4] ),
    .A2(_3296_),
    .B1(\u_s2.u_sync_wbb.m_bl_cnt[5] ),
    .Y(_3308_));
 sky130_fd_sc_hd__a31o_1 _6591_ (.A1(net996),
    .A2(_3307_),
    .A3(_3308_),
    .B1(net489),
    .X(_3309_));
 sky130_fd_sc_hd__a2bb2o_1 _6592_ (.A1_N(_3306_),
    .A2_N(_3309_),
    .B1(\u_s2.u_sync_wbb.m_bl_cnt[5] ),
    .B2(net489),
    .X(_1027_));
 sky130_fd_sc_hd__a31o_1 _6593_ (.A1(net787),
    .A2(net582),
    .A3(_3299_),
    .B1(_1930_),
    .X(_3310_));
 sky130_fd_sc_hd__nand4_1 _6594_ (.A(_1930_),
    .B(net787),
    .C(net582),
    .D(_3299_),
    .Y(_3311_));
 sky130_fd_sc_hd__or2_1 _6595_ (.A(\u_s2.u_sync_wbb.m_bl_cnt[6] ),
    .B(_3307_),
    .X(_3312_));
 sky130_fd_sc_hd__nand2_1 _6596_ (.A(\u_s2.u_sync_wbb.m_bl_cnt[6] ),
    .B(_3307_),
    .Y(_3313_));
 sky130_fd_sc_hd__and3_1 _6597_ (.A(_2921_),
    .B(_3312_),
    .C(_3313_),
    .X(_3314_));
 sky130_fd_sc_hd__a311o_2 _6598_ (.A1(net997),
    .A2(_3310_),
    .A3(_3311_),
    .B1(_3314_),
    .C1(net488),
    .X(_3315_));
 sky130_fd_sc_hd__a21bo_1 _6599_ (.A1(\u_s2.u_sync_wbb.m_bl_cnt[6] ),
    .A2(net489),
    .B1_N(_3315_),
    .X(_1028_));
 sky130_fd_sc_hd__a41o_1 _6600_ (.A1(_1930_),
    .A2(net787),
    .A3(net582),
    .A4(_3299_),
    .B1(_1928_),
    .X(_3316_));
 sky130_fd_sc_hd__or4b_4 _6601_ (.A(_1925_),
    .B(_1933_),
    .C(net783),
    .D_N(net584),
    .X(_3317_));
 sky130_fd_sc_hd__nand2_1 _6602_ (.A(\u_s2.u_sync_wbb.m_bl_cnt[7] ),
    .B(_3312_),
    .Y(_3318_));
 sky130_fd_sc_hd__or2_2 _6603_ (.A(\u_s2.u_sync_wbb.m_bl_cnt[7] ),
    .B(_3312_),
    .X(_3319_));
 sky130_fd_sc_hd__and3_1 _6604_ (.A(_2921_),
    .B(_3318_),
    .C(_3319_),
    .X(_3320_));
 sky130_fd_sc_hd__a311o_1 _6605_ (.A1(net997),
    .A2(_3316_),
    .A3(_3317_),
    .B1(_3320_),
    .C1(net488),
    .X(_3321_));
 sky130_fd_sc_hd__a21bo_1 _6606_ (.A1(\u_s2.u_sync_wbb.m_bl_cnt[7] ),
    .A2(net489),
    .B1_N(_3321_),
    .X(_1029_));
 sky130_fd_sc_hd__nor2_2 _6607_ (.A(net783),
    .B(_1940_),
    .Y(_3322_));
 sky130_fd_sc_hd__a21o_1 _6608_ (.A1(net584),
    .A2(_3322_),
    .B1(net996),
    .X(_3323_));
 sky130_fd_sc_hd__a21o_2 _6609_ (.A1(net790),
    .A2(_3317_),
    .B1(_3323_),
    .X(_3324_));
 sky130_fd_sc_hd__nand2_1 _6610_ (.A(\u_s2.u_sync_wbb.m_bl_cnt[8] ),
    .B(_3319_),
    .Y(_3325_));
 sky130_fd_sc_hd__or2_1 _6611_ (.A(\u_s2.u_sync_wbb.m_bl_cnt[8] ),
    .B(_3319_),
    .X(_3326_));
 sky130_fd_sc_hd__a31oi_1 _6612_ (.A1(net996),
    .A2(_3325_),
    .A3(_3326_),
    .B1(net489),
    .Y(_3327_));
 sky130_fd_sc_hd__a22o_1 _6613_ (.A1(\u_s2.u_sync_wbb.m_bl_cnt[8] ),
    .A2(net489),
    .B1(_3324_),
    .B2(_3327_),
    .X(_1030_));
 sky130_fd_sc_hd__a21oi_1 _6614_ (.A1(_2921_),
    .A2(_3326_),
    .B1(net489),
    .Y(_3328_));
 sky130_fd_sc_hd__a21boi_4 _6615_ (.A1(net582),
    .A2(_3322_),
    .B1_N(net785),
    .Y(_3329_));
 sky130_fd_sc_hd__and3b_2 _6616_ (.A_N(net785),
    .B(net582),
    .C(_3322_),
    .X(_3330_));
 sky130_fd_sc_hd__or3b_1 _6617_ (.A(net997),
    .B(_3326_),
    .C_N(\u_s2.u_sync_wbb.m_bl_cnt[9] ),
    .X(_3331_));
 sky130_fd_sc_hd__o31a_1 _6618_ (.A1(_2921_),
    .A2(_3329_),
    .A3(_3330_),
    .B1(_3331_),
    .X(_3332_));
 sky130_fd_sc_hd__o22a_1 _6619_ (.A1(\u_s2.u_sync_wbb.m_bl_cnt[9] ),
    .A2(_3328_),
    .B1(_3332_),
    .B2(net489),
    .X(_1031_));
 sky130_fd_sc_hd__xnor2_1 _6620_ (.A(\u_s1.u_sync_wbb.u_resp_if.wr_ptr[0] ),
    .B(_3249_),
    .Y(_1032_));
 sky130_fd_sc_hd__a21oi_1 _6621_ (.A1(\u_s1.u_sync_wbb.u_resp_if.wr_ptr[0] ),
    .A2(_3250_),
    .B1(\u_s1.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .Y(_3333_));
 sky130_fd_sc_hd__nor2_1 _6622_ (.A(net491),
    .B(_3333_),
    .Y(_1033_));
 sky130_fd_sc_hd__xor2_1 _6623_ (.A(\u_s1.u_sync_wbb.u_resp_if.wr_ptr[2] ),
    .B(net492),
    .X(_1034_));
 sky130_fd_sc_hd__or2_1 _6624_ (.A(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .B(\u_s1.u_sync_wbb.m_cmd_wr_en ),
    .X(_3334_));
 sky130_fd_sc_hd__and2_1 _6625_ (.A(_2799_),
    .B(_3334_),
    .X(_1035_));
 sky130_fd_sc_hd__nand2_1 _6626_ (.A(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .B(_2799_),
    .Y(_3335_));
 sky130_fd_sc_hd__nand2b_1 _6627_ (.A_N(net752),
    .B(_3335_),
    .Y(_1036_));
 sky130_fd_sc_hd__xor2_1 _6628_ (.A(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[2] ),
    .B(net1004),
    .X(_1037_));
 sky130_fd_sc_hd__or3b_4 _6629_ (.A(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .B(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .C_N(\u_s2.u_sync_wbb.m_cmd_wr_en ),
    .X(_3336_));
 sky130_fd_sc_hd__mux2_1 _6630_ (.A0(net791),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][1] ),
    .S(net974),
    .X(_1038_));
 sky130_fd_sc_hd__mux2_1 _6631_ (.A0(net794),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][2] ),
    .S(net974),
    .X(_1039_));
 sky130_fd_sc_hd__mux2_1 _6632_ (.A0(net792),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][3] ),
    .S(_3336_),
    .X(_1040_));
 sky130_fd_sc_hd__mux2_1 _6633_ (.A0(net795),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][4] ),
    .S(net975),
    .X(_1041_));
 sky130_fd_sc_hd__mux2_1 _6634_ (.A0(net786),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][5] ),
    .S(net969),
    .X(_1042_));
 sky130_fd_sc_hd__mux2_1 _6635_ (.A0(net788),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][6] ),
    .S(net973),
    .X(_1043_));
 sky130_fd_sc_hd__mux2_1 _6636_ (.A0(net789),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][7] ),
    .S(net970),
    .X(_1044_));
 sky130_fd_sc_hd__mux2_1 _6637_ (.A0(net790),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][8] ),
    .S(net971),
    .X(_1045_));
 sky130_fd_sc_hd__mux2_1 _6638_ (.A0(net785),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][9] ),
    .S(net973),
    .X(_1046_));
 sky130_fd_sc_hd__mux2_1 _6639_ (.A0(net677),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][14] ),
    .S(net975),
    .X(_1047_));
 sky130_fd_sc_hd__mux2_1 _6640_ (.A0(net675),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][15] ),
    .S(net975),
    .X(_1048_));
 sky130_fd_sc_hd__mux2_1 _6641_ (.A0(net673),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][16] ),
    .S(net974),
    .X(_1049_));
 sky130_fd_sc_hd__mux2_1 _6642_ (.A0(net672),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][17] ),
    .S(net970),
    .X(_1050_));
 sky130_fd_sc_hd__mux2_1 _6643_ (.A0(net671),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][18] ),
    .S(net972),
    .X(_1051_));
 sky130_fd_sc_hd__mux2_1 _6644_ (.A0(net670),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][19] ),
    .S(net971),
    .X(_1052_));
 sky130_fd_sc_hd__mux2_1 _6645_ (.A0(net669),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][20] ),
    .S(net975),
    .X(_1053_));
 sky130_fd_sc_hd__mux2_1 _6646_ (.A0(net667),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][21] ),
    .S(net973),
    .X(_1054_));
 sky130_fd_sc_hd__mux2_1 _6647_ (.A0(net666),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][22] ),
    .S(net975),
    .X(_1055_));
 sky130_fd_sc_hd__mux2_1 _6648_ (.A0(net665),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][23] ),
    .S(net971),
    .X(_1056_));
 sky130_fd_sc_hd__mux2_1 _6649_ (.A0(net664),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][24] ),
    .S(net971),
    .X(_1057_));
 sky130_fd_sc_hd__mux2_1 _6650_ (.A0(net663),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][25] ),
    .S(_3336_),
    .X(_1058_));
 sky130_fd_sc_hd__mux2_1 _6651_ (.A0(_3164_),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][26] ),
    .S(net970),
    .X(_1059_));
 sky130_fd_sc_hd__mux2_1 _6652_ (.A0(net662),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][27] ),
    .S(net972),
    .X(_1060_));
 sky130_fd_sc_hd__mux2_1 _6653_ (.A0(net661),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][28] ),
    .S(net975),
    .X(_1061_));
 sky130_fd_sc_hd__mux2_1 _6654_ (.A0(net660),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][29] ),
    .S(net969),
    .X(_1062_));
 sky130_fd_sc_hd__mux2_1 _6655_ (.A0(net659),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][30] ),
    .S(net972),
    .X(_1063_));
 sky130_fd_sc_hd__mux2_1 _6656_ (.A0(net658),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][31] ),
    .S(net969),
    .X(_1064_));
 sky130_fd_sc_hd__mux2_1 _6657_ (.A0(net657),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][32] ),
    .S(net973),
    .X(_1065_));
 sky130_fd_sc_hd__mux2_1 _6658_ (.A0(net656),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][33] ),
    .S(net973),
    .X(_1066_));
 sky130_fd_sc_hd__mux2_1 _6659_ (.A0(net655),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][34] ),
    .S(net974),
    .X(_1067_));
 sky130_fd_sc_hd__mux2_1 _6660_ (.A0(net654),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][35] ),
    .S(net973),
    .X(_1068_));
 sky130_fd_sc_hd__mux2_1 _6661_ (.A0(net652),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][36] ),
    .S(net974),
    .X(_1069_));
 sky130_fd_sc_hd__mux2_1 _6662_ (.A0(net651),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][37] ),
    .S(net975),
    .X(_1070_));
 sky130_fd_sc_hd__mux2_1 _6663_ (.A0(_3195_),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][38] ),
    .S(net970),
    .X(_1071_));
 sky130_fd_sc_hd__mux2_1 _6664_ (.A0(net650),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][39] ),
    .S(net969),
    .X(_1072_));
 sky130_fd_sc_hd__mux2_1 _6665_ (.A0(net649),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][40] ),
    .S(net969),
    .X(_1073_));
 sky130_fd_sc_hd__mux2_1 _6666_ (.A0(net648),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][41] ),
    .S(net969),
    .X(_1074_));
 sky130_fd_sc_hd__mux2_1 _6667_ (.A0(net647),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][42] ),
    .S(net971),
    .X(_1075_));
 sky130_fd_sc_hd__mux2_1 _6668_ (.A0(net645),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][43] ),
    .S(net971),
    .X(_1076_));
 sky130_fd_sc_hd__mux2_1 _6669_ (.A0(net644),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][44] ),
    .S(net975),
    .X(_1077_));
 sky130_fd_sc_hd__mux2_1 _6670_ (.A0(net643),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][45] ),
    .S(net973),
    .X(_1078_));
 sky130_fd_sc_hd__mux2_1 _6671_ (.A0(net642),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][46] ),
    .S(net969),
    .X(_1079_));
 sky130_fd_sc_hd__mux2_1 _6672_ (.A0(_3216_),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][47] ),
    .S(net969),
    .X(_1080_));
 sky130_fd_sc_hd__mux2_1 _6673_ (.A0(net641),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][48] ),
    .S(net973),
    .X(_1081_));
 sky130_fd_sc_hd__mux2_1 _6674_ (.A0(net640),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][49] ),
    .S(net969),
    .X(_1082_));
 sky130_fd_sc_hd__mux2_1 _6675_ (.A0(net726),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][50] ),
    .S(net973),
    .X(_1083_));
 sky130_fd_sc_hd__mux2_1 _6676_ (.A0(net585),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][53] ),
    .S(net970),
    .X(_1084_));
 sky130_fd_sc_hd__mux2_1 _6677_ (.A0(net639),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][54] ),
    .S(net973),
    .X(_1085_));
 sky130_fd_sc_hd__mux2_1 _6678_ (.A0(net638),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][55] ),
    .S(net971),
    .X(_1086_));
 sky130_fd_sc_hd__mux2_1 _6679_ (.A0(net637),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][56] ),
    .S(net971),
    .X(_1087_));
 sky130_fd_sc_hd__mux2_1 _6680_ (.A0(net636),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][57] ),
    .S(net971),
    .X(_1088_));
 sky130_fd_sc_hd__mux2_1 _6681_ (.A0(net635),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][58] ),
    .S(net970),
    .X(_1089_));
 sky130_fd_sc_hd__mux2_1 _6682_ (.A0(net633),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][59] ),
    .S(net971),
    .X(_1090_));
 sky130_fd_sc_hd__mux2_1 _6683_ (.A0(net632),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][60] ),
    .S(net970),
    .X(_1091_));
 sky130_fd_sc_hd__mux2_1 _6684_ (.A0(net631),
    .A1(\u_s2.u_sync_wbb.u_cmd_if.mem[0][61] ),
    .S(net969),
    .X(_1092_));
 sky130_fd_sc_hd__or4_1 _6685_ (.A(\u_s1.u_sync_wbb.s_cmd_rd_data_l[7] ),
    .B(\u_s1.u_sync_wbb.s_cmd_rd_data_l[6] ),
    .C(\u_s1.u_sync_wbb.s_cmd_rd_data_l[5] ),
    .D(\u_s1.u_sync_wbb.s_cmd_rd_data_l[4] ),
    .X(_3337_));
 sky130_fd_sc_hd__or4_1 _6686_ (.A(\u_s1.u_sync_wbb.s_cmd_rd_data_l[9] ),
    .B(\u_s1.u_sync_wbb.s_cmd_rd_data_l[8] ),
    .C(net775),
    .D(_3337_),
    .X(_3338_));
 sky130_fd_sc_hd__o41a_1 _6687_ (.A1(\u_s1.u_sync_wbb.s_cmd_rd_data_l[3] ),
    .A2(\u_s1.u_sync_wbb.s_cmd_rd_data_l[2] ),
    .A3(\u_s1.u_sync_wbb.s_cmd_rd_data_l[1] ),
    .A4(_3338_),
    .B1(_1703_),
    .X(_3339_));
 sky130_fd_sc_hd__or4_1 _6688_ (.A(_2792_),
    .B(_2793_),
    .C(_2794_),
    .D(_2795_),
    .X(_3340_));
 sky130_fd_sc_hd__or4b_1 _6689_ (.A(_2790_),
    .B(_3340_),
    .C(_2791_),
    .D_N(net775),
    .X(_3341_));
 sky130_fd_sc_hd__or4_1 _6690_ (.A(_2796_),
    .B(_2797_),
    .C(_2798_),
    .D(_3341_),
    .X(_3342_));
 sky130_fd_sc_hd__a32o_1 _6691_ (.A1(net389),
    .A2(_3339_),
    .A3(_3342_),
    .B1(_1704_),
    .B2(\u_s1.u_sync_wbb.wbs_burst ),
    .X(_1093_));
 sky130_fd_sc_hd__xor2_1 _6692_ (.A(net1361),
    .B(net1506),
    .X(_1094_));
 sky130_fd_sc_hd__a21oi_1 _6693_ (.A1(net1362),
    .A2(net1507),
    .B1(net1355),
    .Y(_3343_));
 sky130_fd_sc_hd__and3_1 _6694_ (.A(net1355),
    .B(net1362),
    .C(net1507),
    .X(_3344_));
 sky130_fd_sc_hd__nor2_1 _6695_ (.A(_3343_),
    .B(_3344_),
    .Y(_1095_));
 sky130_fd_sc_hd__xor2_1 _6696_ (.A(\u_s1.u_sync_wbb.u_cmd_if.rd_ptr[2] ),
    .B(_3344_),
    .X(_1096_));
 sky130_fd_sc_hd__xor2_1 _6697_ (.A(net1350),
    .B(\u_s1.u_sync_wbb.m_resp_rd_en ),
    .X(_1097_));
 sky130_fd_sc_hd__a21oi_1 _6698_ (.A1(net1349),
    .A2(\u_s1.u_sync_wbb.m_resp_rd_en ),
    .B1(net1345),
    .Y(_3345_));
 sky130_fd_sc_hd__and3_1 _6699_ (.A(net1346),
    .B(net1350),
    .C(\u_s1.u_sync_wbb.m_resp_rd_en ),
    .X(_3346_));
 sky130_fd_sc_hd__nor2_1 _6700_ (.A(_3345_),
    .B(_3346_),
    .Y(_1098_));
 sky130_fd_sc_hd__xor2_1 _6701_ (.A(\u_s1.u_sync_wbb.u_resp_if.rd_ptr[2] ),
    .B(_3346_),
    .X(_1099_));
 sky130_fd_sc_hd__nand2_1 _6702_ (.A(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .B(\u_s0.u_sync_wbb.m_cmd_wr_en ),
    .Y(_3347_));
 sky130_fd_sc_hd__and3_1 _6703_ (.A(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .B(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .C(\u_s0.u_sync_wbb.m_cmd_wr_en ),
    .X(_3348_));
 sky130_fd_sc_hd__mux2_1 _6704_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][0] ),
    .A1(_1786_),
    .S(net964),
    .X(_1100_));
 sky130_fd_sc_hd__mux2_1 _6705_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][1] ),
    .A1(_1789_),
    .S(net960),
    .X(_1101_));
 sky130_fd_sc_hd__mux2_1 _6706_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][2] ),
    .A1(_1792_),
    .S(net966),
    .X(_1102_));
 sky130_fd_sc_hd__mux2_1 _6707_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][3] ),
    .A1(_1794_),
    .S(net966),
    .X(_1103_));
 sky130_fd_sc_hd__mux2_1 _6708_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][4] ),
    .A1(_1793_),
    .S(net965),
    .X(_1104_));
 sky130_fd_sc_hd__mux2_1 _6709_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][5] ),
    .A1(net808),
    .S(net965),
    .X(_1105_));
 sky130_fd_sc_hd__mux2_1 _6710_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][6] ),
    .A1(_1797_),
    .S(net965),
    .X(_1106_));
 sky130_fd_sc_hd__mux2_1 _6711_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][7] ),
    .A1(_1796_),
    .S(net966),
    .X(_1107_));
 sky130_fd_sc_hd__mux2_1 _6712_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][8] ),
    .A1(_1799_),
    .S(net966),
    .X(_1108_));
 sky130_fd_sc_hd__mux2_1 _6713_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][9] ),
    .A1(_1787_),
    .S(net964),
    .X(_1109_));
 sky130_fd_sc_hd__mux2_1 _6714_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][14] ),
    .A1(_2948_),
    .S(net962),
    .X(_1110_));
 sky130_fd_sc_hd__mux2_1 _6715_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][15] ),
    .A1(_2951_),
    .S(net960),
    .X(_1111_));
 sky130_fd_sc_hd__mux2_1 _6716_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][16] ),
    .A1(_2954_),
    .S(net959),
    .X(_1112_));
 sky130_fd_sc_hd__mux2_1 _6717_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][17] ),
    .A1(_2957_),
    .S(net959),
    .X(_1113_));
 sky130_fd_sc_hd__mux2_1 _6718_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][18] ),
    .A1(_2960_),
    .S(net965),
    .X(_1114_));
 sky130_fd_sc_hd__mux2_1 _6719_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][19] ),
    .A1(_2962_),
    .S(net965),
    .X(_1115_));
 sky130_fd_sc_hd__mux2_1 _6720_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][20] ),
    .A1(_2964_),
    .S(net966),
    .X(_1116_));
 sky130_fd_sc_hd__mux2_1 _6721_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][21] ),
    .A1(_2966_),
    .S(net965),
    .X(_1117_));
 sky130_fd_sc_hd__mux2_1 _6722_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][22] ),
    .A1(net2007),
    .S(net964),
    .X(_1118_));
 sky130_fd_sc_hd__mux2_1 _6723_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][23] ),
    .A1(_2971_),
    .S(net965),
    .X(_1119_));
 sky130_fd_sc_hd__mux2_1 _6724_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][24] ),
    .A1(_2973_),
    .S(net967),
    .X(_1120_));
 sky130_fd_sc_hd__mux2_1 _6725_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][25] ),
    .A1(_2976_),
    .S(net962),
    .X(_1121_));
 sky130_fd_sc_hd__mux2_1 _6726_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][26] ),
    .A1(_2979_),
    .S(net964),
    .X(_1122_));
 sky130_fd_sc_hd__mux2_1 _6727_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][27] ),
    .A1(_2981_),
    .S(net966),
    .X(_1123_));
 sky130_fd_sc_hd__mux2_1 _6728_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][28] ),
    .A1(_2983_),
    .S(net966),
    .X(_1124_));
 sky130_fd_sc_hd__mux2_1 _6729_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][29] ),
    .A1(_2985_),
    .S(net965),
    .X(_1125_));
 sky130_fd_sc_hd__mux2_1 _6730_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][30] ),
    .A1(_2988_),
    .S(net960),
    .X(_1126_));
 sky130_fd_sc_hd__mux2_1 _6731_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][31] ),
    .A1(_2991_),
    .S(net963),
    .X(_1127_));
 sky130_fd_sc_hd__mux2_1 _6732_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][32] ),
    .A1(_2993_),
    .S(net966),
    .X(_1128_));
 sky130_fd_sc_hd__mux2_1 _6733_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][33] ),
    .A1(_2995_),
    .S(net964),
    .X(_1129_));
 sky130_fd_sc_hd__mux2_1 _6734_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][34] ),
    .A1(_2998_),
    .S(net962),
    .X(_1130_));
 sky130_fd_sc_hd__mux2_1 _6735_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][35] ),
    .A1(_3001_),
    .S(net965),
    .X(_1131_));
 sky130_fd_sc_hd__mux2_1 _6736_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][36] ),
    .A1(_3004_),
    .S(net961),
    .X(_1132_));
 sky130_fd_sc_hd__mux2_1 _6737_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][37] ),
    .A1(net2009),
    .S(net964),
    .X(_1133_));
 sky130_fd_sc_hd__mux2_1 _6738_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][38] ),
    .A1(_3010_),
    .S(net960),
    .X(_1134_));
 sky130_fd_sc_hd__mux2_1 _6739_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][39] ),
    .A1(_3012_),
    .S(net964),
    .X(_1135_));
 sky130_fd_sc_hd__mux2_1 _6740_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][40] ),
    .A1(_3014_),
    .S(net963),
    .X(_1136_));
 sky130_fd_sc_hd__mux2_1 _6741_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][41] ),
    .A1(_3016_),
    .S(net967),
    .X(_1137_));
 sky130_fd_sc_hd__mux2_1 _6742_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][42] ),
    .A1(net2017),
    .S(net968),
    .X(_1138_));
 sky130_fd_sc_hd__mux2_1 _6743_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][43] ),
    .A1(net2038),
    .S(net964),
    .X(_1139_));
 sky130_fd_sc_hd__mux2_1 _6744_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][44] ),
    .A1(_3024_),
    .S(net963),
    .X(_1140_));
 sky130_fd_sc_hd__mux2_1 _6745_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][45] ),
    .A1(_3026_),
    .S(net968),
    .X(_1141_));
 sky130_fd_sc_hd__mux2_1 _6746_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][46] ),
    .A1(_3029_),
    .S(net959),
    .X(_1142_));
 sky130_fd_sc_hd__mux2_1 _6747_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][47] ),
    .A1(_3031_),
    .S(net962),
    .X(_1143_));
 sky130_fd_sc_hd__mux2_1 _6748_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][48] ),
    .A1(_3033_),
    .S(net964),
    .X(_1144_));
 sky130_fd_sc_hd__mux2_1 _6749_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][49] ),
    .A1(net2058),
    .S(net959),
    .X(_1145_));
 sky130_fd_sc_hd__mux2_1 _6750_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][50] ),
    .A1(_1806_),
    .S(net964),
    .X(_1146_));
 sky130_fd_sc_hd__mux2_1 _6751_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][53] ),
    .A1(_3038_),
    .S(net962),
    .X(_1147_));
 sky130_fd_sc_hd__mux2_1 _6752_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][54] ),
    .A1(_3041_),
    .S(net962),
    .X(_1148_));
 sky130_fd_sc_hd__mux2_1 _6753_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][55] ),
    .A1(_3044_),
    .S(net962),
    .X(_1149_));
 sky130_fd_sc_hd__mux2_1 _6754_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][56] ),
    .A1(_3047_),
    .S(net962),
    .X(_1150_));
 sky130_fd_sc_hd__mux2_1 _6755_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][57] ),
    .A1(_3050_),
    .S(net961),
    .X(_1151_));
 sky130_fd_sc_hd__mux2_1 _6756_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][58] ),
    .A1(_3053_),
    .S(net958),
    .X(_1152_));
 sky130_fd_sc_hd__mux2_1 _6757_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][59] ),
    .A1(net2022),
    .S(net962),
    .X(_1153_));
 sky130_fd_sc_hd__mux2_1 _6758_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][60] ),
    .A1(_3059_),
    .S(net963),
    .X(_1154_));
 sky130_fd_sc_hd__mux2_1 _6759_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][61] ),
    .A1(_3062_),
    .S(net962),
    .X(_1155_));
 sky130_fd_sc_hd__mux2_1 _6760_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][62] ),
    .A1(_3065_),
    .S(net960),
    .X(_1156_));
 sky130_fd_sc_hd__mux2_1 _6761_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][63] ),
    .A1(_3068_),
    .S(net963),
    .X(_1157_));
 sky130_fd_sc_hd__mux2_1 _6762_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][64] ),
    .A1(_3071_),
    .S(net960),
    .X(_1158_));
 sky130_fd_sc_hd__mux2_1 _6763_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][65] ),
    .A1(net1998),
    .S(net958),
    .X(_1159_));
 sky130_fd_sc_hd__mux2_1 _6764_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][66] ),
    .A1(net1869),
    .S(net958),
    .X(_1160_));
 sky130_fd_sc_hd__mux2_1 _6765_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][67] ),
    .A1(_3080_),
    .S(net963),
    .X(_1161_));
 sky130_fd_sc_hd__mux2_1 _6766_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][68] ),
    .A1(_3083_),
    .S(net963),
    .X(_1162_));
 sky130_fd_sc_hd__mux2_1 _6767_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][69] ),
    .A1(_3086_),
    .S(net958),
    .X(_1163_));
 sky130_fd_sc_hd__mux2_1 _6768_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][70] ),
    .A1(_3089_),
    .S(net958),
    .X(_1164_));
 sky130_fd_sc_hd__mux2_1 _6769_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][71] ),
    .A1(_3092_),
    .S(net963),
    .X(_1165_));
 sky130_fd_sc_hd__mux2_1 _6770_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][72] ),
    .A1(_3095_),
    .S(net960),
    .X(_1166_));
 sky130_fd_sc_hd__mux2_1 _6771_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][73] ),
    .A1(_3098_),
    .S(net963),
    .X(_1167_));
 sky130_fd_sc_hd__mux2_1 _6772_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][74] ),
    .A1(_3101_),
    .S(net958),
    .X(_1168_));
 sky130_fd_sc_hd__mux2_1 _6773_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][75] ),
    .A1(_3104_),
    .S(net960),
    .X(_1169_));
 sky130_fd_sc_hd__mux2_1 _6774_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][76] ),
    .A1(_3107_),
    .S(net960),
    .X(_1170_));
 sky130_fd_sc_hd__mux2_1 _6775_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][77] ),
    .A1(_3110_),
    .S(net958),
    .X(_1171_));
 sky130_fd_sc_hd__mux2_1 _6776_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][78] ),
    .A1(_3113_),
    .S(net958),
    .X(_1172_));
 sky130_fd_sc_hd__mux2_1 _6777_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][79] ),
    .A1(net1901),
    .S(net960),
    .X(_1173_));
 sky130_fd_sc_hd__mux2_1 _6778_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][80] ),
    .A1(_3119_),
    .S(net958),
    .X(_1174_));
 sky130_fd_sc_hd__mux2_1 _6779_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][81] ),
    .A1(net1867),
    .S(net958),
    .X(_1175_));
 sky130_fd_sc_hd__mux2_1 _6780_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[3][82] ),
    .A1(net1853),
    .S(net959),
    .X(_1176_));
 sky130_fd_sc_hd__and3b_1 _6781_ (.A_N(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .B(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .C(\u_s2.u_sync_wbb.m_cmd_wr_en ),
    .X(_3349_));
 sky130_fd_sc_hd__mux2_1 _6782_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][1] ),
    .A1(net791),
    .S(net955),
    .X(_1177_));
 sky130_fd_sc_hd__mux2_1 _6783_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][2] ),
    .A1(net794),
    .S(net955),
    .X(_1178_));
 sky130_fd_sc_hd__mux2_1 _6784_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][3] ),
    .A1(net792),
    .S(net957),
    .X(_1179_));
 sky130_fd_sc_hd__mux2_1 _6785_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][4] ),
    .A1(net795),
    .S(net956),
    .X(_1180_));
 sky130_fd_sc_hd__mux2_1 _6786_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][5] ),
    .A1(net786),
    .S(net951),
    .X(_1181_));
 sky130_fd_sc_hd__mux2_1 _6787_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][6] ),
    .A1(net788),
    .S(net955),
    .X(_1182_));
 sky130_fd_sc_hd__mux2_1 _6788_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][7] ),
    .A1(net789),
    .S(net952),
    .X(_1183_));
 sky130_fd_sc_hd__mux2_1 _6789_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][8] ),
    .A1(net790),
    .S(net954),
    .X(_1184_));
 sky130_fd_sc_hd__mux2_1 _6790_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][9] ),
    .A1(net785),
    .S(net955),
    .X(_1185_));
 sky130_fd_sc_hd__mux2_1 _6791_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][14] ),
    .A1(net677),
    .S(net957),
    .X(_1186_));
 sky130_fd_sc_hd__mux2_1 _6792_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][15] ),
    .A1(net675),
    .S(net956),
    .X(_1187_));
 sky130_fd_sc_hd__mux2_1 _6793_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][16] ),
    .A1(net673),
    .S(net955),
    .X(_1188_));
 sky130_fd_sc_hd__mux2_1 _6794_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][17] ),
    .A1(net672),
    .S(net952),
    .X(_1189_));
 sky130_fd_sc_hd__mux2_1 _6795_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][18] ),
    .A1(net671),
    .S(net953),
    .X(_1190_));
 sky130_fd_sc_hd__mux2_1 _6796_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][19] ),
    .A1(net670),
    .S(net952),
    .X(_1191_));
 sky130_fd_sc_hd__mux2_1 _6797_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][20] ),
    .A1(net669),
    .S(net956),
    .X(_1192_));
 sky130_fd_sc_hd__mux2_1 _6798_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][21] ),
    .A1(net667),
    .S(net953),
    .X(_1193_));
 sky130_fd_sc_hd__mux2_1 _6799_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][22] ),
    .A1(net666),
    .S(net956),
    .X(_1194_));
 sky130_fd_sc_hd__mux2_1 _6800_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][23] ),
    .A1(net665),
    .S(net952),
    .X(_1195_));
 sky130_fd_sc_hd__mux2_1 _6801_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][24] ),
    .A1(net664),
    .S(net954),
    .X(_1196_));
 sky130_fd_sc_hd__mux2_1 _6802_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][25] ),
    .A1(net663),
    .S(net957),
    .X(_1197_));
 sky130_fd_sc_hd__mux2_1 _6803_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][26] ),
    .A1(_3164_),
    .S(net952),
    .X(_1198_));
 sky130_fd_sc_hd__mux2_1 _6804_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][27] ),
    .A1(net662),
    .S(net953),
    .X(_1199_));
 sky130_fd_sc_hd__mux2_1 _6805_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][28] ),
    .A1(net661),
    .S(net955),
    .X(_1200_));
 sky130_fd_sc_hd__mux2_1 _6806_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][29] ),
    .A1(net660),
    .S(net952),
    .X(_1201_));
 sky130_fd_sc_hd__mux2_1 _6807_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][30] ),
    .A1(net659),
    .S(net953),
    .X(_1202_));
 sky130_fd_sc_hd__mux2_1 _6808_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][31] ),
    .A1(net658),
    .S(net951),
    .X(_1203_));
 sky130_fd_sc_hd__mux2_1 _6809_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][32] ),
    .A1(net657),
    .S(net956),
    .X(_1204_));
 sky130_fd_sc_hd__mux2_1 _6810_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][33] ),
    .A1(net656),
    .S(net955),
    .X(_1205_));
 sky130_fd_sc_hd__mux2_1 _6811_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][34] ),
    .A1(net655),
    .S(net955),
    .X(_1206_));
 sky130_fd_sc_hd__mux2_1 _6812_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][35] ),
    .A1(net654),
    .S(net955),
    .X(_1207_));
 sky130_fd_sc_hd__mux2_1 _6813_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][36] ),
    .A1(net652),
    .S(net956),
    .X(_1208_));
 sky130_fd_sc_hd__mux2_1 _6814_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][37] ),
    .A1(net651),
    .S(net956),
    .X(_1209_));
 sky130_fd_sc_hd__mux2_1 _6815_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][38] ),
    .A1(_3195_),
    .S(net951),
    .X(_1210_));
 sky130_fd_sc_hd__mux2_1 _6816_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][39] ),
    .A1(net650),
    .S(net951),
    .X(_1211_));
 sky130_fd_sc_hd__mux2_1 _6817_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][40] ),
    .A1(net649),
    .S(net953),
    .X(_1212_));
 sky130_fd_sc_hd__mux2_1 _6818_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][41] ),
    .A1(net648),
    .S(net951),
    .X(_1213_));
 sky130_fd_sc_hd__mux2_1 _6819_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][42] ),
    .A1(net647),
    .S(net952),
    .X(_1214_));
 sky130_fd_sc_hd__mux2_1 _6820_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][43] ),
    .A1(net645),
    .S(net953),
    .X(_1215_));
 sky130_fd_sc_hd__mux2_1 _6821_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][44] ),
    .A1(net644),
    .S(net956),
    .X(_1216_));
 sky130_fd_sc_hd__mux2_1 _6822_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][45] ),
    .A1(net643),
    .S(net956),
    .X(_1217_));
 sky130_fd_sc_hd__mux2_1 _6823_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][46] ),
    .A1(net642),
    .S(net951),
    .X(_1218_));
 sky130_fd_sc_hd__mux2_1 _6824_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][47] ),
    .A1(net2029),
    .S(net951),
    .X(_1219_));
 sky130_fd_sc_hd__mux2_1 _6825_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][48] ),
    .A1(net641),
    .S(net954),
    .X(_1220_));
 sky130_fd_sc_hd__mux2_1 _6826_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][49] ),
    .A1(net640),
    .S(net952),
    .X(_1221_));
 sky130_fd_sc_hd__mux2_1 _6827_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][50] ),
    .A1(net726),
    .S(net955),
    .X(_1222_));
 sky130_fd_sc_hd__mux2_1 _6828_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][53] ),
    .A1(net585),
    .S(net954),
    .X(_1223_));
 sky130_fd_sc_hd__mux2_1 _6829_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][54] ),
    .A1(net639),
    .S(net953),
    .X(_1224_));
 sky130_fd_sc_hd__mux2_1 _6830_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][55] ),
    .A1(net638),
    .S(net953),
    .X(_1225_));
 sky130_fd_sc_hd__mux2_1 _6831_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][56] ),
    .A1(net637),
    .S(net951),
    .X(_1226_));
 sky130_fd_sc_hd__mux2_1 _6832_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][57] ),
    .A1(net636),
    .S(net953),
    .X(_1227_));
 sky130_fd_sc_hd__mux2_1 _6833_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][58] ),
    .A1(net635),
    .S(net951),
    .X(_1228_));
 sky130_fd_sc_hd__mux2_1 _6834_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][59] ),
    .A1(net633),
    .S(net953),
    .X(_1229_));
 sky130_fd_sc_hd__mux2_1 _6835_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][60] ),
    .A1(net632),
    .S(net952),
    .X(_1230_));
 sky130_fd_sc_hd__mux2_1 _6836_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[2][61] ),
    .A1(net631),
    .S(net951),
    .X(_1231_));
 sky130_fd_sc_hd__and3b_2 _6837_ (.A_N(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .B(\u_s1.u_sync_wbb.m_cmd_wr_en ),
    .C(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .X(_3350_));
 sky130_fd_sc_hd__mux2_1 _6838_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][1] ),
    .A1(net797),
    .S(net946),
    .X(_1232_));
 sky130_fd_sc_hd__mux2_1 _6839_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][2] ),
    .A1(net798),
    .S(net944),
    .X(_1233_));
 sky130_fd_sc_hd__mux2_1 _6840_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][3] ),
    .A1(_1860_),
    .S(net945),
    .X(_1234_));
 sky130_fd_sc_hd__mux2_1 _6841_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][4] ),
    .A1(_1856_),
    .S(net944),
    .X(_1235_));
 sky130_fd_sc_hd__mux2_1 _6842_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][5] ),
    .A1(_1869_),
    .S(net948),
    .X(_1236_));
 sky130_fd_sc_hd__mux2_1 _6843_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][6] ),
    .A1(_1868_),
    .S(net947),
    .X(_1237_));
 sky130_fd_sc_hd__mux2_1 _6844_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][7] ),
    .A1(_1867_),
    .S(net944),
    .X(_1238_));
 sky130_fd_sc_hd__mux2_1 _6845_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][8] ),
    .A1(_1866_),
    .S(net947),
    .X(_1239_));
 sky130_fd_sc_hd__mux2_1 _6846_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][9] ),
    .A1(_1873_),
    .S(net944),
    .X(_1240_));
 sky130_fd_sc_hd__mux2_1 _6847_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][14] ),
    .A1(net686),
    .S(net948),
    .X(_1241_));
 sky130_fd_sc_hd__mux2_1 _6848_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][15] ),
    .A1(net685),
    .S(net945),
    .X(_1242_));
 sky130_fd_sc_hd__mux2_1 _6849_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][16] ),
    .A1(net684),
    .S(net945),
    .X(_1243_));
 sky130_fd_sc_hd__mux2_1 _6850_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][17] ),
    .A1(net683),
    .S(net947),
    .X(_1244_));
 sky130_fd_sc_hd__mux2_1 _6851_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][18] ),
    .A1(net682),
    .S(net949),
    .X(_1245_));
 sky130_fd_sc_hd__mux2_1 _6852_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][19] ),
    .A1(_2816_),
    .S(net947),
    .X(_1246_));
 sky130_fd_sc_hd__mux2_1 _6853_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][20] ),
    .A1(_2818_),
    .S(net950),
    .X(_1247_));
 sky130_fd_sc_hd__mux2_1 _6854_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][21] ),
    .A1(net681),
    .S(net947),
    .X(_1248_));
 sky130_fd_sc_hd__mux2_1 _6855_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][22] ),
    .A1(_2823_),
    .S(net948),
    .X(_1249_));
 sky130_fd_sc_hd__mux2_1 _6856_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][23] ),
    .A1(_2825_),
    .S(net948),
    .X(_1250_));
 sky130_fd_sc_hd__mux2_1 _6857_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][24] ),
    .A1(_2827_),
    .S(net946),
    .X(_1251_));
 sky130_fd_sc_hd__mux2_1 _6858_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][25] ),
    .A1(_2830_),
    .S(net948),
    .X(_1252_));
 sky130_fd_sc_hd__mux2_1 _6859_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][26] ),
    .A1(_2832_),
    .S(net948),
    .X(_1253_));
 sky130_fd_sc_hd__mux2_1 _6860_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][27] ),
    .A1(_2835_),
    .S(net949),
    .X(_1254_));
 sky130_fd_sc_hd__mux2_1 _6861_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][28] ),
    .A1(_2838_),
    .S(net949),
    .X(_1255_));
 sky130_fd_sc_hd__mux2_1 _6862_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][29] ),
    .A1(_2841_),
    .S(net948),
    .X(_1256_));
 sky130_fd_sc_hd__mux2_1 _6863_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][30] ),
    .A1(_2844_),
    .S(net949),
    .X(_1257_));
 sky130_fd_sc_hd__mux2_1 _6864_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][31] ),
    .A1(_2846_),
    .S(net946),
    .X(_1258_));
 sky130_fd_sc_hd__mux2_1 _6865_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][32] ),
    .A1(_2849_),
    .S(net947),
    .X(_1259_));
 sky130_fd_sc_hd__mux2_1 _6866_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][33] ),
    .A1(_2851_),
    .S(net944),
    .X(_1260_));
 sky130_fd_sc_hd__mux2_1 _6867_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][34] ),
    .A1(_2854_),
    .S(net947),
    .X(_1261_));
 sky130_fd_sc_hd__mux2_1 _6868_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][35] ),
    .A1(_2856_),
    .S(net948),
    .X(_1262_));
 sky130_fd_sc_hd__mux2_1 _6869_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][36] ),
    .A1(_2858_),
    .S(net945),
    .X(_1263_));
 sky130_fd_sc_hd__mux2_1 _6870_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][37] ),
    .A1(_2861_),
    .S(net947),
    .X(_1264_));
 sky130_fd_sc_hd__mux2_1 _6871_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][38] ),
    .A1(_2863_),
    .S(net947),
    .X(_1265_));
 sky130_fd_sc_hd__mux2_1 _6872_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][39] ),
    .A1(_2865_),
    .S(net944),
    .X(_1266_));
 sky130_fd_sc_hd__mux2_1 _6873_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][40] ),
    .A1(_2867_),
    .S(net945),
    .X(_1267_));
 sky130_fd_sc_hd__mux2_1 _6874_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][41] ),
    .A1(_2869_),
    .S(net947),
    .X(_1268_));
 sky130_fd_sc_hd__mux2_1 _6875_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][42] ),
    .A1(net680),
    .S(net948),
    .X(_1269_));
 sky130_fd_sc_hd__mux2_1 _6876_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][43] ),
    .A1(net2080),
    .S(net945),
    .X(_1270_));
 sky130_fd_sc_hd__mux2_1 _6877_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][44] ),
    .A1(_2875_),
    .S(net944),
    .X(_1271_));
 sky130_fd_sc_hd__mux2_1 _6878_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][45] ),
    .A1(_2877_),
    .S(net948),
    .X(_1272_));
 sky130_fd_sc_hd__mux2_1 _6879_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][46] ),
    .A1(net679),
    .S(net949),
    .X(_1273_));
 sky130_fd_sc_hd__mux2_1 _6880_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][47] ),
    .A1(_2881_),
    .S(net944),
    .X(_1274_));
 sky130_fd_sc_hd__mux2_1 _6881_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][48] ),
    .A1(_2883_),
    .S(net944),
    .X(_1275_));
 sky130_fd_sc_hd__mux2_1 _6882_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][49] ),
    .A1(_2885_),
    .S(net946),
    .X(_1276_));
 sky130_fd_sc_hd__mux2_1 _6883_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][50] ),
    .A1(net732),
    .S(net950),
    .X(_1277_));
 sky130_fd_sc_hd__mux2_1 _6884_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][53] ),
    .A1(_2888_),
    .S(net946),
    .X(_1278_));
 sky130_fd_sc_hd__mux2_1 _6885_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][54] ),
    .A1(_2891_),
    .S(net945),
    .X(_1279_));
 sky130_fd_sc_hd__mux2_1 _6886_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][55] ),
    .A1(_2894_),
    .S(net945),
    .X(_1280_));
 sky130_fd_sc_hd__mux2_1 _6887_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][56] ),
    .A1(_2897_),
    .S(net946),
    .X(_1281_));
 sky130_fd_sc_hd__mux2_1 _6888_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][57] ),
    .A1(_2900_),
    .S(net944),
    .X(_1282_));
 sky130_fd_sc_hd__mux2_1 _6889_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][58] ),
    .A1(_2903_),
    .S(net945),
    .X(_1283_));
 sky130_fd_sc_hd__mux2_1 _6890_ (.A0(\u_s1.u_sync_wbb.u_cmd_if.mem[2][59] ),
    .A1(_2906_),
    .S(net945),
    .X(_1284_));
 sky130_fd_sc_hd__and3b_1 _6891_ (.A_N(net619),
    .B(net604),
    .C(net592),
    .X(_3351_));
 sky130_fd_sc_hd__mux2_1 _6892_ (.A0(\u_reg.reg_7[24] ),
    .A1(net695),
    .S(net520),
    .X(_1285_));
 sky130_fd_sc_hd__mux2_1 _6893_ (.A0(\u_reg.reg_7[25] ),
    .A1(net693),
    .S(net520),
    .X(_1286_));
 sky130_fd_sc_hd__mux2_1 _6894_ (.A0(\u_reg.reg_7[26] ),
    .A1(net692),
    .S(net520),
    .X(_1287_));
 sky130_fd_sc_hd__mux2_1 _6895_ (.A0(\u_reg.reg_7[27] ),
    .A1(net691),
    .S(net520),
    .X(_1288_));
 sky130_fd_sc_hd__mux2_1 _6896_ (.A0(\u_reg.reg_7[28] ),
    .A1(net690),
    .S(net520),
    .X(_1289_));
 sky130_fd_sc_hd__mux2_1 _6897_ (.A0(\u_reg.reg_7[29] ),
    .A1(net689),
    .S(net520),
    .X(_1290_));
 sky130_fd_sc_hd__mux2_1 _6898_ (.A0(\u_reg.reg_7[30] ),
    .A1(net688),
    .S(net520),
    .X(_1291_));
 sky130_fd_sc_hd__mux2_1 _6899_ (.A0(\u_reg.reg_7[31] ),
    .A1(net687),
    .S(_3351_),
    .X(_1292_));
 sky130_fd_sc_hd__a21oi_2 _6900_ (.A1(\u_s0.u_sync_wbb.m_state[0] ),
    .A2(net580),
    .B1(_2591_),
    .Y(_3352_));
 sky130_fd_sc_hd__nor2_1 _6901_ (.A(_1784_),
    .B(net1005),
    .Y(_3353_));
 sky130_fd_sc_hd__and3b_1 _6902_ (.A_N(_1784_),
    .B(_1806_),
    .C(_2589_),
    .X(_3354_));
 sky130_fd_sc_hd__or2_1 _6903_ (.A(_1823_),
    .B(_3354_),
    .X(_3355_));
 sky130_fd_sc_hd__nor2_1 _6904_ (.A(_1821_),
    .B(_2591_),
    .Y(_3356_));
 sky130_fd_sc_hd__mux2_1 _6905_ (.A0(\u_s0.u_sync_wbb.wbm_ack_o ),
    .A1(_3355_),
    .S(_3352_),
    .X(_1293_));
 sky130_fd_sc_hd__o31a_1 _6906_ (.A1(_1803_),
    .A2(_1807_),
    .A3(_1913_),
    .B1(_3352_),
    .X(_3357_));
 sky130_fd_sc_hd__o221a_1 _6907_ (.A1(\u_s0.u_sync_wbb.m_state[1] ),
    .A2(_1822_),
    .B1(_1826_),
    .B2(\u_s0.u_sync_wbb.wbm_lack_o ),
    .C1(_2588_),
    .X(_3358_));
 sky130_fd_sc_hd__or2_1 _6908_ (.A(_3354_),
    .B(_3358_),
    .X(_3359_));
 sky130_fd_sc_hd__mux2_1 _6909_ (.A0(\u_s0.u_sync_wbb.wbm_lack_o ),
    .A1(_3359_),
    .S(_3357_),
    .X(_1294_));
 sky130_fd_sc_hd__o32a_1 _6910_ (.A1(_1823_),
    .A2(_2591_),
    .A3(_3353_),
    .B1(_3356_),
    .B2(\u_s0.u_sync_wbb.m_cmd_wr_en ),
    .X(_1295_));
 sky130_fd_sc_hd__o21ai_1 _6911_ (.A1(\u_s0.u_sync_wbb.m_state[1] ),
    .A2(\u_s0.u_sync_wbb.m_state[0] ),
    .B1(_1913_),
    .Y(_3360_));
 sky130_fd_sc_hd__a22o_1 _6912_ (.A1(_1821_),
    .A2(_1913_),
    .B1(_3360_),
    .B2(\u_s0.u_sync_wbb.m_resp_rd_en ),
    .X(_1296_));
 sky130_fd_sc_hd__a221o_1 _6913_ (.A1(\u_s1.u_sync_wbb.m_state[2] ),
    .A2(_1850_),
    .B1(_1892_),
    .B2(\u_s1.u_sync_wbb.m_state[1] ),
    .C1(_3267_),
    .X(_3361_));
 sky130_fd_sc_hd__a211o_1 _6914_ (.A1(_1902_),
    .A2(net976),
    .B1(_3361_),
    .C1(_1903_),
    .X(_3362_));
 sky130_fd_sc_hd__a21oi_4 _6915_ (.A1(net630),
    .A2(_2001_),
    .B1(_1875_),
    .Y(_3363_));
 sky130_fd_sc_hd__and3_1 _6916_ (.A(_1875_),
    .B(net630),
    .C(_2001_),
    .X(_3364_));
 sky130_fd_sc_hd__nand2_1 _6917_ (.A(\u_s1.u_sync_wbb.m_bl_cnt[0] ),
    .B(net977),
    .Y(_3365_));
 sky130_fd_sc_hd__o31a_1 _6918_ (.A1(net977),
    .A2(_3363_),
    .A3(_3364_),
    .B1(_3365_),
    .X(_3366_));
 sky130_fd_sc_hd__mux2_1 _6919_ (.A0(_3366_),
    .A1(\u_s1.u_sync_wbb.m_bl_cnt[0] ),
    .S(net486),
    .X(_1297_));
 sky130_fd_sc_hd__or2_1 _6920_ (.A(_1864_),
    .B(_3363_),
    .X(_3367_));
 sky130_fd_sc_hd__a21oi_1 _6921_ (.A1(_1864_),
    .A2(_3363_),
    .B1(net976),
    .Y(_3368_));
 sky130_fd_sc_hd__o21ai_1 _6922_ (.A1(\u_s1.u_sync_wbb.m_bl_cnt[0] ),
    .A2(\u_s1.u_sync_wbb.m_bl_cnt[1] ),
    .B1(net976),
    .Y(_3369_));
 sky130_fd_sc_hd__a21oi_1 _6923_ (.A1(\u_s1.u_sync_wbb.m_bl_cnt[0] ),
    .A2(\u_s1.u_sync_wbb.m_bl_cnt[1] ),
    .B1(_3369_),
    .Y(_3370_));
 sky130_fd_sc_hd__a21oi_1 _6924_ (.A1(_3367_),
    .A2(_3368_),
    .B1(_3370_),
    .Y(_3371_));
 sky130_fd_sc_hd__mux2_1 _6925_ (.A0(_3371_),
    .A1(\u_s1.u_sync_wbb.m_bl_cnt[1] ),
    .S(net487),
    .X(_1298_));
 sky130_fd_sc_hd__a21oi_1 _6926_ (.A1(_1864_),
    .A2(_3363_),
    .B1(_1859_),
    .Y(_3372_));
 sky130_fd_sc_hd__a31o_1 _6927_ (.A1(_1859_),
    .A2(_1864_),
    .A3(_3363_),
    .B1(net976),
    .X(_3373_));
 sky130_fd_sc_hd__o21ai_1 _6928_ (.A1(\u_s1.u_sync_wbb.m_bl_cnt[0] ),
    .A2(\u_s1.u_sync_wbb.m_bl_cnt[1] ),
    .B1(\u_s1.u_sync_wbb.m_bl_cnt[2] ),
    .Y(_3374_));
 sky130_fd_sc_hd__or3_1 _6929_ (.A(\u_s1.u_sync_wbb.m_bl_cnt[0] ),
    .B(\u_s1.u_sync_wbb.m_bl_cnt[1] ),
    .C(\u_s1.u_sync_wbb.m_bl_cnt[2] ),
    .X(_3375_));
 sky130_fd_sc_hd__nand2_1 _6930_ (.A(_3374_),
    .B(_3375_),
    .Y(_3376_));
 sky130_fd_sc_hd__o22a_1 _6931_ (.A1(_3372_),
    .A2(_3373_),
    .B1(_3376_),
    .B2(net978),
    .X(_3377_));
 sky130_fd_sc_hd__mux2_1 _6932_ (.A0(_3377_),
    .A1(\u_s1.u_sync_wbb.m_bl_cnt[2] ),
    .S(net487),
    .X(_1299_));
 sky130_fd_sc_hd__a31o_1 _6933_ (.A1(_1859_),
    .A2(_1864_),
    .A3(_3363_),
    .B1(_1861_),
    .X(_3378_));
 sky130_fd_sc_hd__or4b_2 _6934_ (.A(net798),
    .B(_1860_),
    .C(net797),
    .D_N(_3363_),
    .X(_3379_));
 sky130_fd_sc_hd__nand2_1 _6935_ (.A(\u_s1.u_sync_wbb.m_bl_cnt[3] ),
    .B(_3375_),
    .Y(_3380_));
 sky130_fd_sc_hd__or4_2 _6936_ (.A(\u_s1.u_sync_wbb.m_bl_cnt[0] ),
    .B(\u_s1.u_sync_wbb.m_bl_cnt[1] ),
    .C(\u_s1.u_sync_wbb.m_bl_cnt[3] ),
    .D(\u_s1.u_sync_wbb.m_bl_cnt[2] ),
    .X(_3381_));
 sky130_fd_sc_hd__and3_1 _6937_ (.A(net976),
    .B(_3380_),
    .C(_3381_),
    .X(_3382_));
 sky130_fd_sc_hd__a31oi_2 _6938_ (.A1(net978),
    .A2(_3378_),
    .A3(_3379_),
    .B1(_3382_),
    .Y(_3383_));
 sky130_fd_sc_hd__mux2_1 _6939_ (.A0(_3383_),
    .A1(\u_s1.u_sync_wbb.m_bl_cnt[3] ),
    .S(net486),
    .X(_1300_));
 sky130_fd_sc_hd__or2_1 _6940_ (.A(_1865_),
    .B(_1875_),
    .X(_3384_));
 sky130_fd_sc_hd__a21oi_4 _6941_ (.A1(net630),
    .A2(_2001_),
    .B1(_3384_),
    .Y(_3385_));
 sky130_fd_sc_hd__a21o_2 _6942_ (.A1(net630),
    .A2(_2001_),
    .B1(_3384_),
    .X(_3386_));
 sky130_fd_sc_hd__a211o_1 _6943_ (.A1(_1856_),
    .A2(_3379_),
    .B1(_3385_),
    .C1(net976),
    .X(_3387_));
 sky130_fd_sc_hd__a21oi_1 _6944_ (.A1(\u_s1.u_sync_wbb.m_bl_cnt[4] ),
    .A2(_3381_),
    .B1(net978),
    .Y(_3388_));
 sky130_fd_sc_hd__o21a_1 _6945_ (.A1(\u_s1.u_sync_wbb.m_bl_cnt[4] ),
    .A2(_3381_),
    .B1(_3388_),
    .X(_3389_));
 sky130_fd_sc_hd__nor2_1 _6946_ (.A(net486),
    .B(_3389_),
    .Y(_3390_));
 sky130_fd_sc_hd__a22o_1 _6947_ (.A1(\u_s1.u_sync_wbb.m_bl_cnt[4] ),
    .A2(net487),
    .B1(_3387_),
    .B2(_3390_),
    .X(_1301_));
 sky130_fd_sc_hd__xnor2_1 _6948_ (.A(_1869_),
    .B(_3386_),
    .Y(_3391_));
 sky130_fd_sc_hd__nor2_1 _6949_ (.A(net977),
    .B(_3391_),
    .Y(_3392_));
 sky130_fd_sc_hd__or3_4 _6950_ (.A(\u_s1.u_sync_wbb.m_bl_cnt[5] ),
    .B(\u_s1.u_sync_wbb.m_bl_cnt[4] ),
    .C(_3381_),
    .X(_3393_));
 sky130_fd_sc_hd__o21ai_1 _6951_ (.A1(\u_s1.u_sync_wbb.m_bl_cnt[4] ),
    .A2(_3381_),
    .B1(\u_s1.u_sync_wbb.m_bl_cnt[5] ),
    .Y(_3394_));
 sky130_fd_sc_hd__a31o_1 _6952_ (.A1(net976),
    .A2(_3393_),
    .A3(_3394_),
    .B1(net487),
    .X(_3395_));
 sky130_fd_sc_hd__a2bb2o_1 _6953_ (.A1_N(_3392_),
    .A2_N(_3395_),
    .B1(\u_s1.u_sync_wbb.m_bl_cnt[5] ),
    .B2(net487),
    .X(_1302_));
 sky130_fd_sc_hd__o21ai_1 _6954_ (.A1(_1869_),
    .A2(_3386_),
    .B1(_1868_),
    .Y(_3396_));
 sky130_fd_sc_hd__o31a_1 _6955_ (.A1(_1868_),
    .A2(_1869_),
    .A3(_3386_),
    .B1(net978),
    .X(_3397_));
 sky130_fd_sc_hd__or2_1 _6956_ (.A(\u_s1.u_sync_wbb.m_bl_cnt[6] ),
    .B(_3393_),
    .X(_3398_));
 sky130_fd_sc_hd__a21oi_1 _6957_ (.A1(\u_s1.u_sync_wbb.m_bl_cnt[6] ),
    .A2(_3393_),
    .B1(net978),
    .Y(_3399_));
 sky130_fd_sc_hd__a22oi_1 _6958_ (.A1(_3396_),
    .A2(_3397_),
    .B1(_3398_),
    .B2(_3399_),
    .Y(_3400_));
 sky130_fd_sc_hd__mux2_1 _6959_ (.A0(_3400_),
    .A1(\u_s1.u_sync_wbb.m_bl_cnt[6] ),
    .S(net486),
    .X(_1303_));
 sky130_fd_sc_hd__o31ai_1 _6960_ (.A1(_1868_),
    .A2(_1869_),
    .A3(_3386_),
    .B1(_1867_),
    .Y(_3401_));
 sky130_fd_sc_hd__or2_1 _6961_ (.A(_1870_),
    .B(_3386_),
    .X(_3402_));
 sky130_fd_sc_hd__nand2_1 _6962_ (.A(\u_s1.u_sync_wbb.m_bl_cnt[7] ),
    .B(_3398_),
    .Y(_3403_));
 sky130_fd_sc_hd__or3_1 _6963_ (.A(\u_s1.u_sync_wbb.m_bl_cnt[7] ),
    .B(\u_s1.u_sync_wbb.m_bl_cnt[6] ),
    .C(_3393_),
    .X(_3404_));
 sky130_fd_sc_hd__and3_1 _6964_ (.A(net977),
    .B(_3403_),
    .C(_3404_),
    .X(_3405_));
 sky130_fd_sc_hd__a311o_1 _6965_ (.A1(net978),
    .A2(_3401_),
    .A3(_3402_),
    .B1(_3405_),
    .C1(net486),
    .X(_3406_));
 sky130_fd_sc_hd__a21bo_1 _6966_ (.A1(\u_s1.u_sync_wbb.m_bl_cnt[7] ),
    .A2(net486),
    .B1_N(_3406_),
    .X(_1304_));
 sky130_fd_sc_hd__a221o_1 _6967_ (.A1(_1871_),
    .A2(_3385_),
    .B1(_3402_),
    .B2(_1866_),
    .C1(net977),
    .X(_3407_));
 sky130_fd_sc_hd__nor2_1 _6968_ (.A(\u_s1.u_sync_wbb.m_bl_cnt[8] ),
    .B(_3404_),
    .Y(_3408_));
 sky130_fd_sc_hd__or2_1 _6969_ (.A(net978),
    .B(_3408_),
    .X(_3409_));
 sky130_fd_sc_hd__a21oi_1 _6970_ (.A1(\u_s1.u_sync_wbb.m_bl_cnt[8] ),
    .A2(_3404_),
    .B1(_3409_),
    .Y(_3410_));
 sky130_fd_sc_hd__nor2_1 _6971_ (.A(net486),
    .B(_3410_),
    .Y(_3411_));
 sky130_fd_sc_hd__a22o_1 _6972_ (.A1(\u_s1.u_sync_wbb.m_bl_cnt[8] ),
    .A2(net486),
    .B1(_3407_),
    .B2(_3411_),
    .X(_1305_));
 sky130_fd_sc_hd__and2b_1 _6973_ (.A_N(net486),
    .B(_3409_),
    .X(_3412_));
 sky130_fd_sc_hd__or3b_1 _6974_ (.A(_1872_),
    .B(_3386_),
    .C_N(_1873_),
    .X(_3413_));
 sky130_fd_sc_hd__a21o_1 _6975_ (.A1(_1871_),
    .A2(_3385_),
    .B1(_1873_),
    .X(_3414_));
 sky130_fd_sc_hd__a21oi_1 _6976_ (.A1(\u_s1.u_sync_wbb.m_bl_cnt[9] ),
    .A2(_3408_),
    .B1(net978),
    .Y(_3415_));
 sky130_fd_sc_hd__a311o_1 _6977_ (.A1(net978),
    .A2(_3413_),
    .A3(_3414_),
    .B1(_3415_),
    .C1(net486),
    .X(_3416_));
 sky130_fd_sc_hd__o21a_1 _6978_ (.A1(\u_s1.u_sync_wbb.m_bl_cnt[9] ),
    .A2(_3412_),
    .B1(_3416_),
    .X(_1306_));
 sky130_fd_sc_hd__xnor2_1 _6979_ (.A(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[0] ),
    .B(_2423_),
    .Y(_1307_));
 sky130_fd_sc_hd__a21oi_1 _6980_ (.A1(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[0] ),
    .A2(_2424_),
    .B1(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[1] ),
    .Y(_3417_));
 sky130_fd_sc_hd__nor2_1 _6981_ (.A(net496),
    .B(_3417_),
    .Y(_1308_));
 sky130_fd_sc_hd__xor2_1 _6982_ (.A(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[2] ),
    .B(net497),
    .X(_1309_));
 sky130_fd_sc_hd__or2_1 _6983_ (.A(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .B(\u_s0.u_sync_wbb.m_cmd_wr_en ),
    .X(_3418_));
 sky130_fd_sc_hd__and2_1 _6984_ (.A(_3347_),
    .B(_3418_),
    .X(_1310_));
 sky130_fd_sc_hd__and2_1 _6985_ (.A(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .B(_3347_),
    .X(_3419_));
 sky130_fd_sc_hd__nor2_1 _6986_ (.A(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .B(_3347_),
    .Y(_3420_));
 sky130_fd_sc_hd__or2_1 _6987_ (.A(_3419_),
    .B(net747),
    .X(_1311_));
 sky130_fd_sc_hd__xor2_1 _6988_ (.A(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[2] ),
    .B(net965),
    .X(_1312_));
 sky130_fd_sc_hd__and3b_1 _6989_ (.A_N(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .B(\u_s2.u_sync_wbb.m_cmd_wr_en ),
    .C(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .X(_3421_));
 sky130_fd_sc_hd__mux2_1 _6990_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][1] ),
    .A1(net791),
    .S(net942),
    .X(_1313_));
 sky130_fd_sc_hd__mux2_1 _6991_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][2] ),
    .A1(net794),
    .S(net943),
    .X(_1314_));
 sky130_fd_sc_hd__mux2_1 _6992_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][3] ),
    .A1(net792),
    .S(net943),
    .X(_1315_));
 sky130_fd_sc_hd__mux2_1 _6993_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][4] ),
    .A1(net795),
    .S(net942),
    .X(_1316_));
 sky130_fd_sc_hd__mux2_1 _6994_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][5] ),
    .A1(net786),
    .S(net937),
    .X(_1317_));
 sky130_fd_sc_hd__mux2_1 _6995_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][6] ),
    .A1(net788),
    .S(net941),
    .X(_1318_));
 sky130_fd_sc_hd__mux2_1 _6996_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][7] ),
    .A1(net789),
    .S(net937),
    .X(_1319_));
 sky130_fd_sc_hd__mux2_1 _6997_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][8] ),
    .A1(net790),
    .S(net939),
    .X(_1320_));
 sky130_fd_sc_hd__mux2_1 _6998_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][9] ),
    .A1(net785),
    .S(net941),
    .X(_1321_));
 sky130_fd_sc_hd__mux2_1 _6999_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][14] ),
    .A1(net677),
    .S(net942),
    .X(_1322_));
 sky130_fd_sc_hd__mux2_1 _7000_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][15] ),
    .A1(net675),
    .S(net942),
    .X(_1323_));
 sky130_fd_sc_hd__mux2_1 _7001_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][16] ),
    .A1(net673),
    .S(net941),
    .X(_1324_));
 sky130_fd_sc_hd__mux2_1 _7002_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][17] ),
    .A1(net672),
    .S(net938),
    .X(_1325_));
 sky130_fd_sc_hd__mux2_1 _7003_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][18] ),
    .A1(net671),
    .S(net940),
    .X(_1326_));
 sky130_fd_sc_hd__mux2_1 _7004_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][19] ),
    .A1(net670),
    .S(net939),
    .X(_1327_));
 sky130_fd_sc_hd__mux2_1 _7005_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][20] ),
    .A1(net669),
    .S(net942),
    .X(_1328_));
 sky130_fd_sc_hd__mux2_1 _7006_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][21] ),
    .A1(net667),
    .S(net941),
    .X(_1329_));
 sky130_fd_sc_hd__mux2_1 _7007_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][22] ),
    .A1(net666),
    .S(net942),
    .X(_1330_));
 sky130_fd_sc_hd__mux2_1 _7008_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][23] ),
    .A1(net665),
    .S(net939),
    .X(_1331_));
 sky130_fd_sc_hd__mux2_1 _7009_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][24] ),
    .A1(net664),
    .S(net939),
    .X(_1332_));
 sky130_fd_sc_hd__mux2_1 _7010_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][25] ),
    .A1(net663),
    .S(net943),
    .X(_1333_));
 sky130_fd_sc_hd__mux2_1 _7011_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][26] ),
    .A1(_3164_),
    .S(net938),
    .X(_1334_));
 sky130_fd_sc_hd__mux2_1 _7012_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][27] ),
    .A1(net662),
    .S(net941),
    .X(_1335_));
 sky130_fd_sc_hd__mux2_1 _7013_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][28] ),
    .A1(net661),
    .S(net942),
    .X(_1336_));
 sky130_fd_sc_hd__mux2_1 _7014_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][29] ),
    .A1(net660),
    .S(net938),
    .X(_1337_));
 sky130_fd_sc_hd__mux2_1 _7015_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][30] ),
    .A1(net659),
    .S(net939),
    .X(_1338_));
 sky130_fd_sc_hd__mux2_1 _7016_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][31] ),
    .A1(net658),
    .S(net937),
    .X(_1339_));
 sky130_fd_sc_hd__mux2_1 _7017_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][32] ),
    .A1(net657),
    .S(net943),
    .X(_1340_));
 sky130_fd_sc_hd__mux2_1 _7018_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][33] ),
    .A1(net656),
    .S(net941),
    .X(_1341_));
 sky130_fd_sc_hd__mux2_1 _7019_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][34] ),
    .A1(net655),
    .S(net943),
    .X(_1342_));
 sky130_fd_sc_hd__mux2_1 _7020_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][35] ),
    .A1(net654),
    .S(net943),
    .X(_1343_));
 sky130_fd_sc_hd__mux2_1 _7021_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][36] ),
    .A1(net652),
    .S(net942),
    .X(_1344_));
 sky130_fd_sc_hd__mux2_1 _7022_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][37] ),
    .A1(net651),
    .S(net942),
    .X(_1345_));
 sky130_fd_sc_hd__mux2_1 _7023_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][38] ),
    .A1(_3195_),
    .S(net937),
    .X(_1346_));
 sky130_fd_sc_hd__mux2_1 _7024_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][39] ),
    .A1(net650),
    .S(net937),
    .X(_1347_));
 sky130_fd_sc_hd__mux2_1 _7025_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][40] ),
    .A1(net649),
    .S(net939),
    .X(_1348_));
 sky130_fd_sc_hd__mux2_1 _7026_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][41] ),
    .A1(net648),
    .S(net937),
    .X(_1349_));
 sky130_fd_sc_hd__mux2_1 _7027_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][42] ),
    .A1(net647),
    .S(net938),
    .X(_1350_));
 sky130_fd_sc_hd__mux2_1 _7028_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][43] ),
    .A1(net645),
    .S(net939),
    .X(_1351_));
 sky130_fd_sc_hd__mux2_1 _7029_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][44] ),
    .A1(net644),
    .S(net942),
    .X(_1352_));
 sky130_fd_sc_hd__mux2_1 _7030_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][45] ),
    .A1(net643),
    .S(net941),
    .X(_1353_));
 sky130_fd_sc_hd__mux2_1 _7031_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][46] ),
    .A1(net642),
    .S(net938),
    .X(_1354_));
 sky130_fd_sc_hd__mux2_1 _7032_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][47] ),
    .A1(_3216_),
    .S(net937),
    .X(_1355_));
 sky130_fd_sc_hd__mux2_1 _7033_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][48] ),
    .A1(net641),
    .S(net941),
    .X(_1356_));
 sky130_fd_sc_hd__mux2_1 _7034_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][49] ),
    .A1(net640),
    .S(net938),
    .X(_1357_));
 sky130_fd_sc_hd__mux2_1 _7035_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][50] ),
    .A1(net726),
    .S(net939),
    .X(_1358_));
 sky130_fd_sc_hd__mux2_1 _7036_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][53] ),
    .A1(net585),
    .S(net940),
    .X(_1359_));
 sky130_fd_sc_hd__mux2_1 _7037_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][54] ),
    .A1(net639),
    .S(net941),
    .X(_1360_));
 sky130_fd_sc_hd__mux2_1 _7038_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][55] ),
    .A1(net638),
    .S(net939),
    .X(_1361_));
 sky130_fd_sc_hd__mux2_1 _7039_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][56] ),
    .A1(net637),
    .S(net939),
    .X(_1362_));
 sky130_fd_sc_hd__mux2_1 _7040_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][57] ),
    .A1(net636),
    .S(net940),
    .X(_1363_));
 sky130_fd_sc_hd__mux2_1 _7041_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][58] ),
    .A1(net635),
    .S(net937),
    .X(_1364_));
 sky130_fd_sc_hd__mux2_1 _7042_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][59] ),
    .A1(net633),
    .S(net941),
    .X(_1365_));
 sky130_fd_sc_hd__mux2_1 _7043_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][60] ),
    .A1(net632),
    .S(net937),
    .X(_1366_));
 sky130_fd_sc_hd__mux2_1 _7044_ (.A0(\u_s2.u_sync_wbb.u_cmd_if.mem[1][61] ),
    .A1(net631),
    .S(net937),
    .X(_1367_));
 sky130_fd_sc_hd__or3_1 _7045_ (.A(net727),
    .B(net333),
    .C(net332),
    .X(_3422_));
 sky130_fd_sc_hd__or4_1 _7046_ (.A(net340),
    .B(net731),
    .C(net730),
    .D(net335),
    .X(_3423_));
 sky130_fd_sc_hd__or4_1 _7047_ (.A(net729),
    .B(net728),
    .C(_3422_),
    .D(_3423_),
    .X(_3424_));
 sky130_fd_sc_hd__a32o_1 _7048_ (.A1(_1705_),
    .A2(net342),
    .A3(_3424_),
    .B1(_1706_),
    .B2(\u_s0.u_sync_wbb.wbs_burst ),
    .X(_1368_));
 sky130_fd_sc_hd__xor2_1 _7049_ (.A(net1337),
    .B(net567),
    .X(_1369_));
 sky130_fd_sc_hd__and3_1 _7050_ (.A(net1339),
    .B(net1329),
    .C(net570),
    .X(_3425_));
 sky130_fd_sc_hd__a21oi_1 _7051_ (.A1(net1340),
    .A2(net569),
    .B1(net1330),
    .Y(_3426_));
 sky130_fd_sc_hd__nor2_1 _7052_ (.A(_3425_),
    .B(_3426_),
    .Y(_1370_));
 sky130_fd_sc_hd__xor2_1 _7053_ (.A(\u_s0.u_sync_wbb.u_cmd_if.rd_ptr[2] ),
    .B(_3425_),
    .X(_1371_));
 sky130_fd_sc_hd__xor2_1 _7054_ (.A(net1320),
    .B(\u_s0.u_sync_wbb.m_resp_rd_en ),
    .X(_1372_));
 sky130_fd_sc_hd__a21oi_1 _7055_ (.A1(net1320),
    .A2(\u_s0.u_sync_wbb.m_resp_rd_en ),
    .B1(net1315),
    .Y(_3427_));
 sky130_fd_sc_hd__and3_1 _7056_ (.A(net1315),
    .B(net1320),
    .C(\u_s0.u_sync_wbb.m_resp_rd_en ),
    .X(_3428_));
 sky130_fd_sc_hd__nor2_1 _7057_ (.A(_3427_),
    .B(_3428_),
    .Y(_1373_));
 sky130_fd_sc_hd__xor2_1 _7058_ (.A(\u_s0.u_sync_wbb.u_resp_if.rd_ptr[2] ),
    .B(_3428_),
    .X(_1374_));
 sky130_fd_sc_hd__a22o_1 _7059_ (.A1(\u_reg.reg_7[0] ),
    .A2(net603),
    .B1(net593),
    .B2(\u_reg.reg_3[0] ),
    .X(_3429_));
 sky130_fd_sc_hd__a221o_1 _7060_ (.A1(\u_reg.reg_4[0] ),
    .A2(net598),
    .B1(net545),
    .B2(\u_dcg_s0.cfg_mode[0] ),
    .C1(_3429_),
    .X(_3430_));
 sky130_fd_sc_hd__and2_4 _7061_ (.A(_2662_),
    .B(_2779_),
    .X(_3431_));
 sky130_fd_sc_hd__nand2_4 _7062_ (.A(_2662_),
    .B(_2779_),
    .Y(_3432_));
 sky130_fd_sc_hd__a22o_1 _7063_ (.A1(\u_reg.reg_6[0] ),
    .A2(net610),
    .B1(net587),
    .B2(\u_reg.reg_2[0] ),
    .X(_3433_));
 sky130_fd_sc_hd__a21o_1 _7064_ (.A1(\u_reg.reg_5[0] ),
    .A2(net621),
    .B1(_3433_),
    .X(_3434_));
 sky130_fd_sc_hd__or3_1 _7065_ (.A(_3430_),
    .B(_3431_),
    .C(_3434_),
    .X(_3435_));
 sky130_fd_sc_hd__a21oi_2 _7066_ (.A1(_1686_),
    .A2(_3431_),
    .B1(net626),
    .Y(_3436_));
 sky130_fd_sc_hd__a22o_1 _7067_ (.A1(\u_reg.reg_rdata[0] ),
    .A2(net626),
    .B1(_3435_),
    .B2(_3436_),
    .X(_1375_));
 sky130_fd_sc_hd__a22o_1 _7068_ (.A1(\u_reg.reg_7[1] ),
    .A2(net603),
    .B1(net593),
    .B2(\u_reg.reg_3[1] ),
    .X(_3437_));
 sky130_fd_sc_hd__a221o_1 _7069_ (.A1(\u_reg.reg_4[1] ),
    .A2(net598),
    .B1(net545),
    .B2(\u_dcg_s0.cfg_mode[1] ),
    .C1(_3437_),
    .X(_3438_));
 sky130_fd_sc_hd__a22o_1 _7070_ (.A1(\u_reg.reg_6[1] ),
    .A2(net610),
    .B1(net587),
    .B2(\u_reg.reg_2[1] ),
    .X(_3439_));
 sky130_fd_sc_hd__a21o_1 _7071_ (.A1(\u_reg.reg_5[1] ),
    .A2(net621),
    .B1(_3439_),
    .X(_3440_));
 sky130_fd_sc_hd__or3_1 _7072_ (.A(_3431_),
    .B(_3438_),
    .C(_3440_),
    .X(_3441_));
 sky130_fd_sc_hd__a21oi_1 _7073_ (.A1(_1690_),
    .A2(_3431_),
    .B1(net626),
    .Y(_3442_));
 sky130_fd_sc_hd__a22o_1 _7074_ (.A1(\u_reg.reg_rdata[1] ),
    .A2(net626),
    .B1(_3441_),
    .B2(_3442_),
    .X(_1376_));
 sky130_fd_sc_hd__or2_1 _7075_ (.A(\u_dcg_s1.cfg_mode[0] ),
    .B(_2662_),
    .X(_3443_));
 sky130_fd_sc_hd__a22o_1 _7076_ (.A1(\u_reg.reg_7[2] ),
    .A2(net603),
    .B1(net587),
    .B2(\u_reg.reg_2[2] ),
    .X(_3444_));
 sky130_fd_sc_hd__a21o_1 _7077_ (.A1(\u_reg.reg_5[2] ),
    .A2(net621),
    .B1(_3444_),
    .X(_3445_));
 sky130_fd_sc_hd__a22o_1 _7078_ (.A1(\u_reg.reg_3[2] ),
    .A2(net593),
    .B1(_2779_),
    .B2(_3443_),
    .X(_3446_));
 sky130_fd_sc_hd__a221o_1 _7079_ (.A1(\u_reg.reg_6[2] ),
    .A2(net610),
    .B1(net598),
    .B2(\u_reg.reg_4[2] ),
    .C1(_3446_),
    .X(_3447_));
 sky130_fd_sc_hd__o221a_1 _7080_ (.A1(m2_wbd_stb_i),
    .A2(net519),
    .B1(_3445_),
    .B2(_3447_),
    .C1(net575),
    .X(_3448_));
 sky130_fd_sc_hd__a21o_1 _7081_ (.A1(\u_reg.reg_rdata[2] ),
    .A2(net626),
    .B1(_3448_),
    .X(_1377_));
 sky130_fd_sc_hd__or2_1 _7082_ (.A(\u_dcg_s1.cfg_mode[1] ),
    .B(_2662_),
    .X(_3449_));
 sky130_fd_sc_hd__a22o_1 _7083_ (.A1(\u_reg.reg_7[3] ),
    .A2(net603),
    .B1(net587),
    .B2(\u_reg.reg_2[3] ),
    .X(_3450_));
 sky130_fd_sc_hd__a21o_1 _7084_ (.A1(\u_reg.reg_6[3] ),
    .A2(net610),
    .B1(_3450_),
    .X(_3451_));
 sky130_fd_sc_hd__a22o_1 _7085_ (.A1(\u_reg.reg_3[3] ),
    .A2(net593),
    .B1(_2779_),
    .B2(_3449_),
    .X(_3452_));
 sky130_fd_sc_hd__a221o_1 _7086_ (.A1(\u_reg.reg_5[3] ),
    .A2(net621),
    .B1(net598),
    .B2(\u_reg.reg_4[3] ),
    .C1(_3452_),
    .X(_3453_));
 sky130_fd_sc_hd__o221a_1 _7087_ (.A1(m3_wbd_stb_i),
    .A2(net519),
    .B1(_3451_),
    .B2(_3453_),
    .C1(net575),
    .X(_3454_));
 sky130_fd_sc_hd__a21o_1 _7088_ (.A1(\u_reg.reg_rdata[3] ),
    .A2(net626),
    .B1(_3454_),
    .X(_1378_));
 sky130_fd_sc_hd__a22o_1 _7089_ (.A1(\u_reg.reg_6[4] ),
    .A2(net610),
    .B1(net546),
    .B2(\u_dcg_s2.cfg_mode[0] ),
    .X(_3455_));
 sky130_fd_sc_hd__a22o_1 _7090_ (.A1(\u_reg.reg_7[4] ),
    .A2(net604),
    .B1(net594),
    .B2(\u_reg.reg_3[4] ),
    .X(_3456_));
 sky130_fd_sc_hd__a221o_1 _7091_ (.A1(\u_reg.reg_4[4] ),
    .A2(net599),
    .B1(net586),
    .B2(\u_reg.reg_2[4] ),
    .C1(_3456_),
    .X(_3457_));
 sky130_fd_sc_hd__a211o_1 _7092_ (.A1(\u_reg.reg_5[4] ),
    .A2(net622),
    .B1(_3455_),
    .C1(_3457_),
    .X(_3458_));
 sky130_fd_sc_hd__mux2_1 _7093_ (.A0(\u_reg.reg_rdata[4] ),
    .A1(_3458_),
    .S(net579),
    .X(_1379_));
 sky130_fd_sc_hd__a22o_1 _7094_ (.A1(\u_reg.reg_6[5] ),
    .A2(net616),
    .B1(net546),
    .B2(\u_dcg_s2.cfg_mode[1] ),
    .X(_3459_));
 sky130_fd_sc_hd__a22o_1 _7095_ (.A1(\u_reg.reg_7[5] ),
    .A2(net604),
    .B1(net594),
    .B2(\u_reg.reg_3[5] ),
    .X(_3460_));
 sky130_fd_sc_hd__a221o_1 _7096_ (.A1(\u_reg.reg_4[5] ),
    .A2(net599),
    .B1(net587),
    .B2(\u_reg.reg_2[5] ),
    .C1(_3460_),
    .X(_3461_));
 sky130_fd_sc_hd__a211o_1 _7097_ (.A1(\u_reg.reg_5[5] ),
    .A2(net622),
    .B1(_3459_),
    .C1(_3461_),
    .X(_3462_));
 sky130_fd_sc_hd__mux2_1 _7098_ (.A0(\u_reg.reg_rdata[5] ),
    .A1(_3462_),
    .S(net576),
    .X(_1380_));
 sky130_fd_sc_hd__a22o_1 _7099_ (.A1(\u_reg.reg_6[6] ),
    .A2(net610),
    .B1(net545),
    .B2(\u_dcg_peri.cfg_mode[0] ),
    .X(_3463_));
 sky130_fd_sc_hd__a22o_1 _7100_ (.A1(\u_reg.reg_4[6] ),
    .A2(net598),
    .B1(net586),
    .B2(\u_reg.reg_2[6] ),
    .X(_3464_));
 sky130_fd_sc_hd__a221o_1 _7101_ (.A1(\u_reg.reg_7[6] ),
    .A2(net603),
    .B1(net593),
    .B2(\u_reg.reg_3[6] ),
    .C1(_3464_),
    .X(_3465_));
 sky130_fd_sc_hd__a211o_2 _7102_ (.A1(\u_reg.reg_5[6] ),
    .A2(net622),
    .B1(_3463_),
    .C1(_3465_),
    .X(_3466_));
 sky130_fd_sc_hd__mux2_1 _7103_ (.A0(\u_reg.reg_rdata[6] ),
    .A1(_3466_),
    .S(net575),
    .X(_1381_));
 sky130_fd_sc_hd__a22o_1 _7104_ (.A1(\u_reg.reg_6[7] ),
    .A2(net610),
    .B1(net545),
    .B2(\u_dcg_peri.cfg_mode[1] ),
    .X(_3467_));
 sky130_fd_sc_hd__a22o_1 _7105_ (.A1(\u_reg.reg_4[7] ),
    .A2(net598),
    .B1(net586),
    .B2(\u_reg.reg_2[7] ),
    .X(_3468_));
 sky130_fd_sc_hd__a221o_2 _7106_ (.A1(\u_reg.reg_7[7] ),
    .A2(net603),
    .B1(net594),
    .B2(\u_reg.reg_3[7] ),
    .C1(_3468_),
    .X(_3469_));
 sky130_fd_sc_hd__a211o_1 _7107_ (.A1(\u_reg.reg_5[7] ),
    .A2(net622),
    .B1(_3467_),
    .C1(_3469_),
    .X(_3470_));
 sky130_fd_sc_hd__mux2_1 _7108_ (.A0(\u_reg.reg_rdata[7] ),
    .A1(_3470_),
    .S(net575),
    .X(_1382_));
 sky130_fd_sc_hd__a22o_1 _7109_ (.A1(\u_reg.reg_7[8] ),
    .A2(net604),
    .B1(net588),
    .B2(\u_reg.reg_2[8] ),
    .X(_3471_));
 sky130_fd_sc_hd__or2_1 _7110_ (.A(\u_dcg_riscv.cfg_mode[0] ),
    .B(_2662_),
    .X(_3472_));
 sky130_fd_sc_hd__a21o_1 _7111_ (.A1(\u_reg.reg_6[8] ),
    .A2(net611),
    .B1(_3471_),
    .X(_3473_));
 sky130_fd_sc_hd__a22o_1 _7112_ (.A1(\u_reg.reg_3[8] ),
    .A2(net594),
    .B1(_2779_),
    .B2(_3472_),
    .X(_3474_));
 sky130_fd_sc_hd__a221o_1 _7113_ (.A1(\u_reg.reg_5[8] ),
    .A2(net622),
    .B1(net599),
    .B2(\u_reg.reg_4[8] ),
    .C1(_3474_),
    .X(_3475_));
 sky130_fd_sc_hd__o221a_2 _7114_ (.A1(\u_dsync.out_data[0] ),
    .A2(net518),
    .B1(_3473_),
    .B2(_3475_),
    .C1(net576),
    .X(_3476_));
 sky130_fd_sc_hd__a21o_1 _7115_ (.A1(\u_reg.reg_rdata[8] ),
    .A2(net626),
    .B1(_3476_),
    .X(_1383_));
 sky130_fd_sc_hd__a22o_1 _7116_ (.A1(\u_reg.reg_7[9] ),
    .A2(net605),
    .B1(net595),
    .B2(\u_reg.reg_3[9] ),
    .X(_3477_));
 sky130_fd_sc_hd__a221o_2 _7117_ (.A1(\u_reg.reg_4[9] ),
    .A2(net601),
    .B1(net547),
    .B2(\u_dcg_riscv.cfg_mode[1] ),
    .C1(_3477_),
    .X(_3478_));
 sky130_fd_sc_hd__a22o_1 _7118_ (.A1(\u_reg.reg_6[9] ),
    .A2(net616),
    .B1(net586),
    .B2(\u_reg.reg_2[9] ),
    .X(_3479_));
 sky130_fd_sc_hd__a21o_1 _7119_ (.A1(\u_reg.reg_5[9] ),
    .A2(net622),
    .B1(_3479_),
    .X(_3480_));
 sky130_fd_sc_hd__or3_2 _7120_ (.A(_3431_),
    .B(net485),
    .C(_3480_),
    .X(_3481_));
 sky130_fd_sc_hd__o21a_1 _7121_ (.A1(\u_dsync.out_data[1] ),
    .A2(net519),
    .B1(net579),
    .X(_3482_));
 sky130_fd_sc_hd__a22o_1 _7122_ (.A1(\u_reg.reg_rdata[9] ),
    .A2(net626),
    .B1(_3481_),
    .B2(_3482_),
    .X(_1384_));
 sky130_fd_sc_hd__a22o_1 _7123_ (.A1(\u_reg.reg_7[10] ),
    .A2(net608),
    .B1(net594),
    .B2(\u_reg.reg_3[10] ),
    .X(_3483_));
 sky130_fd_sc_hd__a221o_1 _7124_ (.A1(\u_reg.reg_4[10] ),
    .A2(net599),
    .B1(net546),
    .B2(\u_reg.cfg_dcg_ctrl[10] ),
    .C1(_3483_),
    .X(_3484_));
 sky130_fd_sc_hd__a22o_1 _7125_ (.A1(\u_reg.reg_6[10] ),
    .A2(net611),
    .B1(net586),
    .B2(\u_reg.reg_2[10] ),
    .X(_3485_));
 sky130_fd_sc_hd__a211o_1 _7126_ (.A1(\u_reg.reg_5[10] ),
    .A2(net624),
    .B1(_3431_),
    .C1(_3485_),
    .X(_3486_));
 sky130_fd_sc_hd__o22a_1 _7127_ (.A1(\u_dsync.out_data[2] ),
    .A2(net518),
    .B1(_3484_),
    .B2(_3486_),
    .X(_3487_));
 sky130_fd_sc_hd__mux2_1 _7128_ (.A0(\u_reg.reg_rdata[10] ),
    .A1(_3487_),
    .S(net574),
    .X(_1385_));
 sky130_fd_sc_hd__a22o_1 _7129_ (.A1(\u_reg.reg_7[11] ),
    .A2(net605),
    .B1(net595),
    .B2(\u_reg.reg_3[11] ),
    .X(_3488_));
 sky130_fd_sc_hd__a221o_1 _7130_ (.A1(\u_reg.reg_4[11] ),
    .A2(net601),
    .B1(net547),
    .B2(\u_reg.cfg_dcg_ctrl[11] ),
    .C1(_3488_),
    .X(_3489_));
 sky130_fd_sc_hd__a22o_1 _7131_ (.A1(\u_reg.reg_6[11] ),
    .A2(net615),
    .B1(net588),
    .B2(\u_reg.reg_2[11] ),
    .X(_3490_));
 sky130_fd_sc_hd__a21o_1 _7132_ (.A1(\u_reg.reg_5[11] ),
    .A2(net623),
    .B1(_3490_),
    .X(_3491_));
 sky130_fd_sc_hd__or3_4 _7133_ (.A(_3431_),
    .B(_3489_),
    .C(_3491_),
    .X(_3492_));
 sky130_fd_sc_hd__o21a_1 _7134_ (.A1(\u_dsync.out_data[3] ),
    .A2(net519),
    .B1(net579),
    .X(_3493_));
 sky130_fd_sc_hd__a22o_1 _7135_ (.A1(\u_reg.reg_rdata[11] ),
    .A2(net626),
    .B1(_3492_),
    .B2(_3493_),
    .X(_1386_));
 sky130_fd_sc_hd__a22o_1 _7136_ (.A1(\u_reg.reg_7[12] ),
    .A2(net604),
    .B1(net596),
    .B2(\u_reg.reg_3[12] ),
    .X(_3494_));
 sky130_fd_sc_hd__a221o_1 _7137_ (.A1(\u_reg.reg_4[12] ),
    .A2(net600),
    .B1(net548),
    .B2(\u_reg.cfg_dcg_ctrl[12] ),
    .C1(_3494_),
    .X(_3495_));
 sky130_fd_sc_hd__a22o_1 _7138_ (.A1(\u_reg.reg_6[12] ),
    .A2(net613),
    .B1(net588),
    .B2(\u_reg.reg_2[12] ),
    .X(_3496_));
 sky130_fd_sc_hd__a211o_1 _7139_ (.A1(\u_reg.reg_5[12] ),
    .A2(net624),
    .B1(_3431_),
    .C1(_3496_),
    .X(_3497_));
 sky130_fd_sc_hd__o22a_1 _7140_ (.A1(\u_dsync.out_data[4] ),
    .A2(_3432_),
    .B1(_3495_),
    .B2(_3497_),
    .X(_3498_));
 sky130_fd_sc_hd__mux2_1 _7141_ (.A0(\u_reg.reg_rdata[12] ),
    .A1(_3498_),
    .S(net577),
    .X(_1387_));
 sky130_fd_sc_hd__a22o_1 _7142_ (.A1(\u_reg.reg_7[13] ),
    .A2(net604),
    .B1(net596),
    .B2(\u_reg.reg_3[13] ),
    .X(_3499_));
 sky130_fd_sc_hd__a221o_1 _7143_ (.A1(\u_reg.reg_4[13] ),
    .A2(net600),
    .B1(net548),
    .B2(\u_reg.cfg_dcg_ctrl[13] ),
    .C1(_3499_),
    .X(_3500_));
 sky130_fd_sc_hd__a22o_1 _7144_ (.A1(\u_reg.reg_6[13] ),
    .A2(net611),
    .B1(net588),
    .B2(\u_reg.reg_2[13] ),
    .X(_3501_));
 sky130_fd_sc_hd__a21o_1 _7145_ (.A1(\u_reg.reg_5[13] ),
    .A2(net623),
    .B1(_3501_),
    .X(_3502_));
 sky130_fd_sc_hd__or3_1 _7146_ (.A(_3431_),
    .B(_3500_),
    .C(_3502_),
    .X(_3503_));
 sky130_fd_sc_hd__o21a_1 _7147_ (.A1(\u_dsync.out_data[5] ),
    .A2(net518),
    .B1(net577),
    .X(_3504_));
 sky130_fd_sc_hd__a22o_1 _7148_ (.A1(\u_reg.reg_rdata[13] ),
    .A2(net627),
    .B1(_3503_),
    .B2(_3504_),
    .X(_1388_));
 sky130_fd_sc_hd__nor2_1 _7149_ (.A(\u_dsync.out_data[6] ),
    .B(net518),
    .Y(_3505_));
 sky130_fd_sc_hd__a22o_1 _7150_ (.A1(\u_reg.reg_7[14] ),
    .A2(net605),
    .B1(net595),
    .B2(\u_reg.reg_3[14] ),
    .X(_3506_));
 sky130_fd_sc_hd__a221oi_4 _7151_ (.A1(\u_reg.reg_4[14] ),
    .A2(net601),
    .B1(net547),
    .B2(\u_reg.cfg_dcg_ctrl[14] ),
    .C1(_3506_),
    .Y(_3507_));
 sky130_fd_sc_hd__a22o_1 _7152_ (.A1(\u_reg.reg_6[14] ),
    .A2(net611),
    .B1(net588),
    .B2(\u_reg.reg_2[14] ),
    .X(_3508_));
 sky130_fd_sc_hd__a21oi_1 _7153_ (.A1(\u_reg.reg_5[14] ),
    .A2(net623),
    .B1(_3508_),
    .Y(_3509_));
 sky130_fd_sc_hd__a31o_1 _7154_ (.A1(net518),
    .A2(_3507_),
    .A3(_3509_),
    .B1(net627),
    .X(_3510_));
 sky130_fd_sc_hd__a2bb2o_1 _7155_ (.A1_N(_3505_),
    .A2_N(_3510_),
    .B1(\u_reg.reg_rdata[14] ),
    .B2(net627),
    .X(_1389_));
 sky130_fd_sc_hd__a22o_1 _7156_ (.A1(\u_reg.reg_7[15] ),
    .A2(net605),
    .B1(net595),
    .B2(\u_reg.reg_3[15] ),
    .X(_3511_));
 sky130_fd_sc_hd__a221o_2 _7157_ (.A1(\u_reg.reg_4[15] ),
    .A2(net601),
    .B1(net547),
    .B2(\u_reg.cfg_dcg_ctrl[15] ),
    .C1(_3511_),
    .X(_3512_));
 sky130_fd_sc_hd__a22o_1 _7158_ (.A1(\u_reg.reg_6[15] ),
    .A2(net611),
    .B1(net588),
    .B2(\u_reg.reg_2[15] ),
    .X(_3513_));
 sky130_fd_sc_hd__a21o_1 _7159_ (.A1(\u_reg.reg_5[15] ),
    .A2(net624),
    .B1(_3513_),
    .X(_3514_));
 sky130_fd_sc_hd__or3_1 _7160_ (.A(_3431_),
    .B(_3512_),
    .C(_3514_),
    .X(_3515_));
 sky130_fd_sc_hd__o21a_1 _7161_ (.A1(\u_dsync.out_data[7] ),
    .A2(net518),
    .B1(net577),
    .X(_3516_));
 sky130_fd_sc_hd__a22o_1 _7162_ (.A1(\u_reg.reg_rdata[15] ),
    .A2(net627),
    .B1(_3515_),
    .B2(_3516_),
    .X(_1390_));
 sky130_fd_sc_hd__a22o_1 _7163_ (.A1(\u_reg.reg_6[16] ),
    .A2(net613),
    .B1(net547),
    .B2(net1824),
    .X(_3517_));
 sky130_fd_sc_hd__a22o_1 _7164_ (.A1(\u_reg.reg_4[16] ),
    .A2(net600),
    .B1(net590),
    .B2(\u_reg.reg_2[16] ),
    .X(_3518_));
 sky130_fd_sc_hd__a221o_1 _7165_ (.A1(\u_reg.reg_7[16] ),
    .A2(net605),
    .B1(net595),
    .B2(\u_reg.reg_3[16] ),
    .C1(_3518_),
    .X(_3519_));
 sky130_fd_sc_hd__a211o_1 _7166_ (.A1(\u_reg.reg_5[16] ),
    .A2(net623),
    .B1(_3517_),
    .C1(_3519_),
    .X(_3520_));
 sky130_fd_sc_hd__mux2_1 _7167_ (.A0(\u_reg.reg_rdata[16] ),
    .A1(net1825),
    .S(net576),
    .X(_1391_));
 sky130_fd_sc_hd__a22o_1 _7168_ (.A1(\u_reg.reg_6[17] ),
    .A2(net613),
    .B1(net547),
    .B2(\u_reg.cfg_dcg_ctrl[17] ),
    .X(_3521_));
 sky130_fd_sc_hd__a22o_1 _7169_ (.A1(\u_reg.reg_7[17] ),
    .A2(net605),
    .B1(net595),
    .B2(\u_reg.reg_3[17] ),
    .X(_3522_));
 sky130_fd_sc_hd__a221o_2 _7170_ (.A1(\u_reg.reg_4[17] ),
    .A2(net601),
    .B1(net590),
    .B2(\u_reg.reg_2[17] ),
    .C1(_3522_),
    .X(_3523_));
 sky130_fd_sc_hd__a211o_1 _7171_ (.A1(net1793),
    .A2(net623),
    .B1(_3521_),
    .C1(_3523_),
    .X(_3524_));
 sky130_fd_sc_hd__mux2_1 _7172_ (.A0(\u_reg.reg_rdata[17] ),
    .A1(net1794),
    .S(net577),
    .X(_1392_));
 sky130_fd_sc_hd__a22o_1 _7173_ (.A1(\u_reg.reg_6[18] ),
    .A2(net610),
    .B1(net545),
    .B2(\u_reg.cfg_dcg_ctrl[18] ),
    .X(_3525_));
 sky130_fd_sc_hd__a22o_1 _7174_ (.A1(\u_reg.reg_4[18] ),
    .A2(net599),
    .B1(net586),
    .B2(\u_reg.reg_2[18] ),
    .X(_3526_));
 sky130_fd_sc_hd__a221o_4 _7175_ (.A1(\u_reg.reg_7[18] ),
    .A2(net603),
    .B1(net593),
    .B2(\u_reg.reg_3[18] ),
    .C1(_3526_),
    .X(_3527_));
 sky130_fd_sc_hd__a211o_1 _7176_ (.A1(\u_reg.reg_5[18] ),
    .A2(net621),
    .B1(_3525_),
    .C1(_3527_),
    .X(_3528_));
 sky130_fd_sc_hd__mux2_1 _7177_ (.A0(\u_reg.reg_rdata[18] ),
    .A1(_3528_),
    .S(net575),
    .X(_1393_));
 sky130_fd_sc_hd__a22o_1 _7178_ (.A1(\u_reg.reg_6[19] ),
    .A2(net616),
    .B1(net545),
    .B2(\u_reg.cfg_dcg_ctrl[19] ),
    .X(_3529_));
 sky130_fd_sc_hd__a22o_1 _7179_ (.A1(\u_reg.reg_7[19] ),
    .A2(net608),
    .B1(net593),
    .B2(\u_reg.reg_3[19] ),
    .X(_3530_));
 sky130_fd_sc_hd__a221o_1 _7180_ (.A1(\u_reg.reg_4[19] ),
    .A2(net598),
    .B1(net586),
    .B2(\u_reg.reg_2[19] ),
    .C1(_3530_),
    .X(_3531_));
 sky130_fd_sc_hd__a211o_2 _7181_ (.A1(\u_reg.reg_5[19] ),
    .A2(net621),
    .B1(_3529_),
    .C1(_3531_),
    .X(_3532_));
 sky130_fd_sc_hd__mux2_1 _7182_ (.A0(\u_reg.reg_rdata[19] ),
    .A1(_3532_),
    .S(net575),
    .X(_1394_));
 sky130_fd_sc_hd__a22o_1 _7183_ (.A1(\u_reg.reg_7[20] ),
    .A2(net604),
    .B1(net596),
    .B2(\u_reg.reg_3[20] ),
    .X(_3533_));
 sky130_fd_sc_hd__a22o_1 _7184_ (.A1(\u_reg.reg_6[20] ),
    .A2(net613),
    .B1(net548),
    .B2(\u_reg.cfg_dcg_ctrl[20] ),
    .X(_3534_));
 sky130_fd_sc_hd__a221o_1 _7185_ (.A1(\u_reg.reg_4[20] ),
    .A2(net600),
    .B1(net591),
    .B2(\u_reg.reg_2[20] ),
    .C1(_3533_),
    .X(_3535_));
 sky130_fd_sc_hd__a211o_1 _7186_ (.A1(\u_reg.reg_5[20] ),
    .A2(net623),
    .B1(_3534_),
    .C1(_3535_),
    .X(_3536_));
 sky130_fd_sc_hd__mux2_1 _7187_ (.A0(\u_reg.reg_rdata[20] ),
    .A1(_3536_),
    .S(net577),
    .X(_1395_));
 sky130_fd_sc_hd__a22o_1 _7188_ (.A1(\u_reg.reg_7[21] ),
    .A2(net604),
    .B1(net596),
    .B2(\u_reg.reg_3[21] ),
    .X(_3537_));
 sky130_fd_sc_hd__a22o_1 _7189_ (.A1(\u_reg.reg_6[21] ),
    .A2(net611),
    .B1(net548),
    .B2(\u_reg.cfg_dcg_ctrl[21] ),
    .X(_3538_));
 sky130_fd_sc_hd__a221o_1 _7190_ (.A1(\u_reg.reg_4[21] ),
    .A2(net600),
    .B1(net588),
    .B2(\u_reg.reg_2[21] ),
    .C1(_3537_),
    .X(_3539_));
 sky130_fd_sc_hd__a211o_1 _7191_ (.A1(\u_reg.reg_5[21] ),
    .A2(net624),
    .B1(_3538_),
    .C1(_3539_),
    .X(_3540_));
 sky130_fd_sc_hd__mux2_1 _7192_ (.A0(\u_reg.reg_rdata[21] ),
    .A1(_3540_),
    .S(net577),
    .X(_1396_));
 sky130_fd_sc_hd__a22o_1 _7193_ (.A1(\u_reg.reg_4[22] ),
    .A2(net599),
    .B1(net586),
    .B2(\u_reg.reg_2[22] ),
    .X(_3541_));
 sky130_fd_sc_hd__a22o_1 _7194_ (.A1(\u_reg.reg_6[22] ),
    .A2(net610),
    .B1(net545),
    .B2(\u_reg.cfg_dcg_ctrl[22] ),
    .X(_3542_));
 sky130_fd_sc_hd__a221o_2 _7195_ (.A1(\u_reg.reg_7[22] ),
    .A2(net603),
    .B1(net593),
    .B2(\u_reg.reg_3[22] ),
    .C1(_3541_),
    .X(_3543_));
 sky130_fd_sc_hd__a211o_1 _7196_ (.A1(\u_reg.reg_5[22] ),
    .A2(net621),
    .B1(_3542_),
    .C1(_3543_),
    .X(_3544_));
 sky130_fd_sc_hd__mux2_1 _7197_ (.A0(net1290),
    .A1(_3544_),
    .S(net575),
    .X(_1397_));
 sky130_fd_sc_hd__and2_1 _7198_ (.A(\u_reg.reg_5[23] ),
    .B(net621),
    .X(_3545_));
 sky130_fd_sc_hd__a221o_1 _7199_ (.A1(\u_reg.reg_4[23] ),
    .A2(net598),
    .B1(net545),
    .B2(\u_reg.cfg_dcg_ctrl[23] ),
    .C1(_3545_),
    .X(_3546_));
 sky130_fd_sc_hd__a22o_1 _7200_ (.A1(\u_reg.reg_7[23] ),
    .A2(net604),
    .B1(net588),
    .B2(\u_reg.reg_2[23] ),
    .X(_3547_));
 sky130_fd_sc_hd__a221o_4 _7201_ (.A1(\u_reg.reg_6[23] ),
    .A2(net611),
    .B1(net594),
    .B2(\u_reg.reg_3[23] ),
    .C1(_3547_),
    .X(_3548_));
 sky130_fd_sc_hd__or3_4 _7202_ (.A(net626),
    .B(_3546_),
    .C(_3548_),
    .X(_3549_));
 sky130_fd_sc_hd__o21a_1 _7203_ (.A1(\u_reg.reg_rdata[23] ),
    .A2(net575),
    .B1(_3549_),
    .X(_1398_));
 sky130_fd_sc_hd__a22o_1 _7204_ (.A1(\u_reg.reg_6[24] ),
    .A2(net613),
    .B1(net547),
    .B2(\u_reg.cfg_dcg_ctrl[24] ),
    .X(_3550_));
 sky130_fd_sc_hd__a22o_1 _7205_ (.A1(\u_reg.reg_7[24] ),
    .A2(net605),
    .B1(net595),
    .B2(\u_reg.reg_3[24] ),
    .X(_3551_));
 sky130_fd_sc_hd__a221o_1 _7206_ (.A1(\u_reg.reg_4[24] ),
    .A2(net601),
    .B1(net590),
    .B2(\u_reg.reg_2[24] ),
    .C1(_3551_),
    .X(_3552_));
 sky130_fd_sc_hd__a211o_1 _7207_ (.A1(\u_reg.reg_5[24] ),
    .A2(net623),
    .B1(_3550_),
    .C1(_3552_),
    .X(_3553_));
 sky130_fd_sc_hd__mux2_1 _7208_ (.A0(\u_reg.reg_rdata[24] ),
    .A1(net480),
    .S(net576),
    .X(_1399_));
 sky130_fd_sc_hd__a22o_1 _7209_ (.A1(\u_reg.reg_4[25] ),
    .A2(net601),
    .B1(net590),
    .B2(\u_reg.reg_2[25] ),
    .X(_3554_));
 sky130_fd_sc_hd__a22o_1 _7210_ (.A1(\u_reg.reg_6[25] ),
    .A2(net613),
    .B1(net547),
    .B2(\u_reg.cfg_dcg_ctrl[25] ),
    .X(_3555_));
 sky130_fd_sc_hd__a221o_1 _7211_ (.A1(\u_reg.reg_7[25] ),
    .A2(net605),
    .B1(net595),
    .B2(\u_reg.reg_3[25] ),
    .C1(_3554_),
    .X(_3556_));
 sky130_fd_sc_hd__a211o_1 _7212_ (.A1(\u_reg.reg_5[25] ),
    .A2(net623),
    .B1(_3555_),
    .C1(_3556_),
    .X(_3557_));
 sky130_fd_sc_hd__mux2_1 _7213_ (.A0(\u_reg.reg_rdata[25] ),
    .A1(net479),
    .S(net576),
    .X(_1400_));
 sky130_fd_sc_hd__a22o_1 _7214_ (.A1(\u_reg.reg_6[26] ),
    .A2(net611),
    .B1(net548),
    .B2(net1820),
    .X(_3558_));
 sky130_fd_sc_hd__a22o_1 _7215_ (.A1(\u_reg.reg_7[26] ),
    .A2(net607),
    .B1(net596),
    .B2(\u_reg.reg_3[26] ),
    .X(_3559_));
 sky130_fd_sc_hd__a221o_1 _7216_ (.A1(\u_reg.reg_4[26] ),
    .A2(net600),
    .B1(net590),
    .B2(\u_reg.reg_2[26] ),
    .C1(_3559_),
    .X(_3560_));
 sky130_fd_sc_hd__a211o_1 _7217_ (.A1(\u_reg.reg_5[26] ),
    .A2(net623),
    .B1(net1821),
    .C1(_3560_),
    .X(_3561_));
 sky130_fd_sc_hd__mux2_1 _7218_ (.A0(\u_reg.reg_rdata[26] ),
    .A1(net1822),
    .S(net576),
    .X(_1401_));
 sky130_fd_sc_hd__a22o_1 _7219_ (.A1(\u_reg.reg_7[27] ),
    .A2(net607),
    .B1(net596),
    .B2(\u_reg.reg_3[27] ),
    .X(_3562_));
 sky130_fd_sc_hd__a22o_1 _7220_ (.A1(\u_reg.reg_6[27] ),
    .A2(net615),
    .B1(net548),
    .B2(\u_reg.cfg_dcg_ctrl[27] ),
    .X(_3563_));
 sky130_fd_sc_hd__a221o_2 _7221_ (.A1(\u_reg.reg_4[27] ),
    .A2(net601),
    .B1(net590),
    .B2(\u_reg.reg_2[27] ),
    .C1(_3562_),
    .X(_3564_));
 sky130_fd_sc_hd__a211o_1 _7222_ (.A1(\u_reg.reg_5[27] ),
    .A2(net624),
    .B1(_3563_),
    .C1(_3564_),
    .X(_3565_));
 sky130_fd_sc_hd__mux2_1 _7223_ (.A0(\u_reg.reg_rdata[27] ),
    .A1(net478),
    .S(net576),
    .X(_1402_));
 sky130_fd_sc_hd__a22o_1 _7224_ (.A1(\u_reg.reg_6[28] ),
    .A2(net613),
    .B1(net548),
    .B2(\u_reg.cfg_dcg_ctrl[28] ),
    .X(_3566_));
 sky130_fd_sc_hd__a22o_1 _7225_ (.A1(\u_reg.reg_4[28] ),
    .A2(net600),
    .B1(net590),
    .B2(\u_reg.reg_2[28] ),
    .X(_3567_));
 sky130_fd_sc_hd__a221o_1 _7226_ (.A1(\u_reg.reg_7[28] ),
    .A2(net607),
    .B1(net596),
    .B2(\u_reg.reg_3[28] ),
    .C1(_3567_),
    .X(_3568_));
 sky130_fd_sc_hd__a211o_2 _7227_ (.A1(\u_reg.reg_5[28] ),
    .A2(net624),
    .B1(_3566_),
    .C1(_3568_),
    .X(_3569_));
 sky130_fd_sc_hd__mux2_1 _7228_ (.A0(\u_reg.reg_rdata[28] ),
    .A1(_3569_),
    .S(net576),
    .X(_1403_));
 sky130_fd_sc_hd__a22o_1 _7229_ (.A1(\u_reg.reg_6[29] ),
    .A2(net613),
    .B1(net547),
    .B2(\u_reg.cfg_dcg_ctrl[29] ),
    .X(_3570_));
 sky130_fd_sc_hd__a22o_1 _7230_ (.A1(\u_reg.reg_4[29] ),
    .A2(net600),
    .B1(net590),
    .B2(\u_reg.reg_2[29] ),
    .X(_3571_));
 sky130_fd_sc_hd__a221o_1 _7231_ (.A1(\u_reg.reg_7[29] ),
    .A2(net605),
    .B1(net595),
    .B2(\u_reg.reg_3[29] ),
    .C1(_3571_),
    .X(_3572_));
 sky130_fd_sc_hd__a211o_2 _7232_ (.A1(\u_reg.reg_5[29] ),
    .A2(net624),
    .B1(_3570_),
    .C1(_3572_),
    .X(_3573_));
 sky130_fd_sc_hd__mux2_1 _7233_ (.A0(\u_reg.reg_rdata[29] ),
    .A1(_3573_),
    .S(net576),
    .X(_1404_));
 sky130_fd_sc_hd__a22o_1 _7234_ (.A1(\u_reg.reg_6[30] ),
    .A2(net615),
    .B1(net547),
    .B2(\u_reg.cfg_dcg_ctrl[30] ),
    .X(_3574_));
 sky130_fd_sc_hd__a22o_1 _7235_ (.A1(\u_reg.reg_4[30] ),
    .A2(net601),
    .B1(net590),
    .B2(\u_reg.reg_2[30] ),
    .X(_3575_));
 sky130_fd_sc_hd__a221o_1 _7236_ (.A1(\u_reg.reg_7[30] ),
    .A2(net605),
    .B1(net595),
    .B2(\u_reg.reg_3[30] ),
    .C1(_3575_),
    .X(_3576_));
 sky130_fd_sc_hd__a211o_1 _7237_ (.A1(\u_reg.reg_5[30] ),
    .A2(net623),
    .B1(_3574_),
    .C1(_3576_),
    .X(_3577_));
 sky130_fd_sc_hd__mux2_1 _7238_ (.A0(\u_reg.reg_rdata[30] ),
    .A1(net477),
    .S(net576),
    .X(_1405_));
 sky130_fd_sc_hd__a22o_1 _7239_ (.A1(\u_reg.reg_4[31] ),
    .A2(net600),
    .B1(net588),
    .B2(\u_reg.reg_2[31] ),
    .X(_3578_));
 sky130_fd_sc_hd__a22o_1 _7240_ (.A1(\u_reg.reg_6[31] ),
    .A2(net611),
    .B1(net546),
    .B2(\u_reg.cfg_dcg_ctrl[31] ),
    .X(_3579_));
 sky130_fd_sc_hd__a221o_1 _7241_ (.A1(\u_reg.reg_7[31] ),
    .A2(net604),
    .B1(net596),
    .B2(\u_reg.reg_3[31] ),
    .C1(_3578_),
    .X(_3580_));
 sky130_fd_sc_hd__a211o_1 _7242_ (.A1(\u_reg.reg_5[31] ),
    .A2(net624),
    .B1(_3579_),
    .C1(_3580_),
    .X(_3581_));
 sky130_fd_sc_hd__mux2_1 _7243_ (.A0(\u_reg.reg_rdata[31] ),
    .A1(_3581_),
    .S(net577),
    .X(_1406_));
 sky130_fd_sc_hd__and3b_4 _7244_ (.A_N(net618),
    .B(_2694_),
    .C(net545),
    .X(_3582_));
 sky130_fd_sc_hd__mux2_1 _7245_ (.A0(\u_dcg_s0.cfg_mode[0] ),
    .A1(_2697_),
    .S(_3582_),
    .X(_1407_));
 sky130_fd_sc_hd__mux2_1 _7246_ (.A0(\u_dcg_s0.cfg_mode[1] ),
    .A1(_2700_),
    .S(_3582_),
    .X(_1408_));
 sky130_fd_sc_hd__mux2_1 _7247_ (.A0(\u_dcg_s1.cfg_mode[0] ),
    .A1(_2703_),
    .S(_3582_),
    .X(_1409_));
 sky130_fd_sc_hd__mux2_1 _7248_ (.A0(\u_dcg_s1.cfg_mode[1] ),
    .A1(_2705_),
    .S(_3582_),
    .X(_1410_));
 sky130_fd_sc_hd__mux2_1 _7249_ (.A0(\u_dcg_s2.cfg_mode[0] ),
    .A1(_2707_),
    .S(_3582_),
    .X(_1411_));
 sky130_fd_sc_hd__mux2_1 _7250_ (.A0(\u_dcg_s2.cfg_mode[1] ),
    .A1(_2709_),
    .S(_3582_),
    .X(_1412_));
 sky130_fd_sc_hd__mux2_1 _7251_ (.A0(\u_dcg_peri.cfg_mode[0] ),
    .A1(_2712_),
    .S(_3582_),
    .X(_1413_));
 sky130_fd_sc_hd__mux2_1 _7252_ (.A0(\u_dcg_peri.cfg_mode[1] ),
    .A1(_2714_),
    .S(_3582_),
    .X(_1414_));
 sky130_fd_sc_hd__and3b_4 _7253_ (.A_N(net618),
    .B(_2694_),
    .C(net587),
    .X(_3583_));
 sky130_fd_sc_hd__mux2_1 _7254_ (.A0(\u_reg.reg_2[0] ),
    .A1(_2697_),
    .S(_3583_),
    .X(_1415_));
 sky130_fd_sc_hd__mux2_1 _7255_ (.A0(\u_reg.reg_2[1] ),
    .A1(_2700_),
    .S(_3583_),
    .X(_1416_));
 sky130_fd_sc_hd__mux2_1 _7256_ (.A0(\u_reg.reg_2[2] ),
    .A1(_2703_),
    .S(_3583_),
    .X(_1417_));
 sky130_fd_sc_hd__mux2_1 _7257_ (.A0(\u_reg.reg_2[3] ),
    .A1(_2705_),
    .S(_3583_),
    .X(_1418_));
 sky130_fd_sc_hd__mux2_1 _7258_ (.A0(\u_reg.reg_2[4] ),
    .A1(_2707_),
    .S(_3583_),
    .X(_1419_));
 sky130_fd_sc_hd__mux2_1 _7259_ (.A0(\u_reg.reg_2[5] ),
    .A1(_2709_),
    .S(_3583_),
    .X(_1420_));
 sky130_fd_sc_hd__mux2_1 _7260_ (.A0(\u_reg.reg_2[6] ),
    .A1(_2712_),
    .S(_3583_),
    .X(_1421_));
 sky130_fd_sc_hd__mux2_1 _7261_ (.A0(\u_reg.reg_2[7] ),
    .A1(_2714_),
    .S(_3583_),
    .X(_1422_));
 sky130_fd_sc_hd__and3b_4 _7262_ (.A_N(net620),
    .B(net617),
    .C(net593),
    .X(_3584_));
 sky130_fd_sc_hd__mux2_1 _7263_ (.A0(\u_reg.reg_3[16] ),
    .A1(net708),
    .S(net517),
    .X(_1423_));
 sky130_fd_sc_hd__mux2_1 _7264_ (.A0(\u_reg.reg_3[17] ),
    .A1(net707),
    .S(net517),
    .X(_1424_));
 sky130_fd_sc_hd__mux2_1 _7265_ (.A0(\u_reg.reg_3[18] ),
    .A1(_2678_),
    .S(_3584_),
    .X(_1425_));
 sky130_fd_sc_hd__mux2_1 _7266_ (.A0(\u_reg.reg_3[19] ),
    .A1(_2681_),
    .S(_3584_),
    .X(_1426_));
 sky130_fd_sc_hd__mux2_1 _7267_ (.A0(\u_reg.reg_3[20] ),
    .A1(net706),
    .S(net517),
    .X(_1427_));
 sky130_fd_sc_hd__mux2_1 _7268_ (.A0(\u_reg.reg_3[21] ),
    .A1(net705),
    .S(net517),
    .X(_1428_));
 sky130_fd_sc_hd__mux2_1 _7269_ (.A0(\u_reg.reg_3[22] ),
    .A1(_2688_),
    .S(_3584_),
    .X(_1429_));
 sky130_fd_sc_hd__mux2_1 _7270_ (.A0(\u_reg.reg_3[23] ),
    .A1(net704),
    .S(_3584_),
    .X(_1430_));
 sky130_fd_sc_hd__and3b_1 _7271_ (.A_N(net619),
    .B(net600),
    .C(net592),
    .X(_3585_));
 sky130_fd_sc_hd__mux2_1 _7272_ (.A0(\u_reg.reg_4[24] ),
    .A1(net695),
    .S(net516),
    .X(_1431_));
 sky130_fd_sc_hd__mux2_1 _7273_ (.A0(\u_reg.reg_4[25] ),
    .A1(net693),
    .S(net516),
    .X(_1432_));
 sky130_fd_sc_hd__mux2_1 _7274_ (.A0(\u_reg.reg_4[26] ),
    .A1(net692),
    .S(net516),
    .X(_1433_));
 sky130_fd_sc_hd__mux2_1 _7275_ (.A0(\u_reg.reg_4[27] ),
    .A1(net691),
    .S(net516),
    .X(_1434_));
 sky130_fd_sc_hd__mux2_1 _7276_ (.A0(\u_reg.reg_4[28] ),
    .A1(net690),
    .S(net516),
    .X(_1435_));
 sky130_fd_sc_hd__mux2_1 _7277_ (.A0(\u_reg.reg_4[29] ),
    .A1(net689),
    .S(net516),
    .X(_1436_));
 sky130_fd_sc_hd__mux2_1 _7278_ (.A0(\u_reg.reg_4[30] ),
    .A1(net688),
    .S(net516),
    .X(_1437_));
 sky130_fd_sc_hd__mux2_1 _7279_ (.A0(\u_reg.reg_4[31] ),
    .A1(net687),
    .S(_3585_),
    .X(_1438_));
 sky130_fd_sc_hd__and4b_2 _7280_ (.A_N(net711),
    .B(net622),
    .C(_2664_),
    .D(net592),
    .X(_3586_));
 sky130_fd_sc_hd__mux2_1 _7281_ (.A0(\u_reg.reg_5[24] ),
    .A1(net695),
    .S(net515),
    .X(_1439_));
 sky130_fd_sc_hd__mux2_1 _7282_ (.A0(\u_reg.reg_5[25] ),
    .A1(net693),
    .S(net515),
    .X(_1440_));
 sky130_fd_sc_hd__mux2_1 _7283_ (.A0(\u_reg.reg_5[26] ),
    .A1(net692),
    .S(net515),
    .X(_1441_));
 sky130_fd_sc_hd__mux2_1 _7284_ (.A0(\u_reg.reg_5[27] ),
    .A1(net691),
    .S(net515),
    .X(_1442_));
 sky130_fd_sc_hd__mux2_1 _7285_ (.A0(\u_reg.reg_5[28] ),
    .A1(net690),
    .S(net515),
    .X(_1443_));
 sky130_fd_sc_hd__mux2_1 _7286_ (.A0(\u_reg.reg_5[29] ),
    .A1(net689),
    .S(net515),
    .X(_1444_));
 sky130_fd_sc_hd__mux2_1 _7287_ (.A0(\u_reg.reg_5[30] ),
    .A1(net688),
    .S(net515),
    .X(_1445_));
 sky130_fd_sc_hd__mux2_1 _7288_ (.A0(\u_reg.reg_5[31] ),
    .A1(net687),
    .S(_3586_),
    .X(_1446_));
 sky130_fd_sc_hd__and3b_4 _7289_ (.A_N(net619),
    .B(net613),
    .C(net592),
    .X(_3587_));
 sky130_fd_sc_hd__mux2_1 _7290_ (.A0(\u_reg.reg_6[24] ),
    .A1(net695),
    .S(_3587_),
    .X(_1447_));
 sky130_fd_sc_hd__mux2_1 _7291_ (.A0(\u_reg.reg_6[25] ),
    .A1(net693),
    .S(_3587_),
    .X(_1448_));
 sky130_fd_sc_hd__mux2_1 _7292_ (.A0(\u_reg.reg_6[26] ),
    .A1(net692),
    .S(_3587_),
    .X(_1449_));
 sky130_fd_sc_hd__mux2_1 _7293_ (.A0(\u_reg.reg_6[27] ),
    .A1(net691),
    .S(_3587_),
    .X(_1450_));
 sky130_fd_sc_hd__mux2_1 _7294_ (.A0(\u_reg.reg_6[28] ),
    .A1(net690),
    .S(_3587_),
    .X(_1451_));
 sky130_fd_sc_hd__mux2_1 _7295_ (.A0(\u_reg.reg_6[29] ),
    .A1(net689),
    .S(_3587_),
    .X(_1452_));
 sky130_fd_sc_hd__mux2_1 _7296_ (.A0(\u_reg.reg_6[30] ),
    .A1(net688),
    .S(_3587_),
    .X(_1453_));
 sky130_fd_sc_hd__mux2_1 _7297_ (.A0(\u_reg.reg_6[31] ),
    .A1(net687),
    .S(_3587_),
    .X(_1454_));
 sky130_fd_sc_hd__nand2_2 _7298_ (.A(net1511),
    .B(net737),
    .Y(_3588_));
 sky130_fd_sc_hd__nor2_1 _7299_ (.A(\u_dcg_s0.hcnt[1] ),
    .B(\u_dcg_s0.hcnt[2] ),
    .Y(_3589_));
 sky130_fd_sc_hd__nand2_1 _7300_ (.A(_1698_),
    .B(_3589_),
    .Y(_3590_));
 sky130_fd_sc_hd__a21o_1 _7301_ (.A1(_1697_),
    .A2(_3590_),
    .B1(_3588_),
    .X(_1455_));
 sky130_fd_sc_hd__xnor2_1 _7302_ (.A(\u_dcg_s0.hcnt[1] ),
    .B(\u_dcg_s0.hcnt[0] ),
    .Y(_3591_));
 sky130_fd_sc_hd__a21o_1 _7303_ (.A1(_3590_),
    .A2(_3591_),
    .B1(_3588_),
    .X(_1456_));
 sky130_fd_sc_hd__o21a_1 _7304_ (.A1(\u_dcg_s0.hcnt[1] ),
    .A2(\u_dcg_s0.hcnt[0] ),
    .B1(\u_dcg_s0.hcnt[2] ),
    .X(_3592_));
 sky130_fd_sc_hd__a311o_1 _7305_ (.A1(_1697_),
    .A2(\u_dcg_s0.hcnt[3] ),
    .A3(_3589_),
    .B1(_3592_),
    .C1(_3588_),
    .X(_1457_));
 sky130_fd_sc_hd__a211oi_1 _7306_ (.A1(_1697_),
    .A2(_3589_),
    .B1(_3588_),
    .C1(_1698_),
    .Y(_1458_));
 sky130_fd_sc_hd__or3b_4 _7307_ (.A(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .B(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .C_N(\u_s1.u_sync_wbb.m_cmd_wr_en ),
    .X(_3593_));
 sky130_fd_sc_hd__mux2_1 _7308_ (.A0(net797),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][1] ),
    .S(net932),
    .X(_1459_));
 sky130_fd_sc_hd__mux2_1 _7309_ (.A0(net798),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][2] ),
    .S(net931),
    .X(_1460_));
 sky130_fd_sc_hd__mux2_1 _7310_ (.A0(_1860_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][3] ),
    .S(net934),
    .X(_1461_));
 sky130_fd_sc_hd__mux2_1 _7311_ (.A0(_1856_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][4] ),
    .S(net932),
    .X(_1462_));
 sky130_fd_sc_hd__mux2_1 _7312_ (.A0(_1869_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][5] ),
    .S(net935),
    .X(_1463_));
 sky130_fd_sc_hd__mux2_1 _7313_ (.A0(_1868_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][6] ),
    .S(net934),
    .X(_1464_));
 sky130_fd_sc_hd__mux2_1 _7314_ (.A0(_1867_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][7] ),
    .S(net931),
    .X(_1465_));
 sky130_fd_sc_hd__mux2_1 _7315_ (.A0(_1866_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][8] ),
    .S(net934),
    .X(_1466_));
 sky130_fd_sc_hd__mux2_1 _7316_ (.A0(_1873_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][9] ),
    .S(net931),
    .X(_1467_));
 sky130_fd_sc_hd__mux2_1 _7317_ (.A0(net686),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][14] ),
    .S(net935),
    .X(_1468_));
 sky130_fd_sc_hd__mux2_1 _7318_ (.A0(net685),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][15] ),
    .S(net932),
    .X(_1469_));
 sky130_fd_sc_hd__mux2_1 _7319_ (.A0(net684),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][16] ),
    .S(net934),
    .X(_1470_));
 sky130_fd_sc_hd__mux2_1 _7320_ (.A0(net683),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][17] ),
    .S(net934),
    .X(_1471_));
 sky130_fd_sc_hd__mux2_1 _7321_ (.A0(net682),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][18] ),
    .S(net935),
    .X(_1472_));
 sky130_fd_sc_hd__mux2_1 _7322_ (.A0(_2816_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][19] ),
    .S(net936),
    .X(_1473_));
 sky130_fd_sc_hd__mux2_1 _7323_ (.A0(_2818_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][20] ),
    .S(net932),
    .X(_1474_));
 sky130_fd_sc_hd__mux2_1 _7324_ (.A0(net681),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][21] ),
    .S(net934),
    .X(_1475_));
 sky130_fd_sc_hd__mux2_1 _7325_ (.A0(_2823_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][22] ),
    .S(net935),
    .X(_1476_));
 sky130_fd_sc_hd__mux2_1 _7326_ (.A0(_2825_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][23] ),
    .S(net935),
    .X(_1477_));
 sky130_fd_sc_hd__mux2_1 _7327_ (.A0(_2827_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][24] ),
    .S(net932),
    .X(_1478_));
 sky130_fd_sc_hd__mux2_1 _7328_ (.A0(_2830_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][25] ),
    .S(net935),
    .X(_1479_));
 sky130_fd_sc_hd__mux2_1 _7329_ (.A0(_2832_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][26] ),
    .S(net936),
    .X(_1480_));
 sky130_fd_sc_hd__mux2_1 _7330_ (.A0(_2835_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][27] ),
    .S(net936),
    .X(_1481_));
 sky130_fd_sc_hd__mux2_1 _7331_ (.A0(_2838_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][28] ),
    .S(net935),
    .X(_1482_));
 sky130_fd_sc_hd__mux2_1 _7332_ (.A0(_2841_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][29] ),
    .S(net936),
    .X(_1483_));
 sky130_fd_sc_hd__mux2_1 _7333_ (.A0(_2844_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][30] ),
    .S(net936),
    .X(_1484_));
 sky130_fd_sc_hd__mux2_1 _7334_ (.A0(_2846_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][31] ),
    .S(net932),
    .X(_1485_));
 sky130_fd_sc_hd__mux2_1 _7335_ (.A0(_2849_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][32] ),
    .S(net934),
    .X(_1486_));
 sky130_fd_sc_hd__mux2_1 _7336_ (.A0(_2851_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][33] ),
    .S(net931),
    .X(_1487_));
 sky130_fd_sc_hd__mux2_1 _7337_ (.A0(_2854_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][34] ),
    .S(net936),
    .X(_1488_));
 sky130_fd_sc_hd__mux2_1 _7338_ (.A0(_2856_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][35] ),
    .S(net935),
    .X(_1489_));
 sky130_fd_sc_hd__mux2_1 _7339_ (.A0(_2858_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][36] ),
    .S(net933),
    .X(_1490_));
 sky130_fd_sc_hd__mux2_1 _7340_ (.A0(_2861_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][37] ),
    .S(net934),
    .X(_1491_));
 sky130_fd_sc_hd__mux2_1 _7341_ (.A0(_2863_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][38] ),
    .S(net934),
    .X(_1492_));
 sky130_fd_sc_hd__mux2_1 _7342_ (.A0(_2865_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][39] ),
    .S(net931),
    .X(_1493_));
 sky130_fd_sc_hd__mux2_1 _7343_ (.A0(_2867_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][40] ),
    .S(net933),
    .X(_1494_));
 sky130_fd_sc_hd__mux2_1 _7344_ (.A0(_2869_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][41] ),
    .S(net934),
    .X(_1495_));
 sky130_fd_sc_hd__mux2_1 _7345_ (.A0(net680),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][42] ),
    .S(net935),
    .X(_1496_));
 sky130_fd_sc_hd__mux2_1 _7346_ (.A0(net2080),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][43] ),
    .S(net932),
    .X(_1497_));
 sky130_fd_sc_hd__mux2_1 _7347_ (.A0(_2875_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][44] ),
    .S(net931),
    .X(_1498_));
 sky130_fd_sc_hd__mux2_1 _7348_ (.A0(_2877_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][45] ),
    .S(net935),
    .X(_1499_));
 sky130_fd_sc_hd__mux2_1 _7349_ (.A0(net679),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][46] ),
    .S(net936),
    .X(_1500_));
 sky130_fd_sc_hd__mux2_1 _7350_ (.A0(_2881_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][47] ),
    .S(net933),
    .X(_1501_));
 sky130_fd_sc_hd__mux2_1 _7351_ (.A0(_2883_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][48] ),
    .S(net931),
    .X(_1502_));
 sky130_fd_sc_hd__mux2_1 _7352_ (.A0(_2885_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][49] ),
    .S(net931),
    .X(_1503_));
 sky130_fd_sc_hd__mux2_1 _7353_ (.A0(net732),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][50] ),
    .S(net936),
    .X(_1504_));
 sky130_fd_sc_hd__mux2_1 _7354_ (.A0(_2888_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][53] ),
    .S(net931),
    .X(_1505_));
 sky130_fd_sc_hd__mux2_1 _7355_ (.A0(_2891_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][54] ),
    .S(net932),
    .X(_1506_));
 sky130_fd_sc_hd__mux2_1 _7356_ (.A0(_2894_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][55] ),
    .S(net932),
    .X(_1507_));
 sky130_fd_sc_hd__mux2_1 _7357_ (.A0(_2897_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][56] ),
    .S(net933),
    .X(_1508_));
 sky130_fd_sc_hd__mux2_1 _7358_ (.A0(_2900_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][57] ),
    .S(net933),
    .X(_1509_));
 sky130_fd_sc_hd__mux2_1 _7359_ (.A0(_2903_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][58] ),
    .S(net932),
    .X(_1510_));
 sky130_fd_sc_hd__mux2_1 _7360_ (.A0(_2906_),
    .A1(\u_s1.u_sync_wbb.u_cmd_if.mem[0][59] ),
    .S(net931),
    .X(_1511_));
 sky130_fd_sc_hd__mux2_1 _7361_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][0] ),
    .A1(_1786_),
    .S(net744),
    .X(_1512_));
 sky130_fd_sc_hd__mux2_1 _7362_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][1] ),
    .A1(_1789_),
    .S(net740),
    .X(_1513_));
 sky130_fd_sc_hd__mux2_1 _7363_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][2] ),
    .A1(_1792_),
    .S(net746),
    .X(_1514_));
 sky130_fd_sc_hd__mux2_1 _7364_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][3] ),
    .A1(_1794_),
    .S(net746),
    .X(_1515_));
 sky130_fd_sc_hd__mux2_1 _7365_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][4] ),
    .A1(_1793_),
    .S(net746),
    .X(_1516_));
 sky130_fd_sc_hd__mux2_1 _7366_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][5] ),
    .A1(net808),
    .S(net746),
    .X(_1517_));
 sky130_fd_sc_hd__mux2_1 _7367_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][6] ),
    .A1(_1797_),
    .S(net746),
    .X(_1518_));
 sky130_fd_sc_hd__mux2_1 _7368_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][7] ),
    .A1(_1796_),
    .S(net747),
    .X(_1519_));
 sky130_fd_sc_hd__mux2_1 _7369_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][8] ),
    .A1(_1799_),
    .S(net746),
    .X(_1520_));
 sky130_fd_sc_hd__mux2_1 _7370_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][9] ),
    .A1(_1787_),
    .S(net745),
    .X(_1521_));
 sky130_fd_sc_hd__mux2_1 _7371_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][14] ),
    .A1(_2948_),
    .S(net743),
    .X(_1522_));
 sky130_fd_sc_hd__mux2_1 _7372_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][15] ),
    .A1(_2951_),
    .S(net740),
    .X(_1523_));
 sky130_fd_sc_hd__mux2_1 _7373_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][16] ),
    .A1(_2954_),
    .S(net741),
    .X(_1524_));
 sky130_fd_sc_hd__mux2_1 _7374_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][17] ),
    .A1(_2957_),
    .S(net741),
    .X(_1525_));
 sky130_fd_sc_hd__mux2_1 _7375_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][18] ),
    .A1(_2960_),
    .S(net747),
    .X(_1526_));
 sky130_fd_sc_hd__mux2_1 _7376_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][19] ),
    .A1(_2962_),
    .S(net746),
    .X(_1527_));
 sky130_fd_sc_hd__mux2_1 _7377_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][20] ),
    .A1(_2964_),
    .S(net747),
    .X(_1528_));
 sky130_fd_sc_hd__mux2_1 _7378_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][21] ),
    .A1(_2966_),
    .S(net747),
    .X(_1529_));
 sky130_fd_sc_hd__mux2_1 _7379_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][22] ),
    .A1(_2969_),
    .S(net744),
    .X(_1530_));
 sky130_fd_sc_hd__mux2_1 _7380_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][23] ),
    .A1(_2971_),
    .S(net744),
    .X(_1531_));
 sky130_fd_sc_hd__mux2_1 _7381_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][24] ),
    .A1(_2973_),
    .S(net745),
    .X(_1532_));
 sky130_fd_sc_hd__mux2_1 _7382_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][25] ),
    .A1(_2976_),
    .S(net743),
    .X(_1533_));
 sky130_fd_sc_hd__mux2_1 _7383_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][26] ),
    .A1(_2979_),
    .S(net745),
    .X(_1534_));
 sky130_fd_sc_hd__mux2_1 _7384_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][27] ),
    .A1(_2981_),
    .S(net746),
    .X(_1535_));
 sky130_fd_sc_hd__mux2_1 _7385_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][28] ),
    .A1(_2983_),
    .S(net746),
    .X(_1536_));
 sky130_fd_sc_hd__mux2_1 _7386_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][29] ),
    .A1(_2985_),
    .S(net747),
    .X(_1537_));
 sky130_fd_sc_hd__mux2_1 _7387_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][30] ),
    .A1(_2988_),
    .S(net740),
    .X(_1538_));
 sky130_fd_sc_hd__mux2_1 _7388_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][31] ),
    .A1(_2991_),
    .S(net742),
    .X(_1539_));
 sky130_fd_sc_hd__mux2_1 _7389_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][32] ),
    .A1(_2993_),
    .S(net747),
    .X(_1540_));
 sky130_fd_sc_hd__mux2_1 _7390_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][33] ),
    .A1(_2995_),
    .S(net744),
    .X(_1541_));
 sky130_fd_sc_hd__mux2_1 _7391_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][34] ),
    .A1(_2998_),
    .S(net742),
    .X(_1542_));
 sky130_fd_sc_hd__mux2_1 _7392_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][35] ),
    .A1(_3001_),
    .S(net746),
    .X(_1543_));
 sky130_fd_sc_hd__mux2_1 _7393_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][36] ),
    .A1(_3004_),
    .S(net741),
    .X(_1544_));
 sky130_fd_sc_hd__mux2_1 _7394_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][37] ),
    .A1(net2009),
    .S(net744),
    .X(_1545_));
 sky130_fd_sc_hd__mux2_1 _7395_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][38] ),
    .A1(_3010_),
    .S(net741),
    .X(_1546_));
 sky130_fd_sc_hd__mux2_1 _7396_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][39] ),
    .A1(_3012_),
    .S(net745),
    .X(_1547_));
 sky130_fd_sc_hd__mux2_1 _7397_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][40] ),
    .A1(_3014_),
    .S(net742),
    .X(_1548_));
 sky130_fd_sc_hd__mux2_1 _7398_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][41] ),
    .A1(_3016_),
    .S(net745),
    .X(_1549_));
 sky130_fd_sc_hd__mux2_1 _7399_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][42] ),
    .A1(net2017),
    .S(net743),
    .X(_1550_));
 sky130_fd_sc_hd__mux2_1 _7400_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][43] ),
    .A1(net2038),
    .S(net744),
    .X(_1551_));
 sky130_fd_sc_hd__mux2_1 _7401_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][44] ),
    .A1(_3024_),
    .S(net743),
    .X(_1552_));
 sky130_fd_sc_hd__mux2_1 _7402_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][45] ),
    .A1(_3026_),
    .S(net743),
    .X(_1553_));
 sky130_fd_sc_hd__mux2_1 _7403_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][46] ),
    .A1(_3029_),
    .S(net741),
    .X(_1554_));
 sky130_fd_sc_hd__mux2_1 _7404_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][47] ),
    .A1(_3031_),
    .S(net743),
    .X(_1555_));
 sky130_fd_sc_hd__mux2_1 _7405_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][48] ),
    .A1(_3033_),
    .S(net744),
    .X(_1556_));
 sky130_fd_sc_hd__mux2_1 _7406_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][49] ),
    .A1(net2058),
    .S(net741),
    .X(_1557_));
 sky130_fd_sc_hd__mux2_1 _7407_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][50] ),
    .A1(_1806_),
    .S(net744),
    .X(_1558_));
 sky130_fd_sc_hd__mux2_1 _7408_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][53] ),
    .A1(_3038_),
    .S(net744),
    .X(_1559_));
 sky130_fd_sc_hd__mux2_1 _7409_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][54] ),
    .A1(_3041_),
    .S(net742),
    .X(_1560_));
 sky130_fd_sc_hd__mux2_1 _7410_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][55] ),
    .A1(_3044_),
    .S(net744),
    .X(_1561_));
 sky130_fd_sc_hd__mux2_1 _7411_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][56] ),
    .A1(_3047_),
    .S(net743),
    .X(_1562_));
 sky130_fd_sc_hd__mux2_1 _7412_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][57] ),
    .A1(_3050_),
    .S(net741),
    .X(_1563_));
 sky130_fd_sc_hd__mux2_1 _7413_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][58] ),
    .A1(_3053_),
    .S(net739),
    .X(_1564_));
 sky130_fd_sc_hd__mux2_1 _7414_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][59] ),
    .A1(net2022),
    .S(net743),
    .X(_1565_));
 sky130_fd_sc_hd__mux2_1 _7415_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][60] ),
    .A1(_3059_),
    .S(net742),
    .X(_1566_));
 sky130_fd_sc_hd__mux2_1 _7416_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][61] ),
    .A1(_3062_),
    .S(net743),
    .X(_1567_));
 sky130_fd_sc_hd__mux2_1 _7417_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][62] ),
    .A1(_3065_),
    .S(net740),
    .X(_1568_));
 sky130_fd_sc_hd__mux2_1 _7418_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][63] ),
    .A1(_3068_),
    .S(net740),
    .X(_1569_));
 sky130_fd_sc_hd__mux2_1 _7419_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][64] ),
    .A1(_3071_),
    .S(net742),
    .X(_1570_));
 sky130_fd_sc_hd__mux2_1 _7420_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][65] ),
    .A1(net1998),
    .S(net739),
    .X(_1571_));
 sky130_fd_sc_hd__mux2_1 _7421_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][66] ),
    .A1(net1869),
    .S(net739),
    .X(_1572_));
 sky130_fd_sc_hd__mux2_1 _7422_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][67] ),
    .A1(_3080_),
    .S(net742),
    .X(_1573_));
 sky130_fd_sc_hd__mux2_1 _7423_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][68] ),
    .A1(_3083_),
    .S(net742),
    .X(_1574_));
 sky130_fd_sc_hd__mux2_1 _7424_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][69] ),
    .A1(_3086_),
    .S(net739),
    .X(_1575_));
 sky130_fd_sc_hd__mux2_1 _7425_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][70] ),
    .A1(_3089_),
    .S(net739),
    .X(_1576_));
 sky130_fd_sc_hd__mux2_1 _7426_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][71] ),
    .A1(_3092_),
    .S(net742),
    .X(_1577_));
 sky130_fd_sc_hd__mux2_1 _7427_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][72] ),
    .A1(_3095_),
    .S(net740),
    .X(_1578_));
 sky130_fd_sc_hd__mux2_1 _7428_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][73] ),
    .A1(_3098_),
    .S(net742),
    .X(_1579_));
 sky130_fd_sc_hd__mux2_1 _7429_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][74] ),
    .A1(_3101_),
    .S(net739),
    .X(_1580_));
 sky130_fd_sc_hd__mux2_1 _7430_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][75] ),
    .A1(_3104_),
    .S(net740),
    .X(_1581_));
 sky130_fd_sc_hd__mux2_1 _7431_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][76] ),
    .A1(_3107_),
    .S(net740),
    .X(_1582_));
 sky130_fd_sc_hd__mux2_1 _7432_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][77] ),
    .A1(net1848),
    .S(net740),
    .X(_1583_));
 sky130_fd_sc_hd__mux2_1 _7433_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][78] ),
    .A1(_3113_),
    .S(net739),
    .X(_1584_));
 sky130_fd_sc_hd__mux2_1 _7434_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][79] ),
    .A1(_3116_),
    .S(net740),
    .X(_1585_));
 sky130_fd_sc_hd__mux2_1 _7435_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][80] ),
    .A1(_3119_),
    .S(net739),
    .X(_1586_));
 sky130_fd_sc_hd__mux2_1 _7436_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][81] ),
    .A1(_3122_),
    .S(net739),
    .X(_1587_));
 sky130_fd_sc_hd__mux2_1 _7437_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[1][82] ),
    .A1(net1853),
    .S(net739),
    .X(_1588_));
 sky130_fd_sc_hd__and3b_4 _7438_ (.A_N(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .B(\u_s0.u_sync_wbb.m_cmd_wr_en ),
    .C(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[1] ),
    .X(_3594_));
 sky130_fd_sc_hd__mux2_1 _7439_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][0] ),
    .A1(_1786_),
    .S(net925),
    .X(_1589_));
 sky130_fd_sc_hd__mux2_1 _7440_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][1] ),
    .A1(_1789_),
    .S(net923),
    .X(_1590_));
 sky130_fd_sc_hd__mux2_1 _7441_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][2] ),
    .A1(_1792_),
    .S(net928),
    .X(_1591_));
 sky130_fd_sc_hd__mux2_1 _7442_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][3] ),
    .A1(_1794_),
    .S(net929),
    .X(_1592_));
 sky130_fd_sc_hd__mux2_1 _7443_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][4] ),
    .A1(_1793_),
    .S(net928),
    .X(_1593_));
 sky130_fd_sc_hd__mux2_1 _7444_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][5] ),
    .A1(net808),
    .S(net928),
    .X(_1594_));
 sky130_fd_sc_hd__mux2_1 _7445_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][6] ),
    .A1(_1797_),
    .S(net928),
    .X(_1595_));
 sky130_fd_sc_hd__mux2_1 _7446_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][7] ),
    .A1(_1796_),
    .S(net929),
    .X(_1596_));
 sky130_fd_sc_hd__mux2_1 _7447_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][8] ),
    .A1(_1799_),
    .S(net929),
    .X(_1597_));
 sky130_fd_sc_hd__mux2_1 _7448_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][9] ),
    .A1(_1787_),
    .S(net927),
    .X(_1598_));
 sky130_fd_sc_hd__mux2_1 _7449_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][14] ),
    .A1(_2948_),
    .S(net925),
    .X(_1599_));
 sky130_fd_sc_hd__mux2_1 _7450_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][15] ),
    .A1(_2951_),
    .S(net923),
    .X(_1600_));
 sky130_fd_sc_hd__mux2_1 _7451_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][16] ),
    .A1(_2954_),
    .S(net922),
    .X(_1601_));
 sky130_fd_sc_hd__mux2_1 _7452_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][17] ),
    .A1(_2957_),
    .S(net922),
    .X(_1602_));
 sky130_fd_sc_hd__mux2_1 _7453_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][18] ),
    .A1(_2960_),
    .S(net928),
    .X(_1603_));
 sky130_fd_sc_hd__mux2_1 _7454_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][19] ),
    .A1(_2962_),
    .S(net928),
    .X(_1604_));
 sky130_fd_sc_hd__mux2_1 _7455_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][20] ),
    .A1(_2964_),
    .S(net929),
    .X(_1605_));
 sky130_fd_sc_hd__mux2_1 _7456_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][21] ),
    .A1(_2966_),
    .S(net928),
    .X(_1606_));
 sky130_fd_sc_hd__mux2_1 _7457_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][22] ),
    .A1(net2007),
    .S(net927),
    .X(_1607_));
 sky130_fd_sc_hd__mux2_1 _7458_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][23] ),
    .A1(_2971_),
    .S(net930),
    .X(_1608_));
 sky130_fd_sc_hd__mux2_1 _7459_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][24] ),
    .A1(_2973_),
    .S(net930),
    .X(_1609_));
 sky130_fd_sc_hd__mux2_1 _7460_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][25] ),
    .A1(_2976_),
    .S(net925),
    .X(_1610_));
 sky130_fd_sc_hd__mux2_1 _7461_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][26] ),
    .A1(_2979_),
    .S(net927),
    .X(_1611_));
 sky130_fd_sc_hd__mux2_1 _7462_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][27] ),
    .A1(_2981_),
    .S(net928),
    .X(_1612_));
 sky130_fd_sc_hd__mux2_1 _7463_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][28] ),
    .A1(_2983_),
    .S(net928),
    .X(_1613_));
 sky130_fd_sc_hd__mux2_1 _7464_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][29] ),
    .A1(_2985_),
    .S(net929),
    .X(_1614_));
 sky130_fd_sc_hd__mux2_1 _7465_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][30] ),
    .A1(_2988_),
    .S(net923),
    .X(_1615_));
 sky130_fd_sc_hd__mux2_1 _7466_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][31] ),
    .A1(_2991_),
    .S(net926),
    .X(_1616_));
 sky130_fd_sc_hd__mux2_1 _7467_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][32] ),
    .A1(_2993_),
    .S(net929),
    .X(_1617_));
 sky130_fd_sc_hd__mux2_1 _7468_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][33] ),
    .A1(_2995_),
    .S(net927),
    .X(_1618_));
 sky130_fd_sc_hd__mux2_1 _7469_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][34] ),
    .A1(net2040),
    .S(net925),
    .X(_1619_));
 sky130_fd_sc_hd__mux2_1 _7470_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][35] ),
    .A1(_3001_),
    .S(net928),
    .X(_1620_));
 sky130_fd_sc_hd__mux2_1 _7471_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][36] ),
    .A1(_3004_),
    .S(net924),
    .X(_1621_));
 sky130_fd_sc_hd__mux2_1 _7472_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][37] ),
    .A1(net2009),
    .S(net927),
    .X(_1622_));
 sky130_fd_sc_hd__mux2_1 _7473_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][38] ),
    .A1(_3010_),
    .S(net924),
    .X(_1623_));
 sky130_fd_sc_hd__mux2_1 _7474_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][39] ),
    .A1(_3012_),
    .S(net930),
    .X(_1624_));
 sky130_fd_sc_hd__mux2_1 _7475_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][40] ),
    .A1(_3014_),
    .S(net926),
    .X(_1625_));
 sky130_fd_sc_hd__mux2_1 _7476_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][41] ),
    .A1(_3016_),
    .S(net930),
    .X(_1626_));
 sky130_fd_sc_hd__mux2_1 _7477_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][42] ),
    .A1(net2017),
    .S(net926),
    .X(_1627_));
 sky130_fd_sc_hd__mux2_1 _7478_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][43] ),
    .A1(net2038),
    .S(net927),
    .X(_1628_));
 sky130_fd_sc_hd__mux2_1 _7479_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][44] ),
    .A1(_3024_),
    .S(net926),
    .X(_1629_));
 sky130_fd_sc_hd__mux2_1 _7480_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][45] ),
    .A1(_3026_),
    .S(net925),
    .X(_1630_));
 sky130_fd_sc_hd__mux2_1 _7481_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][46] ),
    .A1(_3029_),
    .S(net922),
    .X(_1631_));
 sky130_fd_sc_hd__mux2_1 _7482_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][47] ),
    .A1(_3031_),
    .S(net927),
    .X(_1632_));
 sky130_fd_sc_hd__mux2_1 _7483_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][48] ),
    .A1(_3033_),
    .S(net927),
    .X(_1633_));
 sky130_fd_sc_hd__mux2_1 _7484_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][49] ),
    .A1(net2058),
    .S(net922),
    .X(_1634_));
 sky130_fd_sc_hd__mux2_1 _7485_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][50] ),
    .A1(_1806_),
    .S(net927),
    .X(_1635_));
 sky130_fd_sc_hd__mux2_1 _7486_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][53] ),
    .A1(_3038_),
    .S(net925),
    .X(_1636_));
 sky130_fd_sc_hd__mux2_1 _7487_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][54] ),
    .A1(_3041_),
    .S(net925),
    .X(_1637_));
 sky130_fd_sc_hd__mux2_1 _7488_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][55] ),
    .A1(_3044_),
    .S(net925),
    .X(_1638_));
 sky130_fd_sc_hd__mux2_1 _7489_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][56] ),
    .A1(_3047_),
    .S(net927),
    .X(_1639_));
 sky130_fd_sc_hd__mux2_1 _7490_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][57] ),
    .A1(_3050_),
    .S(net924),
    .X(_1640_));
 sky130_fd_sc_hd__mux2_1 _7491_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][58] ),
    .A1(_3053_),
    .S(net921),
    .X(_1641_));
 sky130_fd_sc_hd__mux2_1 _7492_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][59] ),
    .A1(net2022),
    .S(net925),
    .X(_1642_));
 sky130_fd_sc_hd__mux2_1 _7493_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][60] ),
    .A1(_3059_),
    .S(net926),
    .X(_1643_));
 sky130_fd_sc_hd__mux2_1 _7494_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][61] ),
    .A1(_3062_),
    .S(net925),
    .X(_1644_));
 sky130_fd_sc_hd__mux2_1 _7495_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][62] ),
    .A1(_3065_),
    .S(net923),
    .X(_1645_));
 sky130_fd_sc_hd__mux2_1 _7496_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][63] ),
    .A1(_3068_),
    .S(net926),
    .X(_1646_));
 sky130_fd_sc_hd__mux2_1 _7497_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][64] ),
    .A1(net1909),
    .S(net923),
    .X(_1647_));
 sky130_fd_sc_hd__mux2_1 _7498_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][65] ),
    .A1(net1998),
    .S(net921),
    .X(_1648_));
 sky130_fd_sc_hd__mux2_1 _7499_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][66] ),
    .A1(net1869),
    .S(net921),
    .X(_1649_));
 sky130_fd_sc_hd__mux2_1 _7500_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][67] ),
    .A1(_3080_),
    .S(net923),
    .X(_1650_));
 sky130_fd_sc_hd__mux2_1 _7501_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][68] ),
    .A1(_3083_),
    .S(net926),
    .X(_1651_));
 sky130_fd_sc_hd__mux2_1 _7502_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][69] ),
    .A1(_3086_),
    .S(net921),
    .X(_1652_));
 sky130_fd_sc_hd__mux2_1 _7503_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][70] ),
    .A1(_3089_),
    .S(net921),
    .X(_1653_));
 sky130_fd_sc_hd__mux2_1 _7504_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][71] ),
    .A1(_3092_),
    .S(net926),
    .X(_1654_));
 sky130_fd_sc_hd__mux2_1 _7505_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][72] ),
    .A1(_3095_),
    .S(net923),
    .X(_1655_));
 sky130_fd_sc_hd__mux2_1 _7506_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][73] ),
    .A1(_3098_),
    .S(net926),
    .X(_1656_));
 sky130_fd_sc_hd__mux2_1 _7507_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][74] ),
    .A1(_3101_),
    .S(net921),
    .X(_1657_));
 sky130_fd_sc_hd__mux2_1 _7508_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][75] ),
    .A1(_3104_),
    .S(net923),
    .X(_1658_));
 sky130_fd_sc_hd__mux2_1 _7509_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][76] ),
    .A1(_3107_),
    .S(net923),
    .X(_1659_));
 sky130_fd_sc_hd__mux2_1 _7510_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][77] ),
    .A1(_3110_),
    .S(net921),
    .X(_1660_));
 sky130_fd_sc_hd__mux2_1 _7511_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][78] ),
    .A1(_3113_),
    .S(net921),
    .X(_1661_));
 sky130_fd_sc_hd__mux2_1 _7512_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][79] ),
    .A1(net1901),
    .S(net923),
    .X(_1662_));
 sky130_fd_sc_hd__mux2_1 _7513_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][80] ),
    .A1(_3119_),
    .S(net921),
    .X(_1663_));
 sky130_fd_sc_hd__mux2_1 _7514_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][81] ),
    .A1(net1867),
    .S(net921),
    .X(_1664_));
 sky130_fd_sc_hd__mux2_1 _7515_ (.A0(\u_s0.u_sync_wbb.u_cmd_if.mem[2][82] ),
    .A1(net1853),
    .S(net922),
    .X(_1665_));
 sky130_fd_sc_hd__or2_1 _7516_ (.A(\u_dcg_s0.hcnt[0] ),
    .B(_3590_),
    .X(_3595_));
 sky130_fd_sc_hd__a21o_1 _7517_ (.A1(\u_dcg_s0.idle_his ),
    .A2(_3595_),
    .B1(_3588_),
    .X(_1666_));
 sky130_fd_sc_hd__a21o_1 _7518_ (.A1(_2012_),
    .A2(_2022_),
    .B1(_2018_),
    .X(_3596_));
 sky130_fd_sc_hd__and3b_1 _7519_ (.A_N(_2648_),
    .B(net1164),
    .C(m1_wbd_stb_i),
    .X(_3597_));
 sky130_fd_sc_hd__nor2_1 _7520_ (.A(net1210),
    .B(_2022_),
    .Y(_3598_));
 sky130_fd_sc_hd__and2b_1 _7521_ (.A_N(_3598_),
    .B(_3597_),
    .X(_3599_));
 sky130_fd_sc_hd__a21oi_1 _7522_ (.A1(m2_wbd_stb_i),
    .A2(net1161),
    .B1(net1275),
    .Y(_3600_));
 sky130_fd_sc_hd__or2_1 _7523_ (.A(_2648_),
    .B(_3600_),
    .X(_3601_));
 sky130_fd_sc_hd__a31o_1 _7524_ (.A1(net1219),
    .A2(net1275),
    .A3(_2022_),
    .B1(_3601_),
    .X(_3602_));
 sky130_fd_sc_hd__a31o_1 _7525_ (.A1(m3_wbd_stb_i),
    .A2(net1157),
    .A3(_3602_),
    .B1(_3599_),
    .X(_3603_));
 sky130_fd_sc_hd__a22o_1 _7526_ (.A1(net1278),
    .A2(_3596_),
    .B1(_3603_),
    .B2(_2023_),
    .X(_1667_));
 sky130_fd_sc_hd__a31o_1 _7527_ (.A1(m0_wbd_stb_i),
    .A2(net1278),
    .A3(net1147),
    .B1(_3600_),
    .X(_3604_));
 sky130_fd_sc_hd__a211oi_1 _7528_ (.A1(_2016_),
    .A2(_3604_),
    .B1(_3598_),
    .C1(_3597_),
    .Y(_3605_));
 sky130_fd_sc_hd__a22o_1 _7529_ (.A1(net1275),
    .A2(_2018_),
    .B1(_2023_),
    .B2(_3605_),
    .X(_1668_));
 sky130_fd_sc_hd__dfrtp_1 _7530_ (.CLK(\clknet_leaf_30_u_dsync.out_clk ),
    .D(_0010_),
    .RESET_B(net913),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7531_ (.CLK(\clknet_leaf_30_u_dsync.out_clk ),
    .D(_0011_),
    .RESET_B(net913),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7532_ (.CLK(\clknet_leaf_30_u_dsync.out_clk ),
    .D(_0012_),
    .RESET_B(net909),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7533_ (.CLK(\clknet_leaf_29_u_dsync.out_clk ),
    .D(_0013_),
    .RESET_B(net913),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7534_ (.CLK(\clknet_leaf_29_u_dsync.out_clk ),
    .D(_0014_),
    .RESET_B(net913),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7535_ (.CLK(\clknet_leaf_29_u_dsync.out_clk ),
    .D(_0015_),
    .RESET_B(net913),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7536_ (.CLK(\clknet_leaf_29_u_dsync.out_clk ),
    .D(_0016_),
    .RESET_B(net914),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7537_ (.CLK(\clknet_leaf_29_u_dsync.out_clk ),
    .D(_0017_),
    .RESET_B(net913),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7538_ (.CLK(\clknet_leaf_32_u_dsync.out_clk ),
    .D(_0018_),
    .RESET_B(net909),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7539_ (.CLK(\clknet_leaf_54_u_dsync.out_clk ),
    .D(_0019_),
    .RESET_B(net904),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7540_ (.CLK(\clknet_leaf_52_u_dsync.out_clk ),
    .D(_0020_),
    .RESET_B(net916),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7541_ (.CLK(\clknet_leaf_51_u_dsync.out_clk ),
    .D(_0021_),
    .RESET_B(net904),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7542_ (.CLK(\clknet_leaf_53_u_dsync.out_clk ),
    .D(_0022_),
    .RESET_B(net902),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7543_ (.CLK(\clknet_leaf_48_u_dsync.out_clk ),
    .D(_0023_),
    .RESET_B(net915),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7544_ (.CLK(\clknet_leaf_47_u_dsync.out_clk ),
    .D(_0024_),
    .RESET_B(net916),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[19] ));
 sky130_fd_sc_hd__dfrtp_1 _7545_ (.CLK(\clknet_leaf_51_u_dsync.out_clk ),
    .D(_0025_),
    .RESET_B(net915),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[20] ));
 sky130_fd_sc_hd__dfrtp_1 _7546_ (.CLK(\clknet_leaf_42_u_dsync.out_clk ),
    .D(_0026_),
    .RESET_B(net903),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[21] ));
 sky130_fd_sc_hd__dfrtp_1 _7547_ (.CLK(\clknet_leaf_47_u_dsync.out_clk ),
    .D(_0027_),
    .RESET_B(net916),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[22] ));
 sky130_fd_sc_hd__dfrtp_1 _7548_ (.CLK(\clknet_leaf_45_u_dsync.out_clk ),
    .D(_0028_),
    .RESET_B(net915),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[23] ));
 sky130_fd_sc_hd__dfrtp_1 _7549_ (.CLK(\clknet_leaf_49_u_dsync.out_clk ),
    .D(_0029_),
    .RESET_B(net904),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[24] ));
 sky130_fd_sc_hd__dfrtp_1 _7550_ (.CLK(\clknet_leaf_49_u_dsync.out_clk ),
    .D(_0030_),
    .RESET_B(net915),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[25] ));
 sky130_fd_sc_hd__dfrtp_1 _7551_ (.CLK(\clknet_leaf_53_u_dsync.out_clk ),
    .D(_0031_),
    .RESET_B(net902),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[26] ));
 sky130_fd_sc_hd__dfrtp_1 _7552_ (.CLK(\clknet_leaf_54_u_dsync.out_clk ),
    .D(_0032_),
    .RESET_B(net902),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[27] ));
 sky130_fd_sc_hd__dfrtp_1 _7553_ (.CLK(\clknet_leaf_47_u_dsync.out_clk ),
    .D(_0033_),
    .RESET_B(net916),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[28] ));
 sky130_fd_sc_hd__dfrtp_1 _7554_ (.CLK(\clknet_leaf_49_u_dsync.out_clk ),
    .D(_0034_),
    .RESET_B(net903),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[29] ));
 sky130_fd_sc_hd__dfrtp_1 _7555_ (.CLK(\clknet_leaf_54_u_dsync.out_clk ),
    .D(_0035_),
    .RESET_B(net902),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[30] ));
 sky130_fd_sc_hd__dfrtp_1 _7556_ (.CLK(\clknet_leaf_56_u_dsync.out_clk ),
    .D(_0036_),
    .RESET_B(net891),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[31] ));
 sky130_fd_sc_hd__dfrtp_1 _7557_ (.CLK(\clknet_leaf_54_u_dsync.out_clk ),
    .D(_0037_),
    .RESET_B(net904),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[32] ));
 sky130_fd_sc_hd__dfrtp_1 _7558_ (.CLK(\clknet_leaf_53_u_dsync.out_clk ),
    .D(_0038_),
    .RESET_B(net915),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[33] ));
 sky130_fd_sc_hd__dfrtp_1 _7559_ (.CLK(\clknet_leaf_51_u_dsync.out_clk ),
    .D(_0039_),
    .RESET_B(net904),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[34] ));
 sky130_fd_sc_hd__dfrtp_1 _7560_ (.CLK(\clknet_leaf_53_u_dsync.out_clk ),
    .D(_0040_),
    .RESET_B(net905),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[35] ));
 sky130_fd_sc_hd__dfrtp_1 _7561_ (.CLK(\clknet_leaf_51_u_dsync.out_clk ),
    .D(_0041_),
    .RESET_B(net915),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[36] ));
 sky130_fd_sc_hd__dfrtp_1 _7562_ (.CLK(\clknet_leaf_50_u_dsync.out_clk ),
    .D(_0042_),
    .RESET_B(net905),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[37] ));
 sky130_fd_sc_hd__dfrtp_1 _7563_ (.CLK(\clknet_leaf_53_u_dsync.out_clk ),
    .D(_0043_),
    .RESET_B(net904),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[38] ));
 sky130_fd_sc_hd__dfrtp_1 _7564_ (.CLK(\clknet_leaf_56_u_dsync.out_clk ),
    .D(_0044_),
    .RESET_B(net892),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[39] ));
 sky130_fd_sc_hd__dfrtp_1 _7565_ (.CLK(\clknet_leaf_56_u_dsync.out_clk ),
    .D(_0045_),
    .RESET_B(net891),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[40] ));
 sky130_fd_sc_hd__dfrtp_1 _7566_ (.CLK(\clknet_leaf_54_u_dsync.out_clk ),
    .D(_0046_),
    .RESET_B(net902),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[41] ));
 sky130_fd_sc_hd__dfrtp_1 _7567_ (.CLK(\clknet_leaf_56_u_dsync.out_clk ),
    .D(_0047_),
    .RESET_B(net891),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[42] ));
 sky130_fd_sc_hd__dfrtp_1 _7568_ (.CLK(\clknet_leaf_53_u_dsync.out_clk ),
    .D(_0048_),
    .RESET_B(net902),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[43] ));
 sky130_fd_sc_hd__dfrtp_1 _7569_ (.CLK(\clknet_leaf_53_u_dsync.out_clk ),
    .D(_0049_),
    .RESET_B(net915),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[44] ));
 sky130_fd_sc_hd__dfrtp_1 _7570_ (.CLK(\clknet_leaf_54_u_dsync.out_clk ),
    .D(_0050_),
    .RESET_B(net905),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[45] ));
 sky130_fd_sc_hd__dfrtp_1 _7571_ (.CLK(\clknet_leaf_57_u_dsync.out_clk ),
    .D(_0051_),
    .RESET_B(net891),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[46] ));
 sky130_fd_sc_hd__dfrtp_1 _7572_ (.CLK(\clknet_leaf_53_u_dsync.out_clk ),
    .D(_0052_),
    .RESET_B(net905),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[47] ));
 sky130_fd_sc_hd__dfrtp_1 _7573_ (.CLK(\clknet_leaf_50_u_dsync.out_clk ),
    .D(_0053_),
    .RESET_B(net904),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[48] ));
 sky130_fd_sc_hd__dfrtp_1 _7574_ (.CLK(\clknet_leaf_54_u_dsync.out_clk ),
    .D(_0054_),
    .RESET_B(net902),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[49] ));
 sky130_fd_sc_hd__dfrtp_1 _7575_ (.CLK(\clknet_leaf_32_u_dsync.out_clk ),
    .D(_0055_),
    .RESET_B(net904),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[50] ));
 sky130_fd_sc_hd__dfrtp_1 _7576_ (.CLK(\clknet_leaf_31_u_dsync.out_clk ),
    .D(_0056_),
    .RESET_B(net909),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[53] ));
 sky130_fd_sc_hd__dfrtp_1 _7577_ (.CLK(\clknet_leaf_54_u_dsync.out_clk ),
    .D(_0057_),
    .RESET_B(net903),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[54] ));
 sky130_fd_sc_hd__dfrtp_1 _7578_ (.CLK(\clknet_leaf_44_u_dsync.out_clk ),
    .D(_0058_),
    .RESET_B(net904),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[55] ));
 sky130_fd_sc_hd__dfrtp_1 _7579_ (.CLK(\clknet_leaf_56_u_dsync.out_clk ),
    .D(_0059_),
    .RESET_B(net892),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[56] ));
 sky130_fd_sc_hd__dfrtp_1 _7580_ (.CLK(\clknet_leaf_54_u_dsync.out_clk ),
    .D(_0060_),
    .RESET_B(net902),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[57] ));
 sky130_fd_sc_hd__dfrtp_1 _7581_ (.CLK(\clknet_leaf_41_u_dsync.out_clk ),
    .D(_0061_),
    .RESET_B(net891),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[58] ));
 sky130_fd_sc_hd__dfrtp_1 _7582_ (.CLK(\clknet_leaf_31_u_dsync.out_clk ),
    .D(_0062_),
    .RESET_B(net909),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[59] ));
 sky130_fd_sc_hd__dfrtp_1 _7583_ (.CLK(\clknet_leaf_33_u_dsync.out_clk ),
    .D(_0063_),
    .RESET_B(net903),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[60] ));
 sky130_fd_sc_hd__dfrtp_1 _7584_ (.CLK(\clknet_leaf_33_u_dsync.out_clk ),
    .D(net1787),
    .RESET_B(net897),
    .Q(\u_s2.u_sync_wbb.s_cmd_rd_data_l[61] ));
 sky130_fd_sc_hd__dfrtp_4 _7585_ (.CLK(\clknet_leaf_107_u_dsync.out_clk ),
    .D(_0065_),
    .RESET_B(net841),
    .Q(\u_s2.gnt[0] ));
 sky130_fd_sc_hd__dfrtp_4 _7586_ (.CLK(\clknet_leaf_107_u_dsync.out_clk ),
    .D(_0066_),
    .RESET_B(net841),
    .Q(\u_s2.gnt[1] ));
 sky130_fd_sc_hd__dfrtp_2 _7587_ (.CLK(\clknet_leaf_100_u_dsync.out_clk ),
    .D(_0067_),
    .RESET_B(net840),
    .Q(\u_s0.u_sync_wbb.m_bl_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_2 _7588_ (.CLK(\clknet_leaf_100_u_dsync.out_clk ),
    .D(_0068_),
    .RESET_B(net840),
    .Q(\u_s0.u_sync_wbb.m_bl_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_2 _7589_ (.CLK(\clknet_leaf_100_u_dsync.out_clk ),
    .D(_0069_),
    .RESET_B(net840),
    .Q(\u_s0.u_sync_wbb.m_bl_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7590_ (.CLK(\clknet_leaf_99_u_dsync.out_clk ),
    .D(_0070_),
    .RESET_B(net847),
    .Q(\u_s0.u_sync_wbb.m_bl_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_2 _7591_ (.CLK(\clknet_leaf_99_u_dsync.out_clk ),
    .D(_0071_),
    .RESET_B(net847),
    .Q(\u_s0.u_sync_wbb.m_bl_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7592_ (.CLK(\clknet_leaf_98_u_dsync.out_clk ),
    .D(_0072_),
    .RESET_B(net847),
    .Q(\u_s0.u_sync_wbb.m_bl_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7593_ (.CLK(\clknet_leaf_99_u_dsync.out_clk ),
    .D(_0073_),
    .RESET_B(net850),
    .Q(\u_s0.u_sync_wbb.m_bl_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_2 _7594_ (.CLK(\clknet_leaf_6_u_dsync.out_clk ),
    .D(_0074_),
    .RESET_B(net857),
    .Q(\u_s0.u_sync_wbb.m_bl_cnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7595_ (.CLK(\clknet_leaf_97_u_dsync.out_clk ),
    .D(_0075_),
    .RESET_B(net850),
    .Q(\u_s0.u_sync_wbb.m_bl_cnt[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7596_ (.CLK(\clknet_leaf_6_u_dsync.out_clk ),
    .D(_0076_),
    .RESET_B(net850),
    .Q(\u_s0.u_sync_wbb.m_bl_cnt[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7597_ (.CLK(\clknet_leaf_26_u_dsync.out_clk ),
    .D(_0077_),
    .RESET_B(net901),
    .Q(\u_reg.reg_5[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7598_ (.CLK(\clknet_leaf_20_u_dsync.out_clk ),
    .D(_0078_),
    .RESET_B(net895),
    .Q(\u_reg.reg_5[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7599_ (.CLK(\clknet_leaf_2_u_dsync.out_clk ),
    .D(_0079_),
    .RESET_B(net849),
    .Q(\u_reg.reg_5[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7600_ (.CLK(\clknet_leaf_3_u_dsync.out_clk ),
    .D(_0080_),
    .RESET_B(net860),
    .Q(\u_reg.reg_5[19] ));
 sky130_fd_sc_hd__dfrtp_1 _7601_ (.CLK(\clknet_leaf_18_u_dsync.out_clk ),
    .D(_0081_),
    .RESET_B(net888),
    .Q(\u_reg.reg_5[20] ));
 sky130_fd_sc_hd__dfrtp_1 _7602_ (.CLK(\clknet_leaf_18_u_dsync.out_clk ),
    .D(_0082_),
    .RESET_B(net888),
    .Q(\u_reg.reg_5[21] ));
 sky130_fd_sc_hd__dfrtp_1 _7603_ (.CLK(\clknet_leaf_2_u_dsync.out_clk ),
    .D(_0083_),
    .RESET_B(net848),
    .Q(\u_reg.reg_5[22] ));
 sky130_fd_sc_hd__dfrtp_1 _7604_ (.CLK(\clknet_leaf_2_u_dsync.out_clk ),
    .D(_0084_),
    .RESET_B(net855),
    .Q(\u_reg.reg_5[23] ));
 sky130_fd_sc_hd__dfrtp_1 _7605_ (.CLK(\clknet_leaf_1_u_dsync.out_clk ),
    .D(_0085_),
    .RESET_B(net846),
    .Q(\u_reg.reg_6[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7606_ (.CLK(\clknet_leaf_1_u_dsync.out_clk ),
    .D(_0086_),
    .RESET_B(net848),
    .Q(\u_reg.reg_6[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7607_ (.CLK(\clknet_leaf_2_u_dsync.out_clk ),
    .D(_0087_),
    .RESET_B(net849),
    .Q(\u_reg.reg_6[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7608_ (.CLK(\clknet_leaf_1_u_dsync.out_clk ),
    .D(_0088_),
    .RESET_B(net846),
    .Q(\u_reg.reg_6[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7609_ (.CLK(\clknet_leaf_14_u_dsync.out_clk ),
    .D(_0089_),
    .RESET_B(net871),
    .Q(\u_reg.reg_6[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7610_ (.CLK(\clknet_leaf_15_u_dsync.out_clk ),
    .D(_0090_),
    .RESET_B(net874),
    .Q(\u_reg.reg_6[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7611_ (.CLK(\clknet_leaf_3_u_dsync.out_clk ),
    .D(_0091_),
    .RESET_B(net858),
    .Q(\u_reg.reg_6[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7612_ (.CLK(\clknet_leaf_4_u_dsync.out_clk ),
    .D(_0092_),
    .RESET_B(net855),
    .Q(\u_reg.reg_6[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7613_ (.CLK(\clknet_leaf_13_u_dsync.out_clk ),
    .D(_0093_),
    .RESET_B(net882),
    .Q(\u_reg.reg_6[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7614_ (.CLK(\clknet_leaf_13_u_dsync.out_clk ),
    .D(_0094_),
    .RESET_B(net876),
    .Q(\u_reg.reg_6[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7615_ (.CLK(\clknet_leaf_13_u_dsync.out_clk ),
    .D(_0095_),
    .RESET_B(net876),
    .Q(\u_reg.reg_6[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7616_ (.CLK(\clknet_leaf_20_u_dsync.out_clk ),
    .D(_0096_),
    .RESET_B(net896),
    .Q(\u_reg.reg_6[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7617_ (.CLK(\clknet_leaf_13_u_dsync.out_clk ),
    .D(_0097_),
    .RESET_B(net882),
    .Q(\u_reg.reg_6[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7618_ (.CLK(\clknet_leaf_19_u_dsync.out_clk ),
    .D(_0098_),
    .RESET_B(net889),
    .Q(\u_reg.reg_6[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7619_ (.CLK(\clknet_leaf_19_u_dsync.out_clk ),
    .D(_0099_),
    .RESET_B(net889),
    .Q(\u_reg.reg_6[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7620_ (.CLK(\clknet_leaf_19_u_dsync.out_clk ),
    .D(_0100_),
    .RESET_B(net887),
    .Q(\u_reg.reg_6[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7621_ (.CLK(\clknet_leaf_26_u_dsync.out_clk ),
    .D(_0101_),
    .RESET_B(net901),
    .Q(\u_reg.reg_6[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7622_ (.CLK(\clknet_leaf_20_u_dsync.out_clk ),
    .D(_0102_),
    .RESET_B(net899),
    .Q(\u_reg.reg_6[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7623_ (.CLK(\clknet_leaf_2_u_dsync.out_clk ),
    .D(_0103_),
    .RESET_B(net854),
    .Q(\u_reg.reg_6[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7624_ (.CLK(\clknet_leaf_3_u_dsync.out_clk ),
    .D(_0104_),
    .RESET_B(net858),
    .Q(\u_reg.reg_6[19] ));
 sky130_fd_sc_hd__dfrtp_1 _7625_ (.CLK(\clknet_leaf_21_u_dsync.out_clk ),
    .D(_0105_),
    .RESET_B(net898),
    .Q(\u_reg.reg_6[20] ));
 sky130_fd_sc_hd__dfrtp_1 _7626_ (.CLK(\clknet_leaf_18_u_dsync.out_clk ),
    .D(_0106_),
    .RESET_B(net886),
    .Q(\u_reg.reg_6[21] ));
 sky130_fd_sc_hd__dfrtp_1 _7627_ (.CLK(\clknet_leaf_2_u_dsync.out_clk ),
    .D(_0107_),
    .RESET_B(net855),
    .Q(\u_reg.reg_6[22] ));
 sky130_fd_sc_hd__dfrtp_1 _7628_ (.CLK(\clknet_leaf_16_u_dsync.out_clk ),
    .D(_0108_),
    .RESET_B(net876),
    .Q(\u_reg.reg_6[23] ));
 sky130_fd_sc_hd__dfrtp_1 _7629_ (.CLK(\clknet_leaf_4_u_dsync.out_clk ),
    .D(_0109_),
    .RESET_B(net854),
    .Q(\u_reg.reg_7[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7630_ (.CLK(\clknet_leaf_1_u_dsync.out_clk ),
    .D(_0110_),
    .RESET_B(net848),
    .Q(\u_reg.reg_7[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7631_ (.CLK(\clknet_leaf_1_u_dsync.out_clk ),
    .D(_0111_),
    .RESET_B(net847),
    .Q(\u_reg.reg_7[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7632_ (.CLK(\clknet_leaf_1_u_dsync.out_clk ),
    .D(_0112_),
    .RESET_B(net846),
    .Q(\u_reg.reg_7[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7633_ (.CLK(\clknet_leaf_19_u_dsync.out_clk ),
    .D(_0113_),
    .RESET_B(net881),
    .Q(\u_reg.reg_7[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7634_ (.CLK(\clknet_leaf_17_u_dsync.out_clk ),
    .D(_0114_),
    .RESET_B(net881),
    .Q(\u_reg.reg_7[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7635_ (.CLK(\clknet_leaf_3_u_dsync.out_clk ),
    .D(_0115_),
    .RESET_B(net858),
    .Q(\u_reg.reg_7[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7636_ (.CLK(\clknet_leaf_15_u_dsync.out_clk ),
    .D(_0116_),
    .RESET_B(net868),
    .Q(\u_reg.reg_7[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7637_ (.CLK(\clknet_leaf_12_u_dsync.out_clk ),
    .D(_0117_),
    .RESET_B(net882),
    .Q(\u_reg.reg_7[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7638_ (.CLK(\clknet_leaf_25_u_dsync.out_clk ),
    .D(_0118_),
    .RESET_B(net910),
    .Q(\u_reg.reg_7[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7639_ (.CLK(\clknet_leaf_14_u_dsync.out_clk ),
    .D(_0119_),
    .RESET_B(net869),
    .Q(\u_reg.reg_7[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7640_ (.CLK(\clknet_leaf_26_u_dsync.out_clk ),
    .D(_0120_),
    .RESET_B(net898),
    .Q(\u_reg.reg_7[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7641_ (.CLK(\clknet_leaf_20_u_dsync.out_clk ),
    .D(_0121_),
    .RESET_B(net894),
    .Q(\u_reg.reg_7[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7642_ (.CLK(\clknet_leaf_12_u_dsync.out_clk ),
    .D(_0122_),
    .RESET_B(net884),
    .Q(\u_reg.reg_7[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7643_ (.CLK(\clknet_leaf_25_u_dsync.out_clk ),
    .D(_0123_),
    .RESET_B(net907),
    .Q(\u_reg.reg_7[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7644_ (.CLK(\clknet_leaf_25_u_dsync.out_clk ),
    .D(_0124_),
    .RESET_B(net912),
    .Q(\u_reg.reg_7[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7645_ (.CLK(\clknet_leaf_25_u_dsync.out_clk ),
    .D(_0125_),
    .RESET_B(net906),
    .Q(\u_reg.reg_7[16] ));
 sky130_fd_sc_hd__dfrtp_2 _7646_ (.CLK(\clknet_leaf_20_u_dsync.out_clk ),
    .D(_0126_),
    .RESET_B(net898),
    .Q(\u_reg.reg_7[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7647_ (.CLK(\clknet_leaf_16_u_dsync.out_clk ),
    .D(_0127_),
    .RESET_B(net874),
    .Q(\u_reg.reg_7[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7648_ (.CLK(\clknet_leaf_3_u_dsync.out_clk ),
    .D(_0128_),
    .RESET_B(net861),
    .Q(\u_reg.reg_7[19] ));
 sky130_fd_sc_hd__dfrtp_1 _7649_ (.CLK(\clknet_leaf_18_u_dsync.out_clk ),
    .D(_0129_),
    .RESET_B(net888),
    .Q(\u_reg.reg_7[20] ));
 sky130_fd_sc_hd__dfrtp_1 _7650_ (.CLK(\clknet_leaf_18_u_dsync.out_clk ),
    .D(_0130_),
    .RESET_B(net888),
    .Q(\u_reg.reg_7[21] ));
 sky130_fd_sc_hd__dfrtp_1 _7651_ (.CLK(\clknet_leaf_3_u_dsync.out_clk ),
    .D(_0131_),
    .RESET_B(net860),
    .Q(\u_reg.reg_7[22] ));
 sky130_fd_sc_hd__dfrtp_1 _7652_ (.CLK(\clknet_leaf_17_u_dsync.out_clk ),
    .D(_0132_),
    .RESET_B(net883),
    .Q(\u_reg.reg_7[23] ));
 sky130_fd_sc_hd__dfrtp_1 _7653_ (.CLK(\clknet_leaf_4_u_dsync.out_clk ),
    .D(_0133_),
    .RESET_B(net860),
    .Q(\u_reg.reg_5[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7654_ (.CLK(\clknet_leaf_13_u_dsync.out_clk ),
    .D(_0134_),
    .RESET_B(net871),
    .Q(\u_reg.reg_5[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7655_ (.CLK(\clknet_leaf_12_u_dsync.out_clk ),
    .D(_0135_),
    .RESET_B(net882),
    .Q(\u_reg.reg_5[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7656_ (.CLK(\clknet_leaf_26_u_dsync.out_clk ),
    .D(_0136_),
    .RESET_B(net895),
    .Q(\u_reg.reg_5[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7657_ (.CLK(\clknet_leaf_19_u_dsync.out_clk ),
    .D(_0137_),
    .RESET_B(net884),
    .Q(\u_reg.reg_5[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7658_ (.CLK(\clknet_leaf_20_u_dsync.out_clk ),
    .D(_0138_),
    .RESET_B(net894),
    .Q(\u_reg.reg_5[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7659_ (.CLK(\clknet_leaf_20_u_dsync.out_clk ),
    .D(_0139_),
    .RESET_B(net896),
    .Q(\u_reg.reg_5[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7660_ (.CLK(\clknet_leaf_12_u_dsync.out_clk ),
    .D(_0140_),
    .RESET_B(net887),
    .Q(\u_reg.reg_5[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7661_ (.CLK(\clknet_leaf_1_u_dsync.out_clk ),
    .D(_0141_),
    .RESET_B(net846),
    .Q(\u_reg.reg_5[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7662_ (.CLK(\clknet_leaf_1_u_dsync.out_clk ),
    .D(_0142_),
    .RESET_B(net848),
    .Q(\u_reg.reg_5[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7663_ (.CLK(\clknet_leaf_1_u_dsync.out_clk ),
    .D(_0143_),
    .RESET_B(net846),
    .Q(\u_reg.reg_5[2] ));
 sky130_fd_sc_hd__dfrtp_2 _7664_ (.CLK(\clknet_leaf_0_u_dsync.out_clk ),
    .D(_0144_),
    .RESET_B(net840),
    .Q(\u_reg.reg_5[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7665_ (.CLK(\clknet_leaf_15_u_dsync.out_clk ),
    .D(_0145_),
    .RESET_B(net870),
    .Q(\u_reg.reg_5[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7666_ (.CLK(\clknet_leaf_15_u_dsync.out_clk ),
    .D(_0146_),
    .RESET_B(net870),
    .Q(\u_reg.reg_5[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7667_ (.CLK(\clknet_leaf_3_u_dsync.out_clk ),
    .D(_0147_),
    .RESET_B(net855),
    .Q(\u_reg.reg_5[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7668_ (.CLK(\clknet_leaf_3_u_dsync.out_clk ),
    .D(_0148_),
    .RESET_B(net856),
    .Q(\u_reg.reg_5[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7669_ (.CLK(\clknet_leaf_20_u_dsync.out_clk ),
    .D(_0149_),
    .RESET_B(net900),
    .Q(\u_reg.reg_4[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7670_ (.CLK(\clknet_leaf_24_u_dsync.out_clk ),
    .D(_0150_),
    .RESET_B(net907),
    .Q(\u_reg.reg_4[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7671_ (.CLK(\clknet_leaf_16_u_dsync.out_clk ),
    .D(_0151_),
    .RESET_B(net874),
    .Q(\u_reg.reg_4[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7672_ (.CLK(\clknet_leaf_3_u_dsync.out_clk ),
    .D(_0152_),
    .RESET_B(net858),
    .Q(\u_reg.reg_4[19] ));
 sky130_fd_sc_hd__dfrtp_1 _7673_ (.CLK(\clknet_leaf_21_u_dsync.out_clk ),
    .D(_0153_),
    .RESET_B(net895),
    .Q(\u_reg.reg_4[20] ));
 sky130_fd_sc_hd__dfrtp_1 _7674_ (.CLK(\clknet_leaf_18_u_dsync.out_clk ),
    .D(_0154_),
    .RESET_B(net886),
    .Q(\u_reg.reg_4[21] ));
 sky130_fd_sc_hd__dfrtp_1 _7675_ (.CLK(\clknet_leaf_16_u_dsync.out_clk ),
    .D(_0155_),
    .RESET_B(net868),
    .Q(\u_reg.reg_4[22] ));
 sky130_fd_sc_hd__dfrtp_1 _7676_ (.CLK(\clknet_leaf_3_u_dsync.out_clk ),
    .D(_0156_),
    .RESET_B(net858),
    .Q(\u_reg.reg_4[23] ));
 sky130_fd_sc_hd__dfrtp_1 _7677_ (.CLK(\clknet_leaf_14_u_dsync.out_clk ),
    .D(_0157_),
    .RESET_B(net870),
    .Q(\u_reg.reg_4[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7678_ (.CLK(\clknet_leaf_28_u_dsync.out_clk ),
    .D(_0158_),
    .RESET_B(net912),
    .Q(\u_reg.reg_4[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7679_ (.CLK(\clknet_leaf_13_u_dsync.out_clk ),
    .D(_0159_),
    .RESET_B(net874),
    .Q(\u_reg.reg_4[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7680_ (.CLK(\clknet_leaf_26_u_dsync.out_clk ),
    .D(_0160_),
    .RESET_B(net899),
    .Q(\u_reg.reg_4[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7681_ (.CLK(\clknet_leaf_19_u_dsync.out_clk ),
    .D(_0161_),
    .RESET_B(net887),
    .Q(\u_reg.reg_4[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7682_ (.CLK(\clknet_leaf_12_u_dsync.out_clk ),
    .D(_0162_),
    .RESET_B(net884),
    .Q(\u_reg.reg_4[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7683_ (.CLK(\clknet_leaf_25_u_dsync.out_clk ),
    .D(_0163_),
    .RESET_B(net912),
    .Q(\u_reg.reg_4[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7684_ (.CLK(\clknet_leaf_25_u_dsync.out_clk ),
    .D(_0164_),
    .RESET_B(net908),
    .Q(\u_reg.reg_4[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7685_ (.CLK(\clknet_leaf_5_u_dsync.out_clk ),
    .D(_0165_),
    .RESET_B(net856),
    .Q(\u_reg.reg_4[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7686_ (.CLK(\clknet_leaf_5_u_dsync.out_clk ),
    .D(_0166_),
    .RESET_B(net849),
    .Q(\u_reg.reg_4[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7687_ (.CLK(\clknet_leaf_2_u_dsync.out_clk ),
    .D(_0167_),
    .RESET_B(net849),
    .Q(\u_reg.reg_4[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7688_ (.CLK(\clknet_leaf_1_u_dsync.out_clk ),
    .D(_0168_),
    .RESET_B(net849),
    .Q(\u_reg.reg_4[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7689_ (.CLK(\clknet_leaf_15_u_dsync.out_clk ),
    .D(_0169_),
    .RESET_B(net877),
    .Q(\u_reg.reg_4[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7690_ (.CLK(\clknet_leaf_16_u_dsync.out_clk ),
    .D(_0170_),
    .RESET_B(net874),
    .Q(\u_reg.reg_4[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7691_ (.CLK(\clknet_leaf_15_u_dsync.out_clk ),
    .D(_0171_),
    .RESET_B(net868),
    .Q(\u_reg.reg_4[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7692_ (.CLK(\clknet_leaf_15_u_dsync.out_clk ),
    .D(_0172_),
    .RESET_B(net877),
    .Q(\u_reg.reg_4[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7693_ (.CLK(\clknet_leaf_23_u_dsync.out_clk ),
    .D(_0173_),
    .RESET_B(net910),
    .Q(\u_reg.reg_3[24] ));
 sky130_fd_sc_hd__dfrtp_1 _7694_ (.CLK(\clknet_leaf_23_u_dsync.out_clk ),
    .D(_0174_),
    .RESET_B(net911),
    .Q(\u_reg.reg_3[25] ));
 sky130_fd_sc_hd__dfrtp_1 _7695_ (.CLK(\clknet_leaf_21_u_dsync.out_clk ),
    .D(_0175_),
    .RESET_B(net895),
    .Q(\u_reg.reg_3[26] ));
 sky130_fd_sc_hd__dfrtp_1 _7696_ (.CLK(\clknet_leaf_24_u_dsync.out_clk ),
    .D(_0176_),
    .RESET_B(net906),
    .Q(\u_reg.reg_3[27] ));
 sky130_fd_sc_hd__dfrtp_1 _7697_ (.CLK(\clknet_leaf_18_u_dsync.out_clk ),
    .D(_0177_),
    .RESET_B(net888),
    .Q(\u_reg.reg_3[28] ));
 sky130_fd_sc_hd__dfrtp_1 _7698_ (.CLK(\clknet_leaf_22_u_dsync.out_clk ),
    .D(_0178_),
    .RESET_B(net900),
    .Q(\u_reg.reg_3[29] ));
 sky130_fd_sc_hd__dfrtp_1 _7699_ (.CLK(\clknet_leaf_23_u_dsync.out_clk ),
    .D(_0179_),
    .RESET_B(net910),
    .Q(\u_reg.reg_3[30] ));
 sky130_fd_sc_hd__dfrtp_1 _7700_ (.CLK(\clknet_leaf_17_u_dsync.out_clk ),
    .D(_0180_),
    .RESET_B(net883),
    .Q(\u_reg.reg_3[31] ));
 sky130_fd_sc_hd__dfrtp_1 _7701_ (.CLK(\clknet_leaf_14_u_dsync.out_clk ),
    .D(_0181_),
    .RESET_B(net875),
    .Q(\u_reg.reg_3[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7702_ (.CLK(\clknet_leaf_24_u_dsync.out_clk ),
    .D(_0182_),
    .RESET_B(net911),
    .Q(\u_reg.reg_3[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7703_ (.CLK(\clknet_leaf_14_u_dsync.out_clk ),
    .D(_0183_),
    .RESET_B(net871),
    .Q(\u_reg.reg_3[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7704_ (.CLK(\clknet_leaf_26_u_dsync.out_clk ),
    .D(_0184_),
    .RESET_B(net901),
    .Q(\u_reg.reg_3[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7705_ (.CLK(\clknet_leaf_20_u_dsync.out_clk ),
    .D(_0185_),
    .RESET_B(net895),
    .Q(\u_reg.reg_3[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7706_ (.CLK(\clknet_leaf_19_u_dsync.out_clk ),
    .D(_0186_),
    .RESET_B(net887),
    .Q(\u_reg.reg_3[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7707_ (.CLK(\clknet_leaf_25_u_dsync.out_clk ),
    .D(_0187_),
    .RESET_B(net906),
    .Q(\u_reg.reg_3[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7708_ (.CLK(\clknet_leaf_24_u_dsync.out_clk ),
    .D(_0188_),
    .RESET_B(net912),
    .Q(\u_reg.reg_3[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7709_ (.CLK(\clknet_leaf_5_u_dsync.out_clk ),
    .D(_0189_),
    .RESET_B(net856),
    .Q(\u_reg.reg_3[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7710_ (.CLK(\clknet_leaf_2_u_dsync.out_clk ),
    .D(_0190_),
    .RESET_B(net854),
    .Q(\u_reg.reg_3[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7711_ (.CLK(\clknet_leaf_2_u_dsync.out_clk ),
    .D(_0191_),
    .RESET_B(net854),
    .Q(\u_reg.reg_3[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7712_ (.CLK(\clknet_leaf_4_u_dsync.out_clk ),
    .D(_0192_),
    .RESET_B(net854),
    .Q(\u_reg.reg_3[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7713_ (.CLK(\clknet_leaf_18_u_dsync.out_clk ),
    .D(_0193_),
    .RESET_B(net881),
    .Q(\u_reg.reg_3[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7714_ (.CLK(\clknet_leaf_17_u_dsync.out_clk ),
    .D(_0194_),
    .RESET_B(net881),
    .Q(\u_reg.reg_3[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7715_ (.CLK(\clknet_leaf_3_u_dsync.out_clk ),
    .D(_0195_),
    .RESET_B(net858),
    .Q(\u_reg.reg_3[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7716_ (.CLK(\clknet_leaf_15_u_dsync.out_clk ),
    .D(_0196_),
    .RESET_B(net868),
    .Q(\u_reg.reg_3[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7717_ (.CLK(\clknet_leaf_13_u_dsync.out_clk ),
    .D(_0197_),
    .RESET_B(net882),
    .Q(\u_reg.reg_2[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7718_ (.CLK(\clknet_leaf_10_u_dsync.out_clk ),
    .D(_0198_),
    .RESET_B(net875),
    .Q(\u_reg.reg_2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7719_ (.CLK(\clknet_leaf_13_u_dsync.out_clk ),
    .D(_0199_),
    .RESET_B(net876),
    .Q(\u_reg.reg_2[10] ));
 sky130_fd_sc_hd__dfrtp_2 _7720_ (.CLK(\clknet_leaf_12_u_dsync.out_clk ),
    .D(_0200_),
    .RESET_B(net882),
    .Q(\u_reg.reg_2[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7721_ (.CLK(\clknet_leaf_19_u_dsync.out_clk ),
    .D(_0201_),
    .RESET_B(net883),
    .Q(\u_reg.reg_2[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7722_ (.CLK(\clknet_leaf_12_u_dsync.out_clk ),
    .D(_0202_),
    .RESET_B(net888),
    .Q(\u_reg.reg_2[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7723_ (.CLK(\clknet_leaf_19_u_dsync.out_clk ),
    .D(_0203_),
    .RESET_B(net886),
    .Q(\u_reg.reg_2[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7724_ (.CLK(\clknet_leaf_19_u_dsync.out_clk ),
    .D(_0204_),
    .RESET_B(net887),
    .Q(\u_reg.reg_2[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7725_ (.CLK(\clknet_leaf_24_u_dsync.out_clk ),
    .D(_0205_),
    .RESET_B(net907),
    .Q(\u_reg.reg_2[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7726_ (.CLK(\clknet_leaf_24_u_dsync.out_clk ),
    .D(_0206_),
    .RESET_B(net910),
    .Q(\u_reg.reg_2[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7727_ (.CLK(\clknet_leaf_16_u_dsync.out_clk ),
    .D(_0207_),
    .RESET_B(net870),
    .Q(\u_reg.reg_2[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7728_ (.CLK(\clknet_leaf_3_u_dsync.out_clk ),
    .D(_0208_),
    .RESET_B(net858),
    .Q(\u_reg.reg_2[19] ));
 sky130_fd_sc_hd__dfrtp_1 _7729_ (.CLK(\clknet_leaf_21_u_dsync.out_clk ),
    .D(_0209_),
    .RESET_B(net899),
    .Q(\u_reg.reg_2[20] ));
 sky130_fd_sc_hd__dfrtp_1 _7730_ (.CLK(\clknet_leaf_19_u_dsync.out_clk ),
    .D(_0210_),
    .RESET_B(net883),
    .Q(\u_reg.reg_2[21] ));
 sky130_fd_sc_hd__dfrtp_1 _7731_ (.CLK(\clknet_leaf_16_u_dsync.out_clk ),
    .D(_0211_),
    .RESET_B(net868),
    .Q(\u_reg.reg_2[22] ));
 sky130_fd_sc_hd__dfrtp_1 _7732_ (.CLK(\clknet_leaf_17_u_dsync.out_clk ),
    .D(_0212_),
    .RESET_B(net883),
    .Q(\u_reg.reg_2[23] ));
 sky130_fd_sc_hd__dfrtp_1 _7733_ (.CLK(\clknet_leaf_23_u_dsync.out_clk ),
    .D(_0213_),
    .RESET_B(net910),
    .Q(\u_reg.reg_2[24] ));
 sky130_fd_sc_hd__dfrtp_1 _7734_ (.CLK(\clknet_leaf_23_u_dsync.out_clk ),
    .D(_0214_),
    .RESET_B(net910),
    .Q(\u_reg.reg_2[25] ));
 sky130_fd_sc_hd__dfrtp_1 _7735_ (.CLK(\clknet_leaf_21_u_dsync.out_clk ),
    .D(_0215_),
    .RESET_B(net895),
    .Q(\u_reg.reg_2[26] ));
 sky130_fd_sc_hd__dfrtp_1 _7736_ (.CLK(\clknet_leaf_23_u_dsync.out_clk ),
    .D(_0216_),
    .RESET_B(net911),
    .Q(\u_reg.reg_2[27] ));
 sky130_fd_sc_hd__dfrtp_1 _7737_ (.CLK(\clknet_leaf_18_u_dsync.out_clk ),
    .D(_0217_),
    .RESET_B(net888),
    .Q(\u_reg.reg_2[28] ));
 sky130_fd_sc_hd__dfrtp_1 _7738_ (.CLK(\clknet_leaf_21_u_dsync.out_clk ),
    .D(_0218_),
    .RESET_B(net898),
    .Q(\u_reg.reg_2[29] ));
 sky130_fd_sc_hd__dfrtp_1 _7739_ (.CLK(\clknet_leaf_23_u_dsync.out_clk ),
    .D(_0219_),
    .RESET_B(net911),
    .Q(\u_reg.reg_2[30] ));
 sky130_fd_sc_hd__dfrtp_1 _7740_ (.CLK(\clknet_leaf_18_u_dsync.out_clk ),
    .D(_0220_),
    .RESET_B(net888),
    .Q(\u_reg.reg_2[31] ));
 sky130_fd_sc_hd__dfrtp_2 _7741_ (.CLK(\clknet_leaf_13_u_dsync.out_clk ),
    .D(_0221_),
    .RESET_B(net882),
    .Q(\u_dcg_riscv.cfg_mode[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7742_ (.CLK(\clknet_leaf_25_u_dsync.out_clk ),
    .D(_0222_),
    .RESET_B(net908),
    .Q(\u_dcg_riscv.cfg_mode[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7743_ (.CLK(\clknet_leaf_13_u_dsync.out_clk ),
    .D(_0223_),
    .RESET_B(net875),
    .Q(\u_reg.cfg_dcg_ctrl[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7744_ (.CLK(\clknet_leaf_26_u_dsync.out_clk ),
    .D(_0224_),
    .RESET_B(net899),
    .Q(\u_reg.cfg_dcg_ctrl[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7745_ (.CLK(\clknet_leaf_19_u_dsync.out_clk ),
    .D(_0225_),
    .RESET_B(net889),
    .Q(\u_reg.cfg_dcg_ctrl[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7746_ (.CLK(\clknet_leaf_12_u_dsync.out_clk ),
    .D(_0226_),
    .RESET_B(net883),
    .Q(\u_reg.cfg_dcg_ctrl[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7747_ (.CLK(\clknet_leaf_25_u_dsync.out_clk ),
    .D(_0227_),
    .RESET_B(net906),
    .Q(\u_reg.cfg_dcg_ctrl[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7748_ (.CLK(\clknet_leaf_26_u_dsync.out_clk ),
    .D(_0228_),
    .RESET_B(net900),
    .Q(\u_reg.cfg_dcg_ctrl[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7749_ (.CLK(\clknet_leaf_20_u_dsync.out_clk ),
    .D(_0229_),
    .RESET_B(net899),
    .Q(\u_reg.cfg_dcg_ctrl[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7750_ (.CLK(\clknet_leaf_20_u_dsync.out_clk ),
    .D(_0230_),
    .RESET_B(net895),
    .Q(\u_reg.cfg_dcg_ctrl[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7751_ (.CLK(\clknet_leaf_2_u_dsync.out_clk ),
    .D(_0231_),
    .RESET_B(net854),
    .Q(\u_reg.cfg_dcg_ctrl[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7752_ (.CLK(\clknet_leaf_3_u_dsync.out_clk ),
    .D(_0232_),
    .RESET_B(net858),
    .Q(\u_reg.cfg_dcg_ctrl[19] ));
 sky130_fd_sc_hd__dfrtp_1 _7753_ (.CLK(\clknet_leaf_21_u_dsync.out_clk ),
    .D(_0233_),
    .RESET_B(net894),
    .Q(\u_reg.cfg_dcg_ctrl[20] ));
 sky130_fd_sc_hd__dfrtp_1 _7754_ (.CLK(\clknet_leaf_18_u_dsync.out_clk ),
    .D(_0234_),
    .RESET_B(net886),
    .Q(\u_reg.cfg_dcg_ctrl[21] ));
 sky130_fd_sc_hd__dfrtp_1 _7755_ (.CLK(\clknet_leaf_3_u_dsync.out_clk ),
    .D(_0235_),
    .RESET_B(net855),
    .Q(\u_reg.cfg_dcg_ctrl[22] ));
 sky130_fd_sc_hd__dfrtp_1 _7756_ (.CLK(\clknet_leaf_2_u_dsync.out_clk ),
    .D(_0236_),
    .RESET_B(net854),
    .Q(\u_reg.cfg_dcg_ctrl[23] ));
 sky130_fd_sc_hd__dfrtp_1 _7757_ (.CLK(\clknet_leaf_22_u_dsync.out_clk ),
    .D(_0237_),
    .RESET_B(net906),
    .Q(\u_reg.cfg_dcg_ctrl[24] ));
 sky130_fd_sc_hd__dfrtp_1 _7758_ (.CLK(\clknet_leaf_22_u_dsync.out_clk ),
    .D(_0238_),
    .RESET_B(net910),
    .Q(\u_reg.cfg_dcg_ctrl[25] ));
 sky130_fd_sc_hd__dfrtp_1 _7759_ (.CLK(\clknet_leaf_18_u_dsync.out_clk ),
    .D(_0239_),
    .RESET_B(net886),
    .Q(\u_reg.cfg_dcg_ctrl[26] ));
 sky130_fd_sc_hd__dfrtp_1 _7760_ (.CLK(\clknet_leaf_23_u_dsync.out_clk ),
    .D(_0240_),
    .RESET_B(net907),
    .Q(\u_reg.cfg_dcg_ctrl[27] ));
 sky130_fd_sc_hd__dfrtp_1 _7761_ (.CLK(\clknet_leaf_17_u_dsync.out_clk ),
    .D(_0241_),
    .RESET_B(net881),
    .Q(\u_reg.cfg_dcg_ctrl[28] ));
 sky130_fd_sc_hd__dfrtp_1 _7762_ (.CLK(\clknet_leaf_21_u_dsync.out_clk ),
    .D(_0242_),
    .RESET_B(net900),
    .Q(\u_reg.cfg_dcg_ctrl[29] ));
 sky130_fd_sc_hd__dfrtp_1 _7763_ (.CLK(\clknet_leaf_22_u_dsync.out_clk ),
    .D(_0243_),
    .RESET_B(net906),
    .Q(\u_reg.cfg_dcg_ctrl[30] ));
 sky130_fd_sc_hd__dfrtp_1 _7764_ (.CLK(\clknet_leaf_16_u_dsync.out_clk ),
    .D(_0244_),
    .RESET_B(net876),
    .Q(\u_reg.cfg_dcg_ctrl[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7765_ (.CLK(\clknet_leaf_42_u_dsync.out_clk ),
    .D(_0245_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7766_ (.CLK(\clknet_leaf_52_u_dsync.out_clk ),
    .D(_0246_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7767_ (.CLK(\clknet_leaf_51_u_dsync.out_clk ),
    .D(_0247_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7768_ (.CLK(\clknet_leaf_53_u_dsync.out_clk ),
    .D(_0248_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7769_ (.CLK(\clknet_leaf_48_u_dsync.out_clk ),
    .D(_0249_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7770_ (.CLK(\clknet_leaf_48_u_dsync.out_clk ),
    .D(_0250_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7771_ (.CLK(\clknet_leaf_48_u_dsync.out_clk ),
    .D(_0251_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7772_ (.CLK(\clknet_leaf_60_u_dsync.out_clk ),
    .D(_0252_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7773_ (.CLK(\clknet_leaf_49_u_dsync.out_clk ),
    .D(_0253_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7774_ (.CLK(\clknet_leaf_50_u_dsync.out_clk ),
    .D(_0254_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7775_ (.CLK(\clknet_leaf_48_u_dsync.out_clk ),
    .D(_0255_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7776_ (.CLK(\clknet_leaf_62_u_dsync.out_clk ),
    .D(_0256_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7777_ (.CLK(\clknet_leaf_51_u_dsync.out_clk ),
    .D(_0257_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7778_ (.CLK(\clknet_leaf_56_u_dsync.out_clk ),
    .D(_0258_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7779_ (.CLK(\clknet_leaf_55_u_dsync.out_clk ),
    .D(_0259_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7780_ (.CLK(\clknet_leaf_50_u_dsync.out_clk ),
    .D(_0260_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7781_ (.CLK(\clknet_leaf_55_u_dsync.out_clk ),
    .D(_0261_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7782_ (.CLK(\clknet_leaf_51_u_dsync.out_clk ),
    .D(_0262_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7783_ (.CLK(\clknet_leaf_51_u_dsync.out_clk ),
    .D(_0263_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7784_ (.CLK(\clknet_leaf_50_u_dsync.out_clk ),
    .D(_0264_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7785_ (.CLK(\clknet_leaf_50_u_dsync.out_clk ),
    .D(_0265_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7786_ (.CLK(\clknet_leaf_55_u_dsync.out_clk ),
    .D(_0266_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7787_ (.CLK(\clknet_leaf_55_u_dsync.out_clk ),
    .D(_0267_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7788_ (.CLK(\clknet_leaf_50_u_dsync.out_clk ),
    .D(_0268_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7789_ (.CLK(\clknet_leaf_62_u_dsync.out_clk ),
    .D(_0269_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7790_ (.CLK(\clknet_leaf_62_u_dsync.out_clk ),
    .D(_0270_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7791_ (.CLK(\clknet_leaf_63_u_dsync.out_clk ),
    .D(_0271_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7792_ (.CLK(\clknet_leaf_54_u_dsync.out_clk ),
    .D(_0272_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7793_ (.CLK(\clknet_leaf_63_u_dsync.out_clk ),
    .D(_0273_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7794_ (.CLK(\clknet_leaf_60_u_dsync.out_clk ),
    .D(_0274_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7795_ (.CLK(\clknet_leaf_61_u_dsync.out_clk ),
    .D(_0275_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7796_ (.CLK(\clknet_leaf_62_u_dsync.out_clk ),
    .D(_0276_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7797_ (.CLK(\clknet_leaf_42_u_dsync.out_clk ),
    .D(_0277_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7798_ (.CLK(\clknet_leaf_52_u_dsync.out_clk ),
    .D(_0278_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7799_ (.CLK(\clknet_leaf_51_u_dsync.out_clk ),
    .D(_0279_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7800_ (.CLK(\clknet_leaf_52_u_dsync.out_clk ),
    .D(_0280_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7801_ (.CLK(\clknet_leaf_48_u_dsync.out_clk ),
    .D(_0281_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7802_ (.CLK(\clknet_leaf_48_u_dsync.out_clk ),
    .D(_0282_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7803_ (.CLK(\clknet_leaf_48_u_dsync.out_clk ),
    .D(_0283_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7804_ (.CLK(\clknet_leaf_61_u_dsync.out_clk ),
    .D(_0284_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7805_ (.CLK(\clknet_leaf_50_u_dsync.out_clk ),
    .D(_0285_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7806_ (.CLK(\clknet_leaf_54_u_dsync.out_clk ),
    .D(_0286_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7807_ (.CLK(\clknet_leaf_48_u_dsync.out_clk ),
    .D(_0287_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7808_ (.CLK(\clknet_leaf_62_u_dsync.out_clk ),
    .D(_0288_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7809_ (.CLK(\clknet_leaf_49_u_dsync.out_clk ),
    .D(_0289_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7810_ (.CLK(\clknet_leaf_62_u_dsync.out_clk ),
    .D(_0290_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7811_ (.CLK(\clknet_leaf_55_u_dsync.out_clk ),
    .D(_0291_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7812_ (.CLK(\clknet_leaf_50_u_dsync.out_clk ),
    .D(_0292_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7813_ (.CLK(\clknet_leaf_54_u_dsync.out_clk ),
    .D(_0293_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7814_ (.CLK(\clknet_leaf_52_u_dsync.out_clk ),
    .D(_0294_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7815_ (.CLK(\clknet_leaf_51_u_dsync.out_clk ),
    .D(_0295_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7816_ (.CLK(\clknet_leaf_42_u_dsync.out_clk ),
    .D(_0296_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7817_ (.CLK(\clknet_leaf_49_u_dsync.out_clk ),
    .D(_0297_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7818_ (.CLK(\clknet_leaf_63_u_dsync.out_clk ),
    .D(_0298_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7819_ (.CLK(\clknet_leaf_42_u_dsync.out_clk ),
    .D(_0299_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7820_ (.CLK(\clknet_leaf_50_u_dsync.out_clk ),
    .D(_0300_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7821_ (.CLK(\clknet_leaf_63_u_dsync.out_clk ),
    .D(_0301_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7822_ (.CLK(\clknet_leaf_62_u_dsync.out_clk ),
    .D(_0302_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7823_ (.CLK(\clknet_leaf_63_u_dsync.out_clk ),
    .D(_0303_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7824_ (.CLK(\clknet_leaf_54_u_dsync.out_clk ),
    .D(_0304_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7825_ (.CLK(\clknet_leaf_63_u_dsync.out_clk ),
    .D(_0305_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7826_ (.CLK(\clknet_leaf_61_u_dsync.out_clk ),
    .D(_0306_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7827_ (.CLK(\clknet_leaf_62_u_dsync.out_clk ),
    .D(_0307_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7828_ (.CLK(\clknet_leaf_61_u_dsync.out_clk ),
    .D(_0308_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7829_ (.CLK(\clknet_leaf_42_u_dsync.out_clk ),
    .D(_0309_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7830_ (.CLK(\clknet_leaf_52_u_dsync.out_clk ),
    .D(_0310_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7831_ (.CLK(\clknet_leaf_52_u_dsync.out_clk ),
    .D(_0311_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7832_ (.CLK(\clknet_leaf_52_u_dsync.out_clk ),
    .D(_0312_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7833_ (.CLK(\clknet_leaf_47_u_dsync.out_clk ),
    .D(net1780),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7834_ (.CLK(\clknet_leaf_48_u_dsync.out_clk ),
    .D(_0314_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7835_ (.CLK(\clknet_leaf_48_u_dsync.out_clk ),
    .D(_0315_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7836_ (.CLK(\clknet_leaf_62_u_dsync.out_clk ),
    .D(_0316_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7837_ (.CLK(\clknet_leaf_50_u_dsync.out_clk ),
    .D(_0317_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7838_ (.CLK(\clknet_leaf_50_u_dsync.out_clk ),
    .D(_0318_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7839_ (.CLK(\clknet_leaf_47_u_dsync.out_clk ),
    .D(_0319_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7840_ (.CLK(\clknet_leaf_55_u_dsync.out_clk ),
    .D(_0320_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7841_ (.CLK(\clknet_leaf_48_u_dsync.out_clk ),
    .D(_0321_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7842_ (.CLK(\clknet_leaf_62_u_dsync.out_clk ),
    .D(_0322_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7843_ (.CLK(\clknet_leaf_55_u_dsync.out_clk ),
    .D(_0323_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7844_ (.CLK(\clknet_leaf_49_u_dsync.out_clk ),
    .D(_0324_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7845_ (.CLK(\clknet_leaf_50_u_dsync.out_clk ),
    .D(_0325_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7846_ (.CLK(\clknet_leaf_52_u_dsync.out_clk ),
    .D(_0326_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7847_ (.CLK(\clknet_leaf_51_u_dsync.out_clk ),
    .D(_0327_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7848_ (.CLK(\clknet_leaf_49_u_dsync.out_clk ),
    .D(_0328_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7849_ (.CLK(\clknet_leaf_49_u_dsync.out_clk ),
    .D(_0329_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7850_ (.CLK(\clknet_leaf_63_u_dsync.out_clk ),
    .D(_0330_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7851_ (.CLK(\clknet_leaf_42_u_dsync.out_clk ),
    .D(_0331_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7852_ (.CLK(\clknet_leaf_50_u_dsync.out_clk ),
    .D(_0332_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7853_ (.CLK(\clknet_leaf_63_u_dsync.out_clk ),
    .D(_0333_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7854_ (.CLK(\clknet_leaf_63_u_dsync.out_clk ),
    .D(_0334_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7855_ (.CLK(\clknet_leaf_64_u_dsync.out_clk ),
    .D(_0335_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7856_ (.CLK(\clknet_leaf_55_u_dsync.out_clk ),
    .D(_0336_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7857_ (.CLK(\clknet_leaf_41_u_dsync.out_clk ),
    .D(_0337_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7858_ (.CLK(\clknet_leaf_60_u_dsync.out_clk ),
    .D(_0338_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7859_ (.CLK(\clknet_leaf_62_u_dsync.out_clk ),
    .D(_0339_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7860_ (.CLK(\clknet_leaf_61_u_dsync.out_clk ),
    .D(_0340_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7861_ (.CLK(\clknet_leaf_42_u_dsync.out_clk ),
    .D(_0341_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7862_ (.CLK(\clknet_leaf_52_u_dsync.out_clk ),
    .D(_0342_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7863_ (.CLK(\clknet_leaf_51_u_dsync.out_clk ),
    .D(_0343_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7864_ (.CLK(\clknet_leaf_54_u_dsync.out_clk ),
    .D(_0344_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7865_ (.CLK(\clknet_leaf_48_u_dsync.out_clk ),
    .D(_0345_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7866_ (.CLK(\clknet_leaf_48_u_dsync.out_clk ),
    .D(_0346_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7867_ (.CLK(\clknet_leaf_49_u_dsync.out_clk ),
    .D(_0347_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7868_ (.CLK(\clknet_leaf_61_u_dsync.out_clk ),
    .D(_0348_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7869_ (.CLK(\clknet_leaf_49_u_dsync.out_clk ),
    .D(_0349_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7870_ (.CLK(\clknet_leaf_54_u_dsync.out_clk ),
    .D(_0350_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7871_ (.CLK(\clknet_leaf_47_u_dsync.out_clk ),
    .D(net1782),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7872_ (.CLK(\clknet_leaf_62_u_dsync.out_clk ),
    .D(_0352_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7873_ (.CLK(\clknet_leaf_48_u_dsync.out_clk ),
    .D(_0353_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7874_ (.CLK(\clknet_leaf_55_u_dsync.out_clk ),
    .D(_0354_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7875_ (.CLK(\clknet_leaf_55_u_dsync.out_clk ),
    .D(_0355_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7876_ (.CLK(\clknet_leaf_55_u_dsync.out_clk ),
    .D(_0356_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7877_ (.CLK(\clknet_leaf_55_u_dsync.out_clk ),
    .D(_0357_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7878_ (.CLK(\clknet_leaf_52_u_dsync.out_clk ),
    .D(_0358_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7879_ (.CLK(\clknet_leaf_50_u_dsync.out_clk ),
    .D(_0359_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7880_ (.CLK(\clknet_leaf_42_u_dsync.out_clk ),
    .D(_0360_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7881_ (.CLK(\clknet_leaf_49_u_dsync.out_clk ),
    .D(_0361_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7882_ (.CLK(\clknet_leaf_55_u_dsync.out_clk ),
    .D(_0362_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7883_ (.CLK(\clknet_leaf_42_u_dsync.out_clk ),
    .D(_0363_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7884_ (.CLK(\clknet_leaf_54_u_dsync.out_clk ),
    .D(_0364_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7885_ (.CLK(\clknet_leaf_63_u_dsync.out_clk ),
    .D(_0365_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7886_ (.CLK(\clknet_leaf_62_u_dsync.out_clk ),
    .D(_0366_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7887_ (.CLK(\clknet_leaf_64_u_dsync.out_clk ),
    .D(_0367_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7888_ (.CLK(\clknet_leaf_54_u_dsync.out_clk ),
    .D(_0368_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7889_ (.CLK(\clknet_leaf_41_u_dsync.out_clk ),
    .D(_0369_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7890_ (.CLK(\clknet_leaf_61_u_dsync.out_clk ),
    .D(_0370_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7891_ (.CLK(\clknet_leaf_61_u_dsync.out_clk ),
    .D(_0371_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7892_ (.CLK(\clknet_leaf_61_u_dsync.out_clk ),
    .D(_0372_),
    .Q(\u_s2.u_sync_wbb.u_resp_if.mem[3][31] ));
 sky130_fd_sc_hd__dfrtp_1 _7893_ (.CLK(\clknet_leaf_9_u_dsync.out_clk ),
    .D(_0373_),
    .RESET_B(net878),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7894_ (.CLK(\clknet_leaf_9_u_dsync.out_clk ),
    .D(_0374_),
    .RESET_B(net873),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7895_ (.CLK(\clknet_leaf_9_u_dsync.out_clk ),
    .D(_0375_),
    .RESET_B(net878),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7896_ (.CLK(\clknet_leaf_9_u_dsync.out_clk ),
    .D(_0376_),
    .RESET_B(net872),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7897_ (.CLK(\clknet_leaf_10_u_dsync.out_clk ),
    .D(_0377_),
    .RESET_B(net872),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7898_ (.CLK(\clknet_leaf_10_u_dsync.out_clk ),
    .D(_0378_),
    .RESET_B(net873),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7899_ (.CLK(\clknet_leaf_10_u_dsync.out_clk ),
    .D(_0379_),
    .RESET_B(net872),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7900_ (.CLK(\clknet_leaf_10_u_dsync.out_clk ),
    .D(_0380_),
    .RESET_B(net873),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7901_ (.CLK(\clknet_leaf_9_u_dsync.out_clk ),
    .D(_0381_),
    .RESET_B(net872),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7902_ (.CLK(\clknet_leaf_38_u_dsync.out_clk ),
    .D(_0382_),
    .RESET_B(net879),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7903_ (.CLK(\clknet_leaf_96_u_dsync.out_clk ),
    .D(_0383_),
    .RESET_B(net862),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7904_ (.CLK(\clknet_leaf_9_u_dsync.out_clk ),
    .D(_0384_),
    .RESET_B(net872),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7905_ (.CLK(\clknet_leaf_38_u_dsync.out_clk ),
    .D(_0385_),
    .RESET_B(net879),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7906_ (.CLK(\clknet_leaf_68_u_dsync.out_clk ),
    .D(_0386_),
    .RESET_B(net865),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7907_ (.CLK(\clknet_leaf_72_u_dsync.out_clk ),
    .D(_0387_),
    .RESET_B(net864),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[19] ));
 sky130_fd_sc_hd__dfrtp_1 _7908_ (.CLK(\clknet_leaf_64_u_dsync.out_clk ),
    .D(_0388_),
    .RESET_B(net880),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[20] ));
 sky130_fd_sc_hd__dfrtp_1 _7909_ (.CLK(\clknet_leaf_64_u_dsync.out_clk ),
    .D(_0389_),
    .RESET_B(net880),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[21] ));
 sky130_fd_sc_hd__dfrtp_1 _7910_ (.CLK(\clknet_leaf_64_u_dsync.out_clk ),
    .D(_0390_),
    .RESET_B(net879),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[22] ));
 sky130_fd_sc_hd__dfrtp_1 _7911_ (.CLK(\clknet_leaf_68_u_dsync.out_clk ),
    .D(_0391_),
    .RESET_B(net863),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[23] ));
 sky130_fd_sc_hd__dfrtp_1 _7912_ (.CLK(\clknet_leaf_72_u_dsync.out_clk ),
    .D(_0392_),
    .RESET_B(net864),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[24] ));
 sky130_fd_sc_hd__dfrtp_1 _7913_ (.CLK(\clknet_leaf_64_u_dsync.out_clk ),
    .D(_0393_),
    .RESET_B(net880),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[25] ));
 sky130_fd_sc_hd__dfrtp_1 _7914_ (.CLK(\clknet_leaf_64_u_dsync.out_clk ),
    .D(_0394_),
    .RESET_B(net879),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[26] ));
 sky130_fd_sc_hd__dfrtp_1 _7915_ (.CLK(\clknet_leaf_64_u_dsync.out_clk ),
    .D(_0395_),
    .RESET_B(net879),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[27] ));
 sky130_fd_sc_hd__dfrtp_1 _7916_ (.CLK(\clknet_leaf_64_u_dsync.out_clk ),
    .D(_0396_),
    .RESET_B(net880),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[28] ));
 sky130_fd_sc_hd__dfrtp_1 _7917_ (.CLK(\clknet_leaf_61_u_dsync.out_clk ),
    .D(_0397_),
    .RESET_B(net880),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[29] ));
 sky130_fd_sc_hd__dfrtp_1 _7918_ (.CLK(\clknet_leaf_63_u_dsync.out_clk ),
    .D(_0398_),
    .RESET_B(net891),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[30] ));
 sky130_fd_sc_hd__dfrtp_1 _7919_ (.CLK(\clknet_leaf_68_u_dsync.out_clk ),
    .D(_0399_),
    .RESET_B(net863),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[31] ));
 sky130_fd_sc_hd__dfrtp_1 _7920_ (.CLK(\clknet_leaf_68_u_dsync.out_clk ),
    .D(_0400_),
    .RESET_B(net863),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[32] ));
 sky130_fd_sc_hd__dfrtp_1 _7921_ (.CLK(\clknet_leaf_71_u_dsync.out_clk ),
    .D(_0401_),
    .RESET_B(net865),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[33] ));
 sky130_fd_sc_hd__dfrtp_1 _7922_ (.CLK(\clknet_leaf_67_u_dsync.out_clk ),
    .D(_0402_),
    .RESET_B(net863),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[34] ));
 sky130_fd_sc_hd__dfrtp_1 _7923_ (.CLK(\clknet_leaf_61_u_dsync.out_clk ),
    .D(_0403_),
    .RESET_B(net879),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[35] ));
 sky130_fd_sc_hd__dfrtp_1 _7924_ (.CLK(\clknet_leaf_68_u_dsync.out_clk ),
    .D(_0404_),
    .RESET_B(net865),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[36] ));
 sky130_fd_sc_hd__dfrtp_1 _7925_ (.CLK(\clknet_leaf_71_u_dsync.out_clk ),
    .D(_0405_),
    .RESET_B(net862),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[37] ));
 sky130_fd_sc_hd__dfrtp_1 _7926_ (.CLK(\clknet_leaf_61_u_dsync.out_clk ),
    .D(_0406_),
    .RESET_B(net879),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[38] ));
 sky130_fd_sc_hd__dfrtp_1 _7927_ (.CLK(\clknet_leaf_68_u_dsync.out_clk ),
    .D(_0407_),
    .RESET_B(net862),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[39] ));
 sky130_fd_sc_hd__dfrtp_1 _7928_ (.CLK(\clknet_leaf_68_u_dsync.out_clk ),
    .D(_0408_),
    .RESET_B(net862),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[40] ));
 sky130_fd_sc_hd__dfrtp_1 _7929_ (.CLK(\clknet_leaf_64_u_dsync.out_clk ),
    .D(_0409_),
    .RESET_B(net879),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[41] ));
 sky130_fd_sc_hd__dfrtp_1 _7930_ (.CLK(\clknet_leaf_71_u_dsync.out_clk ),
    .D(_0410_),
    .RESET_B(net862),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[42] ));
 sky130_fd_sc_hd__dfrtp_1 _7931_ (.CLK(\clknet_leaf_72_u_dsync.out_clk ),
    .D(_0411_),
    .RESET_B(net864),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[43] ));
 sky130_fd_sc_hd__dfrtp_1 _7932_ (.CLK(\clknet_leaf_71_u_dsync.out_clk ),
    .D(_0412_),
    .RESET_B(net865),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[44] ));
 sky130_fd_sc_hd__dfrtp_1 _7933_ (.CLK(\clknet_leaf_37_u_dsync.out_clk ),
    .D(_0413_),
    .RESET_B(net891),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[45] ));
 sky130_fd_sc_hd__dfrtp_1 _7934_ (.CLK(\clknet_leaf_60_u_dsync.out_clk ),
    .D(_0414_),
    .RESET_B(net879),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[46] ));
 sky130_fd_sc_hd__dfrtp_1 _7935_ (.CLK(\clknet_leaf_68_u_dsync.out_clk ),
    .D(_0415_),
    .RESET_B(net862),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[47] ));
 sky130_fd_sc_hd__dfrtp_1 _7936_ (.CLK(\clknet_leaf_68_u_dsync.out_clk ),
    .D(_0416_),
    .RESET_B(net864),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[48] ));
 sky130_fd_sc_hd__dfrtp_1 _7937_ (.CLK(\clknet_leaf_70_u_dsync.out_clk ),
    .D(_0417_),
    .RESET_B(net852),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[49] ));
 sky130_fd_sc_hd__dfrtp_1 _7938_ (.CLK(\clknet_leaf_66_u_dsync.out_clk ),
    .D(_0418_),
    .RESET_B(net863),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[50] ));
 sky130_fd_sc_hd__dfrtp_1 _7939_ (.CLK(\clknet_leaf_96_u_dsync.out_clk ),
    .D(_0419_),
    .RESET_B(net857),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[53] ));
 sky130_fd_sc_hd__dfrtp_1 _7940_ (.CLK(\clknet_leaf_96_u_dsync.out_clk ),
    .D(_0420_),
    .RESET_B(net863),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[54] ));
 sky130_fd_sc_hd__dfrtp_1 _7941_ (.CLK(\clknet_leaf_96_u_dsync.out_clk ),
    .D(_0421_),
    .RESET_B(net861),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[55] ));
 sky130_fd_sc_hd__dfrtp_1 _7942_ (.CLK(\clknet_leaf_96_u_dsync.out_clk ),
    .D(_0422_),
    .RESET_B(net863),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[56] ));
 sky130_fd_sc_hd__dfrtp_1 _7943_ (.CLK(\clknet_leaf_68_u_dsync.out_clk ),
    .D(_0423_),
    .RESET_B(net862),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[57] ));
 sky130_fd_sc_hd__dfrtp_1 _7944_ (.CLK(\clknet_leaf_96_u_dsync.out_clk ),
    .D(_0424_),
    .RESET_B(net863),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[58] ));
 sky130_fd_sc_hd__dfrtp_1 _7945_ (.CLK(\clknet_leaf_95_u_dsync.out_clk ),
    .D(_0425_),
    .RESET_B(net862),
    .Q(\u_s1.u_sync_wbb.s_cmd_rd_data_l[59] ));
 sky130_fd_sc_hd__dfxtp_1 _7946_ (.CLK(\clknet_leaf_7_u_dsync.out_clk ),
    .D(_0426_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7947_ (.CLK(\clknet_leaf_6_u_dsync.out_clk ),
    .D(_0427_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7948_ (.CLK(\clknet_leaf_10_u_dsync.out_clk ),
    .D(_0428_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7949_ (.CLK(\clknet_leaf_7_u_dsync.out_clk ),
    .D(_0429_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7950_ (.CLK(\clknet_leaf_11_u_dsync.out_clk ),
    .D(_0430_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7951_ (.CLK(\clknet_leaf_10_u_dsync.out_clk ),
    .D(_0431_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7952_ (.CLK(\clknet_leaf_99_u_dsync.out_clk ),
    .D(_0432_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7953_ (.CLK(\clknet_leaf_10_u_dsync.out_clk ),
    .D(_0433_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7954_ (.CLK(\clknet_leaf_6_u_dsync.out_clk ),
    .D(_0434_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7955_ (.CLK(\clknet_leaf_37_u_dsync.out_clk ),
    .D(_0435_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7956_ (.CLK(\clknet_leaf_8_u_dsync.out_clk ),
    .D(_0436_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7957_ (.CLK(\clknet_leaf_9_u_dsync.out_clk ),
    .D(_0437_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7958_ (.CLK(\clknet_leaf_9_u_dsync.out_clk ),
    .D(_0438_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7959_ (.CLK(\clknet_leaf_63_u_dsync.out_clk ),
    .D(_0439_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7960_ (.CLK(\clknet_leaf_65_u_dsync.out_clk ),
    .D(_0440_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7961_ (.CLK(\clknet_leaf_65_u_dsync.out_clk ),
    .D(_0441_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7962_ (.CLK(\clknet_leaf_66_u_dsync.out_clk ),
    .D(_0442_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7963_ (.CLK(\clknet_leaf_39_u_dsync.out_clk ),
    .D(_0443_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7964_ (.CLK(\clknet_leaf_65_u_dsync.out_clk ),
    .D(_0444_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7965_ (.CLK(\clknet_leaf_67_u_dsync.out_clk ),
    .D(_0445_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7966_ (.CLK(\clknet_leaf_39_u_dsync.out_clk ),
    .D(_0446_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7967_ (.CLK(\clknet_leaf_65_u_dsync.out_clk ),
    .D(_0447_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7968_ (.CLK(\clknet_leaf_64_u_dsync.out_clk ),
    .D(_0448_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7969_ (.CLK(\clknet_leaf_41_u_dsync.out_clk ),
    .D(_0449_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7970_ (.CLK(\clknet_leaf_39_u_dsync.out_clk ),
    .D(_0450_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7971_ (.CLK(\clknet_leaf_39_u_dsync.out_clk ),
    .D(_0451_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7972_ (.CLK(\clknet_leaf_67_u_dsync.out_clk ),
    .D(_0452_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7973_ (.CLK(\clknet_leaf_38_u_dsync.out_clk ),
    .D(_0453_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][32] ));
 sky130_fd_sc_hd__dfxtp_1 _7974_ (.CLK(\clknet_leaf_68_u_dsync.out_clk ),
    .D(_0454_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][33] ));
 sky130_fd_sc_hd__dfxtp_1 _7975_ (.CLK(\clknet_leaf_39_u_dsync.out_clk ),
    .D(_0455_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][34] ));
 sky130_fd_sc_hd__dfxtp_1 _7976_ (.CLK(\clknet_leaf_38_u_dsync.out_clk ),
    .D(_0456_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][35] ));
 sky130_fd_sc_hd__dfxtp_1 _7977_ (.CLK(\clknet_leaf_67_u_dsync.out_clk ),
    .D(_0457_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][36] ));
 sky130_fd_sc_hd__dfxtp_1 _7978_ (.CLK(\clknet_leaf_38_u_dsync.out_clk ),
    .D(_0458_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][37] ));
 sky130_fd_sc_hd__dfxtp_1 _7979_ (.CLK(\clknet_leaf_65_u_dsync.out_clk ),
    .D(_0459_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][38] ));
 sky130_fd_sc_hd__dfxtp_1 _7980_ (.CLK(\clknet_leaf_69_u_dsync.out_clk ),
    .D(_0460_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][39] ));
 sky130_fd_sc_hd__dfxtp_1 _7981_ (.CLK(\clknet_leaf_66_u_dsync.out_clk ),
    .D(_0461_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][40] ));
 sky130_fd_sc_hd__dfxtp_1 _7982_ (.CLK(\clknet_leaf_66_u_dsync.out_clk ),
    .D(_0462_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][41] ));
 sky130_fd_sc_hd__dfxtp_1 _7983_ (.CLK(\clknet_leaf_38_u_dsync.out_clk ),
    .D(_0463_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][42] ));
 sky130_fd_sc_hd__dfxtp_1 _7984_ (.CLK(\clknet_leaf_66_u_dsync.out_clk ),
    .D(_0464_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][43] ));
 sky130_fd_sc_hd__dfxtp_1 _7985_ (.CLK(\clknet_leaf_95_u_dsync.out_clk ),
    .D(_0465_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][44] ));
 sky130_fd_sc_hd__dfxtp_1 _7986_ (.CLK(\clknet_leaf_37_u_dsync.out_clk ),
    .D(_0466_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][45] ));
 sky130_fd_sc_hd__dfxtp_1 _7987_ (.CLK(\clknet_leaf_37_u_dsync.out_clk ),
    .D(_0467_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][46] ));
 sky130_fd_sc_hd__dfxtp_1 _7988_ (.CLK(\clknet_leaf_69_u_dsync.out_clk ),
    .D(_0468_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][47] ));
 sky130_fd_sc_hd__dfxtp_1 _7989_ (.CLK(\clknet_leaf_95_u_dsync.out_clk ),
    .D(_0469_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][48] ));
 sky130_fd_sc_hd__dfxtp_1 _7990_ (.CLK(\clknet_leaf_95_u_dsync.out_clk ),
    .D(_0470_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][49] ));
 sky130_fd_sc_hd__dfxtp_1 _7991_ (.CLK(\clknet_leaf_9_u_dsync.out_clk ),
    .D(_0471_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][50] ));
 sky130_fd_sc_hd__dfxtp_1 _7992_ (.CLK(\clknet_leaf_8_u_dsync.out_clk ),
    .D(_0472_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][53] ));
 sky130_fd_sc_hd__dfxtp_1 _7993_ (.CLK(\clknet_leaf_8_u_dsync.out_clk ),
    .D(_0473_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][54] ));
 sky130_fd_sc_hd__dfxtp_1 _7994_ (.CLK(\clknet_leaf_7_u_dsync.out_clk ),
    .D(_0474_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][55] ));
 sky130_fd_sc_hd__dfxtp_1 _7995_ (.CLK(\clknet_leaf_7_u_dsync.out_clk ),
    .D(_0475_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][56] ));
 sky130_fd_sc_hd__dfxtp_1 _7996_ (.CLK(\clknet_leaf_96_u_dsync.out_clk ),
    .D(_0476_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][57] ));
 sky130_fd_sc_hd__dfxtp_1 _7997_ (.CLK(\clknet_leaf_7_u_dsync.out_clk ),
    .D(_0477_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][58] ));
 sky130_fd_sc_hd__dfxtp_1 _7998_ (.CLK(\clknet_leaf_8_u_dsync.out_clk ),
    .D(_0478_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[3][59] ));
 sky130_fd_sc_hd__dfrtp_1 _7999_ (.CLK(\clknet_leaf_0_u_dsync.out_clk ),
    .D(_0479_),
    .RESET_B(net840),
    .Q(\u_s1.gnt[0] ));
 sky130_fd_sc_hd__dfrtp_2 _8000_ (.CLK(\clknet_leaf_1_u_dsync.out_clk ),
    .D(_0480_),
    .RESET_B(net846),
    .Q(\u_s1.gnt[1] ));
 sky130_fd_sc_hd__dfrtp_4 _8001_ (.CLK(\clknet_leaf_12_u_dsync.out_clk ),
    .D(_0481_),
    .RESET_B(net890),
    .Q(\u_s2.u_sync_wbb.wbm_ack_o ));
 sky130_fd_sc_hd__dfrtp_1 _8002_ (.CLK(\clknet_leaf_12_u_dsync.out_clk ),
    .D(_0482_),
    .RESET_B(net890),
    .Q(\u_s2.u_sync_wbb.wbm_lack_o ));
 sky130_fd_sc_hd__dfrtp_4 _8003_ (.CLK(\clknet_leaf_34_u_dsync.out_clk ),
    .D(net1819),
    .RESET_B(net897),
    .Q(\u_s2.u_sync_wbb.m_cmd_wr_en ));
 sky130_fd_sc_hd__dfrtp_4 _8004_ (.CLK(\clknet_leaf_28_u_dsync.out_clk ),
    .D(_0484_),
    .RESET_B(net909),
    .Q(\u_s2.u_sync_wbb.m_resp_rd_en ));
 sky130_fd_sc_hd__dfrtp_1 _8005_ (.CLK(\clknet_leaf_31_u_dsync.out_clk ),
    .D(net1499),
    .RESET_B(net909),
    .Q(\u_s2.u_sync_wbb.wbs_ack_f ));
 sky130_fd_sc_hd__dfrtp_1 _8006_ (.CLK(\clknet_leaf_31_u_dsync.out_clk ),
    .D(net438),
    .RESET_B(net913),
    .Q(\u_s2.u_sync_wbb.wbs_stb_l ));
 sky130_fd_sc_hd__dfrtp_1 _8007_ (.CLK(\clknet_leaf_49_u_dsync.out_clk ),
    .D(_0485_),
    .RESET_B(net904),
    .Q(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_4 _8008_ (.CLK(\clknet_leaf_47_u_dsync.out_clk ),
    .D(_0486_),
    .RESET_B(net915),
    .Q(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_4 _8009_ (.CLK(\clknet_leaf_46_u_dsync.out_clk ),
    .D(_0487_),
    .RESET_B(net916),
    .Q(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_4 _8010_ (.CLK(\clknet_leaf_30_u_dsync.out_clk ),
    .D(_0488_),
    .RESET_B(net914),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_2 _8011_ (.CLK(\clknet_leaf_28_u_dsync.out_clk ),
    .D(_0489_),
    .RESET_B(net909),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_4 _8012_ (.CLK(\clknet_leaf_31_u_dsync.out_clk ),
    .D(_0490_),
    .RESET_B(net913),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.wr_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8013_ (.CLK(\clknet_leaf_30_u_dsync.out_clk ),
    .D(_0491_),
    .RESET_B(net909),
    .Q(\u_s2.u_sync_wbb.wbs_burst ));
 sky130_fd_sc_hd__dfrtp_1 _8014_ (.CLK(\clknet_leaf_30_u_dsync.out_clk ),
    .D(_0492_),
    .RESET_B(net914),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_4 _8015_ (.CLK(\clknet_leaf_31_u_dsync.out_clk ),
    .D(_0493_),
    .RESET_B(net914),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_4 _8016_ (.CLK(\clknet_leaf_30_u_dsync.out_clk ),
    .D(_0494_),
    .RESET_B(net913),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.rd_ptr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8017_ (.CLK(\clknet_leaf_7_u_dsync.out_clk ),
    .D(_0495_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8018_ (.CLK(\clknet_leaf_6_u_dsync.out_clk ),
    .D(_0496_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8019_ (.CLK(\clknet_leaf_10_u_dsync.out_clk ),
    .D(_0497_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8020_ (.CLK(\clknet_leaf_7_u_dsync.out_clk ),
    .D(_0498_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8021_ (.CLK(\clknet_leaf_9_u_dsync.out_clk ),
    .D(_0499_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8022_ (.CLK(\clknet_leaf_10_u_dsync.out_clk ),
    .D(_0500_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8023_ (.CLK(\clknet_leaf_6_u_dsync.out_clk ),
    .D(_0501_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8024_ (.CLK(\clknet_leaf_7_u_dsync.out_clk ),
    .D(_0502_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8025_ (.CLK(\clknet_leaf_6_u_dsync.out_clk ),
    .D(_0503_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8026_ (.CLK(\clknet_leaf_37_u_dsync.out_clk ),
    .D(_0504_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8027_ (.CLK(\clknet_leaf_8_u_dsync.out_clk ),
    .D(_0505_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8028_ (.CLK(\clknet_leaf_9_u_dsync.out_clk ),
    .D(_0506_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8029_ (.CLK(\clknet_leaf_37_u_dsync.out_clk ),
    .D(_0507_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8030_ (.CLK(\clknet_leaf_41_u_dsync.out_clk ),
    .D(_0508_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8031_ (.CLK(\clknet_leaf_65_u_dsync.out_clk ),
    .D(_0509_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8032_ (.CLK(\clknet_leaf_65_u_dsync.out_clk ),
    .D(_0510_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8033_ (.CLK(\clknet_leaf_65_u_dsync.out_clk ),
    .D(_0511_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8034_ (.CLK(\clknet_leaf_65_u_dsync.out_clk ),
    .D(_0512_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8035_ (.CLK(\clknet_leaf_64_u_dsync.out_clk ),
    .D(_0513_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8036_ (.CLK(\clknet_leaf_67_u_dsync.out_clk ),
    .D(_0514_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8037_ (.CLK(\clknet_leaf_39_u_dsync.out_clk ),
    .D(_0515_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8038_ (.CLK(\clknet_leaf_65_u_dsync.out_clk ),
    .D(_0516_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8039_ (.CLK(\clknet_leaf_64_u_dsync.out_clk ),
    .D(_0517_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8040_ (.CLK(\clknet_leaf_41_u_dsync.out_clk ),
    .D(_0518_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8041_ (.CLK(\clknet_leaf_39_u_dsync.out_clk ),
    .D(_0519_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8042_ (.CLK(\clknet_leaf_39_u_dsync.out_clk ),
    .D(_0520_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8043_ (.CLK(\clknet_leaf_67_u_dsync.out_clk ),
    .D(_0521_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8044_ (.CLK(\clknet_leaf_38_u_dsync.out_clk ),
    .D(_0522_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _8045_ (.CLK(\clknet_leaf_68_u_dsync.out_clk ),
    .D(_0523_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _8046_ (.CLK(\clknet_leaf_65_u_dsync.out_clk ),
    .D(_0524_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _8047_ (.CLK(\clknet_leaf_37_u_dsync.out_clk ),
    .D(_0525_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _8048_ (.CLK(\clknet_leaf_67_u_dsync.out_clk ),
    .D(_0526_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _8049_ (.CLK(\clknet_leaf_38_u_dsync.out_clk ),
    .D(_0527_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _8050_ (.CLK(\clknet_leaf_65_u_dsync.out_clk ),
    .D(_0528_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _8051_ (.CLK(\clknet_leaf_69_u_dsync.out_clk ),
    .D(_0529_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _8052_ (.CLK(\clknet_leaf_67_u_dsync.out_clk ),
    .D(_0530_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _8053_ (.CLK(\clknet_leaf_67_u_dsync.out_clk ),
    .D(_0531_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _8054_ (.CLK(\clknet_leaf_38_u_dsync.out_clk ),
    .D(_0532_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _8055_ (.CLK(\clknet_leaf_66_u_dsync.out_clk ),
    .D(_0533_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _8056_ (.CLK(\clknet_leaf_95_u_dsync.out_clk ),
    .D(_0534_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _8057_ (.CLK(\clknet_leaf_37_u_dsync.out_clk ),
    .D(_0535_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _8058_ (.CLK(\clknet_leaf_37_u_dsync.out_clk ),
    .D(_0536_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _8059_ (.CLK(\clknet_leaf_68_u_dsync.out_clk ),
    .D(_0537_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][47] ));
 sky130_fd_sc_hd__dfxtp_1 _8060_ (.CLK(\clknet_leaf_95_u_dsync.out_clk ),
    .D(_0538_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][48] ));
 sky130_fd_sc_hd__dfxtp_1 _8061_ (.CLK(\clknet_leaf_67_u_dsync.out_clk ),
    .D(_0539_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][49] ));
 sky130_fd_sc_hd__dfxtp_1 _8062_ (.CLK(\clknet_leaf_38_u_dsync.out_clk ),
    .D(_0540_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][50] ));
 sky130_fd_sc_hd__dfxtp_1 _8063_ (.CLK(\clknet_leaf_96_u_dsync.out_clk ),
    .D(_0541_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][53] ));
 sky130_fd_sc_hd__dfxtp_1 _8064_ (.CLK(\clknet_leaf_8_u_dsync.out_clk ),
    .D(_0542_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][54] ));
 sky130_fd_sc_hd__dfxtp_1 _8065_ (.CLK(\clknet_leaf_6_u_dsync.out_clk ),
    .D(_0543_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][55] ));
 sky130_fd_sc_hd__dfxtp_1 _8066_ (.CLK(\clknet_leaf_7_u_dsync.out_clk ),
    .D(_0544_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][56] ));
 sky130_fd_sc_hd__dfxtp_1 _8067_ (.CLK(\clknet_leaf_96_u_dsync.out_clk ),
    .D(_0545_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][57] ));
 sky130_fd_sc_hd__dfxtp_1 _8068_ (.CLK(\clknet_leaf_8_u_dsync.out_clk ),
    .D(_0546_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][58] ));
 sky130_fd_sc_hd__dfxtp_1 _8069_ (.CLK(\clknet_leaf_97_u_dsync.out_clk ),
    .D(_0547_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[1][59] ));
 sky130_fd_sc_hd__dfxtp_1 _8070_ (.CLK(\clknet_leaf_100_u_dsync.out_clk ),
    .D(_0548_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8071_ (.CLK(\clknet_leaf_105_u_dsync.out_clk ),
    .D(_0549_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8072_ (.CLK(\clknet_leaf_6_u_dsync.out_clk ),
    .D(_0550_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8073_ (.CLK(\clknet_leaf_97_u_dsync.out_clk ),
    .D(_0551_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8074_ (.CLK(\clknet_leaf_94_u_dsync.out_clk ),
    .D(_0552_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8075_ (.CLK(\clknet_leaf_97_u_dsync.out_clk ),
    .D(_0553_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8076_ (.CLK(\clknet_leaf_97_u_dsync.out_clk ),
    .D(_0554_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8077_ (.CLK(\clknet_leaf_97_u_dsync.out_clk ),
    .D(_0555_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8078_ (.CLK(\clknet_leaf_98_u_dsync.out_clk ),
    .D(_0556_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8079_ (.CLK(\clknet_leaf_101_u_dsync.out_clk ),
    .D(_0557_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8080_ (.CLK(\clknet_leaf_100_u_dsync.out_clk ),
    .D(_0558_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8081_ (.CLK(\clknet_leaf_90_u_dsync.out_clk ),
    .D(_0559_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8082_ (.CLK(\clknet_leaf_88_u_dsync.out_clk ),
    .D(_0560_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8083_ (.CLK(\clknet_leaf_89_u_dsync.out_clk ),
    .D(_0561_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8084_ (.CLK(\clknet_leaf_70_u_dsync.out_clk ),
    .D(_0562_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8085_ (.CLK(\clknet_leaf_70_u_dsync.out_clk ),
    .D(_0563_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8086_ (.CLK(\clknet_leaf_70_u_dsync.out_clk ),
    .D(_0564_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8087_ (.CLK(\clknet_leaf_93_u_dsync.out_clk ),
    .D(_0565_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8088_ (.CLK(\clknet_leaf_86_u_dsync.out_clk ),
    .D(_0566_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8089_ (.CLK(\clknet_leaf_93_u_dsync.out_clk ),
    .D(_0567_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8090_ (.CLK(\clknet_leaf_93_u_dsync.out_clk ),
    .D(_0568_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8091_ (.CLK(\clknet_leaf_86_u_dsync.out_clk ),
    .D(_0569_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8092_ (.CLK(\clknet_leaf_86_u_dsync.out_clk ),
    .D(_0570_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8093_ (.CLK(\clknet_leaf_69_u_dsync.out_clk ),
    .D(_0571_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8094_ (.CLK(\clknet_leaf_93_u_dsync.out_clk ),
    .D(_0572_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8095_ (.CLK(\clknet_leaf_69_u_dsync.out_clk ),
    .D(_0573_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8096_ (.CLK(\clknet_leaf_88_u_dsync.out_clk ),
    .D(_0574_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8097_ (.CLK(\clknet_leaf_87_u_dsync.out_clk ),
    .D(_0575_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8098_ (.CLK(\clknet_leaf_94_u_dsync.out_clk ),
    .D(_0576_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _8099_ (.CLK(\clknet_leaf_92_u_dsync.out_clk ),
    .D(_0577_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _8100_ (.CLK(\clknet_leaf_87_u_dsync.out_clk ),
    .D(_0578_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _8101_ (.CLK(\clknet_leaf_94_u_dsync.out_clk ),
    .D(_0579_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _8102_ (.CLK(\clknet_leaf_89_u_dsync.out_clk ),
    .D(_0580_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _8103_ (.CLK(\clknet_leaf_92_u_dsync.out_clk ),
    .D(_0581_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _8104_ (.CLK(\clknet_leaf_87_u_dsync.out_clk ),
    .D(_0582_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _8105_ (.CLK(\clknet_leaf_92_u_dsync.out_clk ),
    .D(_0583_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _8106_ (.CLK(\clknet_leaf_87_u_dsync.out_clk ),
    .D(_0584_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _8107_ (.CLK(\clknet_leaf_91_u_dsync.out_clk ),
    .D(_0585_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _8108_ (.CLK(\clknet_leaf_92_u_dsync.out_clk ),
    .D(_0586_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _8109_ (.CLK(\clknet_leaf_91_u_dsync.out_clk ),
    .D(_0587_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _8110_ (.CLK(\clknet_leaf_90_u_dsync.out_clk ),
    .D(_0588_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _8111_ (.CLK(\clknet_leaf_101_u_dsync.out_clk ),
    .D(_0589_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _8112_ (.CLK(\clknet_leaf_88_u_dsync.out_clk ),
    .D(_0590_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _8113_ (.CLK(\clknet_leaf_86_u_dsync.out_clk ),
    .D(_0591_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][47] ));
 sky130_fd_sc_hd__dfxtp_1 _8114_ (.CLK(\clknet_leaf_91_u_dsync.out_clk ),
    .D(_0592_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][48] ));
 sky130_fd_sc_hd__dfxtp_1 _8115_ (.CLK(\clknet_leaf_90_u_dsync.out_clk ),
    .D(_0593_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][49] ));
 sky130_fd_sc_hd__dfxtp_1 _8116_ (.CLK(\clknet_leaf_91_u_dsync.out_clk ),
    .D(_0594_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][50] ));
 sky130_fd_sc_hd__dfxtp_1 _8117_ (.CLK(\clknet_leaf_100_u_dsync.out_clk ),
    .D(_0595_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][53] ));
 sky130_fd_sc_hd__dfxtp_1 _8118_ (.CLK(\clknet_leaf_106_u_dsync.out_clk ),
    .D(_0596_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][54] ));
 sky130_fd_sc_hd__dfxtp_1 _8119_ (.CLK(\clknet_leaf_101_u_dsync.out_clk ),
    .D(_0597_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][55] ));
 sky130_fd_sc_hd__dfxtp_1 _8120_ (.CLK(\clknet_leaf_100_u_dsync.out_clk ),
    .D(_0598_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][56] ));
 sky130_fd_sc_hd__dfxtp_1 _8121_ (.CLK(\clknet_leaf_90_u_dsync.out_clk ),
    .D(_0599_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][57] ));
 sky130_fd_sc_hd__dfxtp_1 _8122_ (.CLK(\clknet_leaf_88_u_dsync.out_clk ),
    .D(_0600_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][58] ));
 sky130_fd_sc_hd__dfxtp_1 _8123_ (.CLK(\clknet_leaf_101_u_dsync.out_clk ),
    .D(_0601_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][59] ));
 sky130_fd_sc_hd__dfxtp_1 _8124_ (.CLK(\clknet_leaf_105_u_dsync.out_clk ),
    .D(_0602_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][60] ));
 sky130_fd_sc_hd__dfxtp_1 _8125_ (.CLK(\clknet_leaf_106_u_dsync.out_clk ),
    .D(_0603_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][61] ));
 sky130_fd_sc_hd__dfxtp_1 _8126_ (.CLK(\clknet_leaf_107_u_dsync.out_clk ),
    .D(_0604_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][62] ));
 sky130_fd_sc_hd__dfxtp_1 _8127_ (.CLK(\clknet_leaf_107_u_dsync.out_clk ),
    .D(_0605_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][63] ));
 sky130_fd_sc_hd__dfxtp_1 _8128_ (.CLK(\clknet_leaf_107_u_dsync.out_clk ),
    .D(_0606_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][64] ));
 sky130_fd_sc_hd__dfxtp_1 _8129_ (.CLK(\clknet_leaf_108_u_dsync.out_clk ),
    .D(_0607_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][65] ));
 sky130_fd_sc_hd__dfxtp_1 _8130_ (.CLK(\clknet_leaf_107_u_dsync.out_clk ),
    .D(_0608_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][66] ));
 sky130_fd_sc_hd__dfxtp_1 _8131_ (.CLK(\clknet_leaf_102_u_dsync.out_clk ),
    .D(_0609_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][67] ));
 sky130_fd_sc_hd__dfxtp_1 _8132_ (.CLK(\clknet_leaf_102_u_dsync.out_clk ),
    .D(_0610_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][68] ));
 sky130_fd_sc_hd__dfxtp_1 _8133_ (.CLK(\clknet_leaf_103_u_dsync.out_clk ),
    .D(_0611_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][69] ));
 sky130_fd_sc_hd__dfxtp_1 _8134_ (.CLK(\clknet_leaf_90_u_dsync.out_clk ),
    .D(_0612_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][70] ));
 sky130_fd_sc_hd__dfxtp_1 _8135_ (.CLK(\clknet_leaf_106_u_dsync.out_clk ),
    .D(_0613_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][71] ));
 sky130_fd_sc_hd__dfxtp_1 _8136_ (.CLK(\clknet_leaf_102_u_dsync.out_clk ),
    .D(_0614_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][72] ));
 sky130_fd_sc_hd__dfxtp_1 _8137_ (.CLK(\clknet_leaf_102_u_dsync.out_clk ),
    .D(_0615_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][73] ));
 sky130_fd_sc_hd__dfxtp_1 _8138_ (.CLK(\clknet_leaf_103_u_dsync.out_clk ),
    .D(_0616_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][74] ));
 sky130_fd_sc_hd__dfxtp_1 _8139_ (.CLK(\clknet_leaf_104_u_dsync.out_clk ),
    .D(_0617_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][75] ));
 sky130_fd_sc_hd__dfxtp_1 _8140_ (.CLK(\clknet_leaf_104_u_dsync.out_clk ),
    .D(_0618_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][76] ));
 sky130_fd_sc_hd__dfxtp_1 _8141_ (.CLK(\clknet_leaf_103_u_dsync.out_clk ),
    .D(_0619_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][77] ));
 sky130_fd_sc_hd__dfxtp_1 _8142_ (.CLK(\clknet_leaf_104_u_dsync.out_clk ),
    .D(_0620_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][78] ));
 sky130_fd_sc_hd__dfxtp_1 _8143_ (.CLK(\clknet_leaf_103_u_dsync.out_clk ),
    .D(_0621_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][79] ));
 sky130_fd_sc_hd__dfxtp_1 _8144_ (.CLK(\clknet_leaf_105_u_dsync.out_clk ),
    .D(_0622_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][80] ));
 sky130_fd_sc_hd__dfxtp_1 _8145_ (.CLK(\clknet_leaf_105_u_dsync.out_clk ),
    .D(_0623_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][81] ));
 sky130_fd_sc_hd__dfxtp_1 _8146_ (.CLK(\clknet_leaf_103_u_dsync.out_clk ),
    .D(_0624_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[0][82] ));
 sky130_fd_sc_hd__dfrtp_1 _8147_ (.CLK(\clknet_leaf_48_u_dsync.out_clk ),
    .D(_0625_),
    .RESET_B(net916),
    .Q(\u_s2.u_sync_wbb.u_resp_if.rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_4 _8148_ (.CLK(\clknet_leaf_47_u_dsync.out_clk ),
    .D(_0626_),
    .RESET_B(net915),
    .Q(\u_s2.u_sync_wbb.u_resp_if.rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_2 _8149_ (.CLK(\clknet_leaf_46_u_dsync.out_clk ),
    .D(_0627_),
    .RESET_B(net915),
    .Q(\u_s2.u_sync_wbb.u_resp_if.rd_ptr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8150_ (.CLK(\clknet_leaf_80_u_dsync.out_clk ),
    .D(_0628_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8151_ (.CLK(\clknet_leaf_79_u_dsync.out_clk ),
    .D(_0629_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8152_ (.CLK(\clknet_leaf_75_u_dsync.out_clk ),
    .D(_0630_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8153_ (.CLK(\clknet_leaf_79_u_dsync.out_clk ),
    .D(_0631_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8154_ (.CLK(\clknet_leaf_75_u_dsync.out_clk ),
    .D(_0632_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8155_ (.CLK(\clknet_leaf_75_u_dsync.out_clk ),
    .D(_0633_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8156_ (.CLK(\clknet_leaf_76_u_dsync.out_clk ),
    .D(_0634_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8157_ (.CLK(\clknet_leaf_76_u_dsync.out_clk ),
    .D(_0635_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8158_ (.CLK(\clknet_leaf_79_u_dsync.out_clk ),
    .D(_0636_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8159_ (.CLK(\clknet_leaf_78_u_dsync.out_clk ),
    .D(_0637_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8160_ (.CLK(\clknet_leaf_79_u_dsync.out_clk ),
    .D(_0638_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8161_ (.CLK(\clknet_leaf_80_u_dsync.out_clk ),
    .D(_0639_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8162_ (.CLK(\clknet_leaf_80_u_dsync.out_clk ),
    .D(_0640_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8163_ (.CLK(\clknet_leaf_78_u_dsync.out_clk ),
    .D(_0641_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8164_ (.CLK(\clknet_leaf_81_u_dsync.out_clk ),
    .D(_0642_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8165_ (.CLK(\clknet_leaf_76_u_dsync.out_clk ),
    .D(_0643_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8166_ (.CLK(\clknet_leaf_82_u_dsync.out_clk ),
    .D(_0644_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8167_ (.CLK(\clknet_leaf_76_u_dsync.out_clk ),
    .D(_0645_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8168_ (.CLK(\clknet_leaf_76_u_dsync.out_clk ),
    .D(_0646_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8169_ (.CLK(\clknet_leaf_80_u_dsync.out_clk ),
    .D(_0647_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8170_ (.CLK(\clknet_leaf_81_u_dsync.out_clk ),
    .D(_0648_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8171_ (.CLK(\clknet_leaf_77_u_dsync.out_clk ),
    .D(_0649_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8172_ (.CLK(\clknet_leaf_82_u_dsync.out_clk ),
    .D(_0650_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8173_ (.CLK(\clknet_leaf_85_u_dsync.out_clk ),
    .D(_0651_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8174_ (.CLK(\clknet_leaf_79_u_dsync.out_clk ),
    .D(_0652_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8175_ (.CLK(\clknet_leaf_85_u_dsync.out_clk ),
    .D(_0653_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8176_ (.CLK(\clknet_leaf_80_u_dsync.out_clk ),
    .D(_0654_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8177_ (.CLK(\clknet_leaf_82_u_dsync.out_clk ),
    .D(_0655_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8178_ (.CLK(\clknet_leaf_80_u_dsync.out_clk ),
    .D(_0656_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8179_ (.CLK(\clknet_leaf_81_u_dsync.out_clk ),
    .D(_0657_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8180_ (.CLK(\clknet_leaf_83_u_dsync.out_clk ),
    .D(_0658_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8181_ (.CLK(\clknet_leaf_79_u_dsync.out_clk ),
    .D(_0659_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8182_ (.CLK(\clknet_leaf_80_u_dsync.out_clk ),
    .D(_0660_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8183_ (.CLK(\clknet_leaf_78_u_dsync.out_clk ),
    .D(_0661_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8184_ (.CLK(\clknet_leaf_76_u_dsync.out_clk ),
    .D(_0662_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8185_ (.CLK(\clknet_leaf_79_u_dsync.out_clk ),
    .D(_0663_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8186_ (.CLK(\clknet_leaf_75_u_dsync.out_clk ),
    .D(_0664_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8187_ (.CLK(\clknet_leaf_75_u_dsync.out_clk ),
    .D(_0665_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8188_ (.CLK(\clknet_leaf_76_u_dsync.out_clk ),
    .D(_0666_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8189_ (.CLK(\clknet_leaf_76_u_dsync.out_clk ),
    .D(_0667_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8190_ (.CLK(\clknet_leaf_79_u_dsync.out_clk ),
    .D(_0668_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8191_ (.CLK(\clknet_leaf_78_u_dsync.out_clk ),
    .D(_0669_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8192_ (.CLK(\clknet_leaf_79_u_dsync.out_clk ),
    .D(_0670_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8193_ (.CLK(\clknet_leaf_80_u_dsync.out_clk ),
    .D(_0671_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8194_ (.CLK(\clknet_leaf_81_u_dsync.out_clk ),
    .D(_0672_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8195_ (.CLK(\clknet_leaf_85_u_dsync.out_clk ),
    .D(_0673_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8196_ (.CLK(\clknet_leaf_81_u_dsync.out_clk ),
    .D(_0674_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8197_ (.CLK(\clknet_leaf_79_u_dsync.out_clk ),
    .D(_0675_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8198_ (.CLK(\clknet_leaf_81_u_dsync.out_clk ),
    .D(_0676_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8199_ (.CLK(\clknet_leaf_76_u_dsync.out_clk ),
    .D(_0677_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8200_ (.CLK(\clknet_leaf_76_u_dsync.out_clk ),
    .D(_0678_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8201_ (.CLK(\clknet_leaf_80_u_dsync.out_clk ),
    .D(_0679_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8202_ (.CLK(\clknet_leaf_81_u_dsync.out_clk ),
    .D(_0680_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8203_ (.CLK(\clknet_leaf_71_u_dsync.out_clk ),
    .D(_0681_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8204_ (.CLK(\clknet_leaf_82_u_dsync.out_clk ),
    .D(_0682_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8205_ (.CLK(\clknet_leaf_85_u_dsync.out_clk ),
    .D(_0683_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8206_ (.CLK(\clknet_leaf_79_u_dsync.out_clk ),
    .D(_0684_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8207_ (.CLK(\clknet_leaf_78_u_dsync.out_clk ),
    .D(_0685_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8208_ (.CLK(\clknet_leaf_79_u_dsync.out_clk ),
    .D(_0686_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8209_ (.CLK(\clknet_leaf_82_u_dsync.out_clk ),
    .D(_0687_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8210_ (.CLK(\clknet_leaf_80_u_dsync.out_clk ),
    .D(_0688_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8211_ (.CLK(\clknet_leaf_81_u_dsync.out_clk ),
    .D(_0689_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8212_ (.CLK(\clknet_leaf_82_u_dsync.out_clk ),
    .D(_0690_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8213_ (.CLK(\clknet_leaf_79_u_dsync.out_clk ),
    .D(_0691_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8214_ (.CLK(\clknet_leaf_85_u_dsync.out_clk ),
    .D(_0692_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8215_ (.CLK(\clknet_leaf_78_u_dsync.out_clk ),
    .D(_0693_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8216_ (.CLK(\clknet_leaf_76_u_dsync.out_clk ),
    .D(_0694_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8217_ (.CLK(\clknet_leaf_79_u_dsync.out_clk ),
    .D(_0695_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8218_ (.CLK(\clknet_leaf_76_u_dsync.out_clk ),
    .D(_0696_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8219_ (.CLK(\clknet_leaf_75_u_dsync.out_clk ),
    .D(_0697_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8220_ (.CLK(\clknet_leaf_76_u_dsync.out_clk ),
    .D(_0698_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8221_ (.CLK(\clknet_leaf_76_u_dsync.out_clk ),
    .D(_0699_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8222_ (.CLK(\clknet_leaf_79_u_dsync.out_clk ),
    .D(_0700_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8223_ (.CLK(\clknet_leaf_78_u_dsync.out_clk ),
    .D(_0701_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8224_ (.CLK(\clknet_leaf_79_u_dsync.out_clk ),
    .D(_0702_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8225_ (.CLK(\clknet_leaf_80_u_dsync.out_clk ),
    .D(_0703_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8226_ (.CLK(\clknet_leaf_81_u_dsync.out_clk ),
    .D(_0704_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8227_ (.CLK(\clknet_leaf_85_u_dsync.out_clk ),
    .D(_0705_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8228_ (.CLK(\clknet_leaf_80_u_dsync.out_clk ),
    .D(_0706_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8229_ (.CLK(\clknet_leaf_76_u_dsync.out_clk ),
    .D(_0707_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8230_ (.CLK(\clknet_leaf_82_u_dsync.out_clk ),
    .D(_0708_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8231_ (.CLK(\clknet_leaf_77_u_dsync.out_clk ),
    .D(_0709_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8232_ (.CLK(\clknet_leaf_77_u_dsync.out_clk ),
    .D(_0710_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8233_ (.CLK(\clknet_leaf_80_u_dsync.out_clk ),
    .D(_0711_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8234_ (.CLK(\clknet_leaf_81_u_dsync.out_clk ),
    .D(_0712_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8235_ (.CLK(\clknet_leaf_71_u_dsync.out_clk ),
    .D(_0713_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8236_ (.CLK(\clknet_leaf_82_u_dsync.out_clk ),
    .D(_0714_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8237_ (.CLK(\clknet_leaf_84_u_dsync.out_clk ),
    .D(_0715_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8238_ (.CLK(\clknet_leaf_79_u_dsync.out_clk ),
    .D(_0716_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8239_ (.CLK(\clknet_leaf_78_u_dsync.out_clk ),
    .D(_0717_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8240_ (.CLK(\clknet_leaf_78_u_dsync.out_clk ),
    .D(_0718_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8241_ (.CLK(\clknet_leaf_85_u_dsync.out_clk ),
    .D(_0719_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8242_ (.CLK(\clknet_leaf_82_u_dsync.out_clk ),
    .D(_0720_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8243_ (.CLK(\clknet_leaf_81_u_dsync.out_clk ),
    .D(_0721_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8244_ (.CLK(\clknet_leaf_83_u_dsync.out_clk ),
    .D(_0722_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8245_ (.CLK(\clknet_leaf_78_u_dsync.out_clk ),
    .D(_0723_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8246_ (.CLK(\clknet_leaf_80_u_dsync.out_clk ),
    .D(_0724_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8247_ (.CLK(\clknet_leaf_78_u_dsync.out_clk ),
    .D(_0725_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8248_ (.CLK(\clknet_leaf_76_u_dsync.out_clk ),
    .D(_0726_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8249_ (.CLK(\clknet_leaf_79_u_dsync.out_clk ),
    .D(_0727_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8250_ (.CLK(\clknet_leaf_75_u_dsync.out_clk ),
    .D(_0728_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8251_ (.CLK(\clknet_leaf_75_u_dsync.out_clk ),
    .D(_0729_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8252_ (.CLK(\clknet_leaf_76_u_dsync.out_clk ),
    .D(_0730_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8253_ (.CLK(\clknet_leaf_76_u_dsync.out_clk ),
    .D(_0731_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8254_ (.CLK(\clknet_leaf_79_u_dsync.out_clk ),
    .D(_0732_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8255_ (.CLK(\clknet_leaf_77_u_dsync.out_clk ),
    .D(_0733_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8256_ (.CLK(\clknet_leaf_80_u_dsync.out_clk ),
    .D(_0734_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8257_ (.CLK(\clknet_leaf_80_u_dsync.out_clk ),
    .D(_0735_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8258_ (.CLK(\clknet_leaf_80_u_dsync.out_clk ),
    .D(_0736_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8259_ (.CLK(\clknet_leaf_85_u_dsync.out_clk ),
    .D(_0737_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8260_ (.CLK(\clknet_leaf_80_u_dsync.out_clk ),
    .D(_0738_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8261_ (.CLK(\clknet_leaf_76_u_dsync.out_clk ),
    .D(_0739_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8262_ (.CLK(\clknet_leaf_82_u_dsync.out_clk ),
    .D(_0740_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8263_ (.CLK(\clknet_leaf_76_u_dsync.out_clk ),
    .D(_0741_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8264_ (.CLK(\clknet_leaf_77_u_dsync.out_clk ),
    .D(_0742_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8265_ (.CLK(\clknet_leaf_80_u_dsync.out_clk ),
    .D(_0743_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8266_ (.CLK(\clknet_leaf_80_u_dsync.out_clk ),
    .D(_0744_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8267_ (.CLK(\clknet_leaf_71_u_dsync.out_clk ),
    .D(_0745_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8268_ (.CLK(\clknet_leaf_82_u_dsync.out_clk ),
    .D(_0746_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8269_ (.CLK(\clknet_leaf_84_u_dsync.out_clk ),
    .D(_0747_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8270_ (.CLK(\clknet_leaf_79_u_dsync.out_clk ),
    .D(_0748_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8271_ (.CLK(\clknet_leaf_78_u_dsync.out_clk ),
    .D(_0749_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8272_ (.CLK(\clknet_leaf_78_u_dsync.out_clk ),
    .D(_0750_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8273_ (.CLK(\clknet_leaf_83_u_dsync.out_clk ),
    .D(_0751_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8274_ (.CLK(\clknet_leaf_82_u_dsync.out_clk ),
    .D(_0752_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8275_ (.CLK(\clknet_leaf_81_u_dsync.out_clk ),
    .D(_0753_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8276_ (.CLK(\clknet_leaf_83_u_dsync.out_clk ),
    .D(_0754_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8277_ (.CLK(\clknet_leaf_78_u_dsync.out_clk ),
    .D(_0755_),
    .Q(\u_s0.u_sync_wbb.u_resp_if.mem[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8278_ (.CLK(\clknet_leaf_28_u_dsync.out_clk ),
    .D(_0756_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8279_ (.CLK(\clknet_leaf_30_u_dsync.out_clk ),
    .D(_0757_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8280_ (.CLK(\clknet_leaf_28_u_dsync.out_clk ),
    .D(_0758_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8281_ (.CLK(\clknet_leaf_29_u_dsync.out_clk ),
    .D(_0759_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8282_ (.CLK(\clknet_leaf_35_u_dsync.out_clk ),
    .D(_0760_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8283_ (.CLK(\clknet_leaf_28_u_dsync.out_clk ),
    .D(_0761_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8284_ (.CLK(\clknet_leaf_35_u_dsync.out_clk ),
    .D(_0762_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8285_ (.CLK(\clknet_leaf_33_u_dsync.out_clk ),
    .D(_0763_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8286_ (.CLK(\clknet_leaf_27_u_dsync.out_clk ),
    .D(_0764_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8287_ (.CLK(\clknet_leaf_31_u_dsync.out_clk ),
    .D(_0765_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8288_ (.CLK(\clknet_leaf_30_u_dsync.out_clk ),
    .D(_0766_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8289_ (.CLK(\clknet_leaf_32_u_dsync.out_clk ),
    .D(_0767_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8290_ (.CLK(\clknet_leaf_36_u_dsync.out_clk ),
    .D(_0768_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8291_ (.CLK(\clknet_leaf_43_u_dsync.out_clk ),
    .D(_0769_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8292_ (.CLK(\clknet_leaf_43_u_dsync.out_clk ),
    .D(_0770_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8293_ (.CLK(\clknet_leaf_45_u_dsync.out_clk ),
    .D(_0771_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8294_ (.CLK(\clknet_leaf_43_u_dsync.out_clk ),
    .D(_0772_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8295_ (.CLK(\clknet_leaf_48_u_dsync.out_clk ),
    .D(_0773_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8296_ (.CLK(\clknet_leaf_43_u_dsync.out_clk ),
    .D(_0774_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8297_ (.CLK(\clknet_leaf_43_u_dsync.out_clk ),
    .D(_0775_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8298_ (.CLK(\clknet_leaf_46_u_dsync.out_clk ),
    .D(_0776_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8299_ (.CLK(\clknet_leaf_41_u_dsync.out_clk ),
    .D(_0777_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8300_ (.CLK(\clknet_leaf_44_u_dsync.out_clk ),
    .D(_0778_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8301_ (.CLK(\clknet_leaf_47_u_dsync.out_clk ),
    .D(_0779_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8302_ (.CLK(\clknet_leaf_40_u_dsync.out_clk ),
    .D(_0780_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8303_ (.CLK(\clknet_leaf_44_u_dsync.out_clk ),
    .D(_0781_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8304_ (.CLK(\clknet_leaf_40_u_dsync.out_clk ),
    .D(_0782_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8305_ (.CLK(\clknet_leaf_45_u_dsync.out_clk ),
    .D(_0783_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][32] ));
 sky130_fd_sc_hd__dfxtp_1 _8306_ (.CLK(\clknet_leaf_43_u_dsync.out_clk ),
    .D(_0784_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][33] ));
 sky130_fd_sc_hd__dfxtp_1 _8307_ (.CLK(\clknet_leaf_45_u_dsync.out_clk ),
    .D(_0785_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][34] ));
 sky130_fd_sc_hd__dfxtp_1 _8308_ (.CLK(\clknet_leaf_32_u_dsync.out_clk ),
    .D(_0786_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][35] ));
 sky130_fd_sc_hd__dfxtp_1 _8309_ (.CLK(\clknet_leaf_45_u_dsync.out_clk ),
    .D(_0787_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][36] ));
 sky130_fd_sc_hd__dfxtp_1 _8310_ (.CLK(\clknet_leaf_31_u_dsync.out_clk ),
    .D(_0788_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][37] ));
 sky130_fd_sc_hd__dfxtp_1 _8311_ (.CLK(\clknet_leaf_40_u_dsync.out_clk ),
    .D(_0789_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][38] ));
 sky130_fd_sc_hd__dfxtp_1 _8312_ (.CLK(\clknet_leaf_41_u_dsync.out_clk ),
    .D(_0790_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][39] ));
 sky130_fd_sc_hd__dfxtp_1 _8313_ (.CLK(\clknet_leaf_44_u_dsync.out_clk ),
    .D(_0791_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][40] ));
 sky130_fd_sc_hd__dfxtp_1 _8314_ (.CLK(\clknet_leaf_39_u_dsync.out_clk ),
    .D(_0792_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][41] ));
 sky130_fd_sc_hd__dfxtp_1 _8315_ (.CLK(\clknet_leaf_33_u_dsync.out_clk ),
    .D(_0793_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][42] ));
 sky130_fd_sc_hd__dfxtp_1 _8316_ (.CLK(\clknet_leaf_33_u_dsync.out_clk ),
    .D(_0794_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][43] ));
 sky130_fd_sc_hd__dfxtp_1 _8317_ (.CLK(\clknet_leaf_46_u_dsync.out_clk ),
    .D(_0795_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][44] ));
 sky130_fd_sc_hd__dfxtp_1 _8318_ (.CLK(\clknet_leaf_31_u_dsync.out_clk ),
    .D(_0796_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][45] ));
 sky130_fd_sc_hd__dfxtp_1 _8319_ (.CLK(\clknet_leaf_36_u_dsync.out_clk ),
    .D(_0797_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][46] ));
 sky130_fd_sc_hd__dfxtp_1 _8320_ (.CLK(\clknet_leaf_36_u_dsync.out_clk ),
    .D(_0798_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][47] ));
 sky130_fd_sc_hd__dfxtp_1 _8321_ (.CLK(\clknet_leaf_33_u_dsync.out_clk ),
    .D(_0799_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][48] ));
 sky130_fd_sc_hd__dfxtp_1 _8322_ (.CLK(\clknet_leaf_36_u_dsync.out_clk ),
    .D(_0800_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][49] ));
 sky130_fd_sc_hd__dfxtp_1 _8323_ (.CLK(\clknet_leaf_31_u_dsync.out_clk ),
    .D(_0801_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][50] ));
 sky130_fd_sc_hd__dfxtp_1 _8324_ (.CLK(\clknet_leaf_33_u_dsync.out_clk ),
    .D(_0802_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][53] ));
 sky130_fd_sc_hd__dfxtp_1 _8325_ (.CLK(\clknet_leaf_27_u_dsync.out_clk ),
    .D(_0803_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][54] ));
 sky130_fd_sc_hd__dfxtp_1 _8326_ (.CLK(\clknet_leaf_33_u_dsync.out_clk ),
    .D(_0804_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][55] ));
 sky130_fd_sc_hd__dfxtp_1 _8327_ (.CLK(\clknet_leaf_33_u_dsync.out_clk ),
    .D(_0805_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][56] ));
 sky130_fd_sc_hd__dfxtp_1 _8328_ (.CLK(\clknet_leaf_34_u_dsync.out_clk ),
    .D(_0806_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][57] ));
 sky130_fd_sc_hd__dfxtp_1 _8329_ (.CLK(\clknet_leaf_35_u_dsync.out_clk ),
    .D(_0807_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][58] ));
 sky130_fd_sc_hd__dfxtp_1 _8330_ (.CLK(\clknet_leaf_34_u_dsync.out_clk ),
    .D(_0808_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][59] ));
 sky130_fd_sc_hd__dfxtp_1 _8331_ (.CLK(\clknet_leaf_35_u_dsync.out_clk ),
    .D(_0809_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][60] ));
 sky130_fd_sc_hd__dfxtp_1 _8332_ (.CLK(\clknet_leaf_35_u_dsync.out_clk ),
    .D(_0810_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[3][61] ));
 sky130_fd_sc_hd__dfrtp_1 _8333_ (.CLK(\clknet_leaf_86_u_dsync.out_clk ),
    .D(_0811_),
    .RESET_B(net842),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8334_ (.CLK(\clknet_leaf_83_u_dsync.out_clk ),
    .D(_0812_),
    .RESET_B(net838),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8335_ (.CLK(\clknet_leaf_84_u_dsync.out_clk ),
    .D(_0813_),
    .RESET_B(net838),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8336_ (.CLK(\clknet_leaf_70_u_dsync.out_clk ),
    .D(_0814_),
    .RESET_B(net852),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8337_ (.CLK(\clknet_leaf_87_u_dsync.out_clk ),
    .D(_0815_),
    .RESET_B(net838),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8338_ (.CLK(\clknet_leaf_77_u_dsync.out_clk ),
    .D(_0816_),
    .RESET_B(net852),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[5] ));
 sky130_fd_sc_hd__dfrtp_1 _8339_ (.CLK(\clknet_leaf_70_u_dsync.out_clk ),
    .D(_0817_),
    .RESET_B(net851),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[6] ));
 sky130_fd_sc_hd__dfrtp_1 _8340_ (.CLK(\clknet_leaf_71_u_dsync.out_clk ),
    .D(_0818_),
    .RESET_B(net852),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[7] ));
 sky130_fd_sc_hd__dfrtp_1 _8341_ (.CLK(\clknet_leaf_70_u_dsync.out_clk ),
    .D(_0819_),
    .RESET_B(net852),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[8] ));
 sky130_fd_sc_hd__dfrtp_1 _8342_ (.CLK(\clknet_leaf_78_u_dsync.out_clk ),
    .D(_0820_),
    .RESET_B(net844),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[9] ));
 sky130_fd_sc_hd__dfrtp_1 _8343_ (.CLK(\clknet_leaf_78_u_dsync.out_clk ),
    .D(_0821_),
    .RESET_B(net842),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[14] ));
 sky130_fd_sc_hd__dfrtp_1 _8344_ (.CLK(\clknet_leaf_89_u_dsync.out_clk ),
    .D(_0822_),
    .RESET_B(net837),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[15] ));
 sky130_fd_sc_hd__dfrtp_1 _8345_ (.CLK(\clknet_leaf_83_u_dsync.out_clk ),
    .D(_0823_),
    .RESET_B(net836),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[16] ));
 sky130_fd_sc_hd__dfrtp_1 _8346_ (.CLK(\clknet_leaf_88_u_dsync.out_clk ),
    .D(_0824_),
    .RESET_B(net834),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[17] ));
 sky130_fd_sc_hd__dfrtp_1 _8347_ (.CLK(\clknet_leaf_70_u_dsync.out_clk ),
    .D(_0825_),
    .RESET_B(net851),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[18] ));
 sky130_fd_sc_hd__dfrtp_1 _8348_ (.CLK(\clknet_leaf_77_u_dsync.out_clk ),
    .D(_0826_),
    .RESET_B(net851),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[19] ));
 sky130_fd_sc_hd__dfrtp_1 _8349_ (.CLK(\clknet_leaf_70_u_dsync.out_clk ),
    .D(_0827_),
    .RESET_B(net852),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[20] ));
 sky130_fd_sc_hd__dfrtp_1 _8350_ (.CLK(\clknet_leaf_93_u_dsync.out_clk ),
    .D(_0828_),
    .RESET_B(net851),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[21] ));
 sky130_fd_sc_hd__dfrtp_1 _8351_ (.CLK(\clknet_leaf_86_u_dsync.out_clk ),
    .D(_0829_),
    .RESET_B(net844),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[22] ));
 sky130_fd_sc_hd__dfrtp_1 _8352_ (.CLK(\clknet_leaf_86_u_dsync.out_clk ),
    .D(_0830_),
    .RESET_B(net842),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[23] ));
 sky130_fd_sc_hd__dfrtp_1 _8353_ (.CLK(\clknet_leaf_70_u_dsync.out_clk ),
    .D(_0831_),
    .RESET_B(net853),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[24] ));
 sky130_fd_sc_hd__dfrtp_1 _8354_ (.CLK(\clknet_leaf_84_u_dsync.out_clk ),
    .D(_0832_),
    .RESET_B(net836),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[25] ));
 sky130_fd_sc_hd__dfrtp_1 _8355_ (.CLK(\clknet_leaf_85_u_dsync.out_clk ),
    .D(_0833_),
    .RESET_B(net843),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[26] ));
 sky130_fd_sc_hd__dfrtp_1 _8356_ (.CLK(\clknet_leaf_69_u_dsync.out_clk ),
    .D(_0834_),
    .RESET_B(net852),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[27] ));
 sky130_fd_sc_hd__dfrtp_1 _8357_ (.CLK(\clknet_leaf_85_u_dsync.out_clk ),
    .D(_0835_),
    .RESET_B(net843),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[28] ));
 sky130_fd_sc_hd__dfrtp_1 _8358_ (.CLK(\clknet_leaf_68_u_dsync.out_clk ),
    .D(_0836_),
    .RESET_B(net862),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[29] ));
 sky130_fd_sc_hd__dfrtp_1 _8359_ (.CLK(\clknet_leaf_87_u_dsync.out_clk ),
    .D(_0837_),
    .RESET_B(net838),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[30] ));
 sky130_fd_sc_hd__dfrtp_1 _8360_ (.CLK(\clknet_leaf_84_u_dsync.out_clk ),
    .D(_0838_),
    .RESET_B(net838),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[31] ));
 sky130_fd_sc_hd__dfrtp_1 _8361_ (.CLK(\clknet_leaf_70_u_dsync.out_clk ),
    .D(_0839_),
    .RESET_B(net852),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[32] ));
 sky130_fd_sc_hd__dfrtp_1 _8362_ (.CLK(\clknet_leaf_85_u_dsync.out_clk ),
    .D(_0840_),
    .RESET_B(net842),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[33] ));
 sky130_fd_sc_hd__dfrtp_1 _8363_ (.CLK(\clknet_leaf_87_u_dsync.out_clk ),
    .D(_0841_),
    .RESET_B(net837),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[34] ));
 sky130_fd_sc_hd__dfrtp_1 _8364_ (.CLK(\clknet_leaf_85_u_dsync.out_clk ),
    .D(_0842_),
    .RESET_B(net842),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[35] ));
 sky130_fd_sc_hd__dfrtp_1 _8365_ (.CLK(\clknet_leaf_87_u_dsync.out_clk ),
    .D(_0843_),
    .RESET_B(net839),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[36] ));
 sky130_fd_sc_hd__dfrtp_1 _8366_ (.CLK(\clknet_leaf_86_u_dsync.out_clk ),
    .D(_0844_),
    .RESET_B(net844),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[37] ));
 sky130_fd_sc_hd__dfrtp_1 _8367_ (.CLK(\clknet_leaf_84_u_dsync.out_clk ),
    .D(_0845_),
    .RESET_B(net836),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[38] ));
 sky130_fd_sc_hd__dfrtp_1 _8368_ (.CLK(\clknet_leaf_78_u_dsync.out_clk ),
    .D(_0846_),
    .RESET_B(net844),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[39] ));
 sky130_fd_sc_hd__dfrtp_1 _8369_ (.CLK(\clknet_leaf_87_u_dsync.out_clk ),
    .D(_0847_),
    .RESET_B(net839),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[40] ));
 sky130_fd_sc_hd__dfrtp_1 _8370_ (.CLK(\clknet_leaf_84_u_dsync.out_clk ),
    .D(_0848_),
    .RESET_B(net838),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[41] ));
 sky130_fd_sc_hd__dfrtp_1 _8371_ (.CLK(\clknet_leaf_87_u_dsync.out_clk ),
    .D(_0849_),
    .RESET_B(net839),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[42] ));
 sky130_fd_sc_hd__dfrtp_1 _8372_ (.CLK(\clknet_leaf_86_u_dsync.out_clk ),
    .D(_0850_),
    .RESET_B(net843),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[43] ));
 sky130_fd_sc_hd__dfrtp_1 _8373_ (.CLK(\clknet_leaf_92_u_dsync.out_clk ),
    .D(_0851_),
    .RESET_B(net843),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[44] ));
 sky130_fd_sc_hd__dfrtp_1 _8374_ (.CLK(\clknet_leaf_85_u_dsync.out_clk ),
    .D(_0852_),
    .RESET_B(net842),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[45] ));
 sky130_fd_sc_hd__dfrtp_1 _8375_ (.CLK(\clknet_leaf_88_u_dsync.out_clk ),
    .D(_0853_),
    .RESET_B(net837),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[46] ));
 sky130_fd_sc_hd__dfrtp_1 _8376_ (.CLK(\clknet_leaf_85_u_dsync.out_clk ),
    .D(_0854_),
    .RESET_B(net838),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[47] ));
 sky130_fd_sc_hd__dfrtp_1 _8377_ (.CLK(\clknet_leaf_78_u_dsync.out_clk ),
    .D(_0855_),
    .RESET_B(net844),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[48] ));
 sky130_fd_sc_hd__dfrtp_1 _8378_ (.CLK(\clknet_leaf_84_u_dsync.out_clk ),
    .D(_0856_),
    .RESET_B(net838),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[49] ));
 sky130_fd_sc_hd__dfrtp_1 _8379_ (.CLK(\clknet_leaf_94_u_dsync.out_clk ),
    .D(_0857_),
    .RESET_B(net851),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[50] ));
 sky130_fd_sc_hd__dfrtp_1 _8380_ (.CLK(\clknet_leaf_84_u_dsync.out_clk ),
    .D(_0858_),
    .RESET_B(net838),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[53] ));
 sky130_fd_sc_hd__dfrtp_1 _8381_ (.CLK(\clknet_leaf_85_u_dsync.out_clk ),
    .D(_0859_),
    .RESET_B(net842),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[54] ));
 sky130_fd_sc_hd__dfrtp_1 _8382_ (.CLK(\clknet_leaf_78_u_dsync.out_clk ),
    .D(_0860_),
    .RESET_B(net842),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[55] ));
 sky130_fd_sc_hd__dfrtp_1 _8383_ (.CLK(\clknet_leaf_85_u_dsync.out_clk ),
    .D(_0861_),
    .RESET_B(net843),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[56] ));
 sky130_fd_sc_hd__dfrtp_1 _8384_ (.CLK(\clknet_leaf_89_u_dsync.out_clk ),
    .D(_0862_),
    .RESET_B(net837),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[57] ));
 sky130_fd_sc_hd__dfrtp_1 _8385_ (.CLK(\clknet_leaf_84_u_dsync.out_clk ),
    .D(_0863_),
    .RESET_B(net834),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[58] ));
 sky130_fd_sc_hd__dfrtp_1 _8386_ (.CLK(\clknet_leaf_85_u_dsync.out_clk ),
    .D(_0864_),
    .RESET_B(net843),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[59] ));
 sky130_fd_sc_hd__dfrtp_1 _8387_ (.CLK(\clknet_leaf_83_u_dsync.out_clk ),
    .D(_0865_),
    .RESET_B(net836),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[60] ));
 sky130_fd_sc_hd__dfrtp_1 _8388_ (.CLK(\clknet_leaf_88_u_dsync.out_clk ),
    .D(_0866_),
    .RESET_B(net834),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[61] ));
 sky130_fd_sc_hd__dfrtp_1 _8389_ (.CLK(\clknet_leaf_82_u_dsync.out_clk ),
    .D(_0867_),
    .RESET_B(net834),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[62] ));
 sky130_fd_sc_hd__dfrtp_1 _8390_ (.CLK(\clknet_leaf_83_u_dsync.out_clk ),
    .D(_0868_),
    .RESET_B(net836),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[63] ));
 sky130_fd_sc_hd__dfrtp_1 _8391_ (.CLK(\clknet_leaf_85_u_dsync.out_clk ),
    .D(_0869_),
    .RESET_B(net842),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[64] ));
 sky130_fd_sc_hd__dfrtp_1 _8392_ (.CLK(\clknet_leaf_88_u_dsync.out_clk ),
    .D(_0870_),
    .RESET_B(net837),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[65] ));
 sky130_fd_sc_hd__dfrtp_1 _8393_ (.CLK(\clknet_leaf_83_u_dsync.out_clk ),
    .D(_0871_),
    .RESET_B(net834),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[66] ));
 sky130_fd_sc_hd__dfrtp_1 _8394_ (.CLK(\clknet_leaf_89_u_dsync.out_clk ),
    .D(_0872_),
    .RESET_B(net837),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[67] ));
 sky130_fd_sc_hd__dfrtp_1 _8395_ (.CLK(\clknet_leaf_89_u_dsync.out_clk ),
    .D(_0873_),
    .RESET_B(net837),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[68] ));
 sky130_fd_sc_hd__dfrtp_1 _8396_ (.CLK(\clknet_leaf_88_u_dsync.out_clk ),
    .D(_0874_),
    .RESET_B(net837),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[69] ));
 sky130_fd_sc_hd__dfrtp_1 _8397_ (.CLK(\clknet_leaf_83_u_dsync.out_clk ),
    .D(_0875_),
    .RESET_B(net834),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[70] ));
 sky130_fd_sc_hd__dfrtp_1 _8398_ (.CLK(\clknet_leaf_88_u_dsync.out_clk ),
    .D(_0876_),
    .RESET_B(net836),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[71] ));
 sky130_fd_sc_hd__dfrtp_1 _8399_ (.CLK(\clknet_leaf_88_u_dsync.out_clk ),
    .D(_0877_),
    .RESET_B(net837),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[72] ));
 sky130_fd_sc_hd__dfrtp_1 _8400_ (.CLK(\clknet_leaf_84_u_dsync.out_clk ),
    .D(_0878_),
    .RESET_B(net839),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[73] ));
 sky130_fd_sc_hd__dfrtp_1 _8401_ (.CLK(\clknet_leaf_83_u_dsync.out_clk ),
    .D(_0879_),
    .RESET_B(net834),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[74] ));
 sky130_fd_sc_hd__dfrtp_1 _8402_ (.CLK(\clknet_leaf_84_u_dsync.out_clk ),
    .D(_0880_),
    .RESET_B(net836),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[75] ));
 sky130_fd_sc_hd__dfrtp_1 _8403_ (.CLK(\clknet_leaf_83_u_dsync.out_clk ),
    .D(_0881_),
    .RESET_B(net835),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[76] ));
 sky130_fd_sc_hd__dfrtp_1 _8404_ (.CLK(\clknet_leaf_83_u_dsync.out_clk ),
    .D(_0882_),
    .RESET_B(net835),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[77] ));
 sky130_fd_sc_hd__dfrtp_1 _8405_ (.CLK(\clknet_leaf_83_u_dsync.out_clk ),
    .D(_0883_),
    .RESET_B(net834),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[78] ));
 sky130_fd_sc_hd__dfrtp_1 _8406_ (.CLK(\clknet_leaf_84_u_dsync.out_clk ),
    .D(_0884_),
    .RESET_B(net834),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[79] ));
 sky130_fd_sc_hd__dfrtp_1 _8407_ (.CLK(\clknet_leaf_83_u_dsync.out_clk ),
    .D(_0885_),
    .RESET_B(net835),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[80] ));
 sky130_fd_sc_hd__dfrtp_1 _8408_ (.CLK(\clknet_leaf_84_u_dsync.out_clk ),
    .D(_0886_),
    .RESET_B(net834),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[81] ));
 sky130_fd_sc_hd__dfrtp_1 _8409_ (.CLK(\clknet_leaf_83_u_dsync.out_clk ),
    .D(_0887_),
    .RESET_B(net835),
    .Q(\u_s0.u_sync_wbb.s_cmd_rd_data_l[82] ));
 sky130_fd_sc_hd__dfstp_2 _8410_ (.CLK(\clknet_leaf_11_u_dsync.out_clk ),
    .D(_0003_),
    .SET_B(net885),
    .Q(\u_s1.u_sync_wbb.m_state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _8411_ (.CLK(\clknet_leaf_10_u_dsync.out_clk ),
    .D(net1926),
    .RESET_B(net872),
    .Q(\u_s1.u_sync_wbb.m_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8412_ (.CLK(\clknet_leaf_10_u_dsync.out_clk ),
    .D(_0005_),
    .RESET_B(net878),
    .Q(\u_s1.u_sync_wbb.m_state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8413_ (.CLK(\clknet_leaf_58_u_dsync.out_clk ),
    .D(_0888_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8414_ (.CLK(\clknet_leaf_62_u_dsync.out_clk ),
    .D(_0889_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8415_ (.CLK(\clknet_leaf_57_u_dsync.out_clk ),
    .D(_0890_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8416_ (.CLK(\clknet_leaf_73_u_dsync.out_clk ),
    .D(_0891_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8417_ (.CLK(\clknet_leaf_60_u_dsync.out_clk ),
    .D(_0892_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8418_ (.CLK(\clknet_leaf_56_u_dsync.out_clk ),
    .D(_0893_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8419_ (.CLK(\clknet_leaf_56_u_dsync.out_clk ),
    .D(_0894_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8420_ (.CLK(\clknet_leaf_60_u_dsync.out_clk ),
    .D(_0895_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8421_ (.CLK(\clknet_leaf_58_u_dsync.out_clk ),
    .D(_0896_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8422_ (.CLK(\clknet_leaf_59_u_dsync.out_clk ),
    .D(_0897_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8423_ (.CLK(\clknet_leaf_75_u_dsync.out_clk ),
    .D(_0898_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8424_ (.CLK(\clknet_leaf_74_u_dsync.out_clk ),
    .D(_0899_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8425_ (.CLK(\clknet_leaf_59_u_dsync.out_clk ),
    .D(_0900_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8426_ (.CLK(\clknet_leaf_72_u_dsync.out_clk ),
    .D(_0901_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8427_ (.CLK(\clknet_leaf_59_u_dsync.out_clk ),
    .D(_0902_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8428_ (.CLK(\clknet_leaf_59_u_dsync.out_clk ),
    .D(_0903_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8429_ (.CLK(\clknet_leaf_59_u_dsync.out_clk ),
    .D(_0904_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8430_ (.CLK(\clknet_leaf_71_u_dsync.out_clk ),
    .D(_0905_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8431_ (.CLK(\clknet_leaf_58_u_dsync.out_clk ),
    .D(_0906_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8432_ (.CLK(\clknet_leaf_77_u_dsync.out_clk ),
    .D(_0907_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8433_ (.CLK(\clknet_leaf_73_u_dsync.out_clk ),
    .D(_0908_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8434_ (.CLK(\clknet_leaf_59_u_dsync.out_clk ),
    .D(_0909_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8435_ (.CLK(\clknet_leaf_73_u_dsync.out_clk ),
    .D(_0910_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8436_ (.CLK(\clknet_leaf_74_u_dsync.out_clk ),
    .D(_0911_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8437_ (.CLK(\clknet_leaf_74_u_dsync.out_clk ),
    .D(_0912_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8438_ (.CLK(\clknet_leaf_73_u_dsync.out_clk ),
    .D(_0913_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8439_ (.CLK(\clknet_leaf_75_u_dsync.out_clk ),
    .D(_0914_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8440_ (.CLK(\clknet_leaf_71_u_dsync.out_clk ),
    .D(_0915_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8441_ (.CLK(\clknet_leaf_71_u_dsync.out_clk ),
    .D(_0916_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8442_ (.CLK(\clknet_leaf_73_u_dsync.out_clk ),
    .D(_0917_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8443_ (.CLK(\clknet_leaf_71_u_dsync.out_clk ),
    .D(_0918_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8444_ (.CLK(\clknet_leaf_72_u_dsync.out_clk ),
    .D(_0919_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8445_ (.CLK(\clknet_leaf_59_u_dsync.out_clk ),
    .D(_0920_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8446_ (.CLK(\clknet_leaf_61_u_dsync.out_clk ),
    .D(_0921_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8447_ (.CLK(\clknet_leaf_56_u_dsync.out_clk ),
    .D(_0922_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8448_ (.CLK(\clknet_leaf_74_u_dsync.out_clk ),
    .D(_0923_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8449_ (.CLK(\clknet_leaf_60_u_dsync.out_clk ),
    .D(_0924_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8450_ (.CLK(\clknet_leaf_62_u_dsync.out_clk ),
    .D(_0925_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8451_ (.CLK(\clknet_leaf_56_u_dsync.out_clk ),
    .D(_0926_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8452_ (.CLK(\clknet_leaf_60_u_dsync.out_clk ),
    .D(_0927_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8453_ (.CLK(\clknet_leaf_57_u_dsync.out_clk ),
    .D(_0928_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8454_ (.CLK(\clknet_leaf_59_u_dsync.out_clk ),
    .D(_0929_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8455_ (.CLK(\clknet_leaf_74_u_dsync.out_clk ),
    .D(_0930_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8456_ (.CLK(\clknet_leaf_73_u_dsync.out_clk ),
    .D(_0931_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8457_ (.CLK(\clknet_leaf_60_u_dsync.out_clk ),
    .D(_0932_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8458_ (.CLK(\clknet_leaf_72_u_dsync.out_clk ),
    .D(_0933_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8459_ (.CLK(\clknet_leaf_59_u_dsync.out_clk ),
    .D(_0934_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8460_ (.CLK(\clknet_leaf_60_u_dsync.out_clk ),
    .D(_0935_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8461_ (.CLK(\clknet_leaf_60_u_dsync.out_clk ),
    .D(_0936_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8462_ (.CLK(\clknet_leaf_72_u_dsync.out_clk ),
    .D(_0937_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8463_ (.CLK(\clknet_leaf_60_u_dsync.out_clk ),
    .D(_0938_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8464_ (.CLK(\clknet_leaf_71_u_dsync.out_clk ),
    .D(_0939_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8465_ (.CLK(\clknet_leaf_72_u_dsync.out_clk ),
    .D(_0940_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8466_ (.CLK(\clknet_leaf_74_u_dsync.out_clk ),
    .D(_0941_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8467_ (.CLK(\clknet_leaf_75_u_dsync.out_clk ),
    .D(_0942_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8468_ (.CLK(\clknet_leaf_73_u_dsync.out_clk ),
    .D(_0943_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8469_ (.CLK(\clknet_leaf_75_u_dsync.out_clk ),
    .D(_0944_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8470_ (.CLK(\clknet_leaf_73_u_dsync.out_clk ),
    .D(_0945_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8471_ (.CLK(\clknet_leaf_75_u_dsync.out_clk ),
    .D(_0946_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8472_ (.CLK(\clknet_leaf_71_u_dsync.out_clk ),
    .D(_0947_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8473_ (.CLK(\clknet_leaf_71_u_dsync.out_clk ),
    .D(_0948_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8474_ (.CLK(\clknet_leaf_73_u_dsync.out_clk ),
    .D(_0949_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8475_ (.CLK(\clknet_leaf_71_u_dsync.out_clk ),
    .D(_0950_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8476_ (.CLK(\clknet_leaf_72_u_dsync.out_clk ),
    .D(_0951_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8477_ (.CLK(\clknet_leaf_58_u_dsync.out_clk ),
    .D(_0952_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8478_ (.CLK(\clknet_leaf_61_u_dsync.out_clk ),
    .D(_0953_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8479_ (.CLK(\clknet_leaf_60_u_dsync.out_clk ),
    .D(_0954_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8480_ (.CLK(\clknet_leaf_74_u_dsync.out_clk ),
    .D(_0955_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8481_ (.CLK(\clknet_leaf_60_u_dsync.out_clk ),
    .D(_0956_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8482_ (.CLK(\clknet_leaf_58_u_dsync.out_clk ),
    .D(_0957_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8483_ (.CLK(\clknet_leaf_56_u_dsync.out_clk ),
    .D(_0958_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8484_ (.CLK(\clknet_leaf_60_u_dsync.out_clk ),
    .D(_0959_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8485_ (.CLK(\clknet_leaf_58_u_dsync.out_clk ),
    .D(_0960_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8486_ (.CLK(\clknet_leaf_59_u_dsync.out_clk ),
    .D(_0961_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8487_ (.CLK(\clknet_leaf_75_u_dsync.out_clk ),
    .D(_0962_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8488_ (.CLK(\clknet_leaf_74_u_dsync.out_clk ),
    .D(_0963_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8489_ (.CLK(\clknet_leaf_60_u_dsync.out_clk ),
    .D(_0964_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8490_ (.CLK(\clknet_leaf_72_u_dsync.out_clk ),
    .D(_0965_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8491_ (.CLK(\clknet_leaf_59_u_dsync.out_clk ),
    .D(_0966_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8492_ (.CLK(\clknet_leaf_59_u_dsync.out_clk ),
    .D(_0967_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8493_ (.CLK(\clknet_leaf_59_u_dsync.out_clk ),
    .D(_0968_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8494_ (.CLK(\clknet_leaf_71_u_dsync.out_clk ),
    .D(_0969_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8495_ (.CLK(\clknet_leaf_58_u_dsync.out_clk ),
    .D(_0970_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8496_ (.CLK(\clknet_leaf_75_u_dsync.out_clk ),
    .D(_0971_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8497_ (.CLK(\clknet_leaf_73_u_dsync.out_clk ),
    .D(_0972_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8498_ (.CLK(\clknet_leaf_74_u_dsync.out_clk ),
    .D(_0973_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8499_ (.CLK(\clknet_leaf_74_u_dsync.out_clk ),
    .D(_0974_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8500_ (.CLK(\clknet_leaf_74_u_dsync.out_clk ),
    .D(_0975_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8501_ (.CLK(\clknet_leaf_74_u_dsync.out_clk ),
    .D(_0976_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8502_ (.CLK(\clknet_leaf_73_u_dsync.out_clk ),
    .D(_0977_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8503_ (.CLK(\clknet_leaf_75_u_dsync.out_clk ),
    .D(_0978_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8504_ (.CLK(\clknet_leaf_72_u_dsync.out_clk ),
    .D(_0979_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8505_ (.CLK(\clknet_leaf_72_u_dsync.out_clk ),
    .D(_0980_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8506_ (.CLK(\clknet_leaf_73_u_dsync.out_clk ),
    .D(_0981_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8507_ (.CLK(\clknet_leaf_71_u_dsync.out_clk ),
    .D(_0982_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8508_ (.CLK(\clknet_leaf_72_u_dsync.out_clk ),
    .D(_0983_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8509_ (.CLK(\clknet_leaf_58_u_dsync.out_clk ),
    .D(_0984_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8510_ (.CLK(\clknet_leaf_60_u_dsync.out_clk ),
    .D(_0985_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8511_ (.CLK(\clknet_leaf_57_u_dsync.out_clk ),
    .D(_0986_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8512_ (.CLK(\clknet_leaf_74_u_dsync.out_clk ),
    .D(_0987_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8513_ (.CLK(\clknet_leaf_59_u_dsync.out_clk ),
    .D(_0988_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8514_ (.CLK(\clknet_leaf_58_u_dsync.out_clk ),
    .D(_0989_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8515_ (.CLK(\clknet_leaf_57_u_dsync.out_clk ),
    .D(_0990_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8516_ (.CLK(\clknet_leaf_60_u_dsync.out_clk ),
    .D(_0991_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8517_ (.CLK(\clknet_leaf_58_u_dsync.out_clk ),
    .D(_0992_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8518_ (.CLK(\clknet_leaf_59_u_dsync.out_clk ),
    .D(_0993_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8519_ (.CLK(\clknet_leaf_75_u_dsync.out_clk ),
    .D(_0994_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8520_ (.CLK(\clknet_leaf_74_u_dsync.out_clk ),
    .D(_0995_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8521_ (.CLK(\clknet_leaf_59_u_dsync.out_clk ),
    .D(_0996_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8522_ (.CLK(\clknet_leaf_72_u_dsync.out_clk ),
    .D(_0997_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8523_ (.CLK(\clknet_leaf_59_u_dsync.out_clk ),
    .D(_0998_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8524_ (.CLK(\clknet_leaf_60_u_dsync.out_clk ),
    .D(_0999_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8525_ (.CLK(\clknet_leaf_59_u_dsync.out_clk ),
    .D(_1000_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8526_ (.CLK(\clknet_leaf_72_u_dsync.out_clk ),
    .D(_1001_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8527_ (.CLK(\clknet_leaf_58_u_dsync.out_clk ),
    .D(_1002_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8528_ (.CLK(\clknet_leaf_74_u_dsync.out_clk ),
    .D(_1003_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8529_ (.CLK(\clknet_leaf_73_u_dsync.out_clk ),
    .D(_1004_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8530_ (.CLK(\clknet_leaf_74_u_dsync.out_clk ),
    .D(_1005_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8531_ (.CLK(\clknet_leaf_74_u_dsync.out_clk ),
    .D(_1006_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8532_ (.CLK(\clknet_leaf_74_u_dsync.out_clk ),
    .D(_1007_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8533_ (.CLK(\clknet_leaf_75_u_dsync.out_clk ),
    .D(_1008_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8534_ (.CLK(\clknet_leaf_73_u_dsync.out_clk ),
    .D(_1009_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8535_ (.CLK(\clknet_leaf_75_u_dsync.out_clk ),
    .D(_1010_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8536_ (.CLK(\clknet_leaf_73_u_dsync.out_clk ),
    .D(_1011_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8537_ (.CLK(\clknet_leaf_72_u_dsync.out_clk ),
    .D(_1012_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8538_ (.CLK(\clknet_leaf_74_u_dsync.out_clk ),
    .D(_1013_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8539_ (.CLK(\clknet_leaf_72_u_dsync.out_clk ),
    .D(_1014_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8540_ (.CLK(\clknet_leaf_73_u_dsync.out_clk ),
    .D(_1015_),
    .Q(\u_s1.u_sync_wbb.u_resp_if.mem[0][31] ));
 sky130_fd_sc_hd__dfrtp_4 _8541_ (.CLK(\clknet_leaf_107_u_dsync.out_clk ),
    .D(_1016_),
    .RESET_B(net845),
    .Q(\u_s0.gnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8542_ (.CLK(\clknet_leaf_109_u_dsync.out_clk ),
    .D(_1017_),
    .RESET_B(net845),
    .Q(\u_s0.gnt[1] ));
 sky130_fd_sc_hd__dfrtp_4 _8543_ (.CLK(\clknet_leaf_14_u_dsync.out_clk ),
    .D(_1018_),
    .RESET_B(net870),
    .Q(\u_s1.u_sync_wbb.wbm_ack_o ));
 sky130_fd_sc_hd__dfrtp_4 _8544_ (.CLK(\clknet_leaf_14_u_dsync.out_clk ),
    .D(_1019_),
    .RESET_B(net868),
    .Q(\u_s1.u_sync_wbb.wbm_lack_o ));
 sky130_fd_sc_hd__dfrtp_2 _8545_ (.CLK(\clknet_leaf_11_u_dsync.out_clk ),
    .D(_1020_),
    .RESET_B(net878),
    .Q(\u_s1.u_sync_wbb.m_cmd_wr_en ));
 sky130_fd_sc_hd__dfrtp_4 _8546_ (.CLK(\clknet_leaf_10_u_dsync.out_clk ),
    .D(_1021_),
    .RESET_B(net878),
    .Q(\u_s1.u_sync_wbb.m_resp_rd_en ));
 sky130_fd_sc_hd__dfrtp_2 _8547_ (.CLK(\clknet_leaf_27_u_dsync.out_clk ),
    .D(net1800),
    .RESET_B(net918),
    .Q(\u_s2.u_sync_wbb.m_bl_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8548_ (.CLK(\clknet_leaf_26_u_dsync.out_clk ),
    .D(_1023_),
    .RESET_B(net898),
    .Q(\u_s2.u_sync_wbb.m_bl_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8549_ (.CLK(\clknet_leaf_27_u_dsync.out_clk ),
    .D(_1024_),
    .RESET_B(net894),
    .Q(\u_s2.u_sync_wbb.m_bl_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8550_ (.CLK(\clknet_leaf_34_u_dsync.out_clk ),
    .D(_1025_),
    .RESET_B(net897),
    .Q(\u_s2.u_sync_wbb.m_bl_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_2 _8551_ (.CLK(\clknet_leaf_34_u_dsync.out_clk ),
    .D(_1026_),
    .RESET_B(net897),
    .Q(\u_s2.u_sync_wbb.m_bl_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_2 _8552_ (.CLK(\clknet_leaf_28_u_dsync.out_clk ),
    .D(_1027_),
    .RESET_B(net909),
    .Q(\u_s2.u_sync_wbb.m_bl_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_2 _8553_ (.CLK(\clknet_leaf_28_u_dsync.out_clk ),
    .D(_1028_),
    .RESET_B(net917),
    .Q(\u_s2.u_sync_wbb.m_bl_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _8554_ (.CLK(\clknet_leaf_27_u_dsync.out_clk ),
    .D(_1029_),
    .RESET_B(net898),
    .Q(\u_s2.u_sync_wbb.m_bl_cnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _8555_ (.CLK(\clknet_leaf_28_u_dsync.out_clk ),
    .D(_1030_),
    .RESET_B(net909),
    .Q(\u_s2.u_sync_wbb.m_bl_cnt[8] ));
 sky130_fd_sc_hd__dfrtp_1 _8556_ (.CLK(\clknet_leaf_28_u_dsync.out_clk ),
    .D(_1031_),
    .RESET_B(net913),
    .Q(\u_s2.u_sync_wbb.m_bl_cnt[9] ));
 sky130_fd_sc_hd__dfrtp_1 _8557_ (.CLK(\clknet_leaf_8_u_dsync.out_clk ),
    .D(net1505),
    .RESET_B(net861),
    .Q(\u_s1.u_sync_wbb.wbs_ack_f ));
 sky130_fd_sc_hd__dfrtp_1 _8558_ (.CLK(\clknet_leaf_9_u_dsync.out_clk ),
    .D(net389),
    .RESET_B(net872),
    .Q(\u_s1.u_sync_wbb.wbs_stb_l ));
 sky130_fd_sc_hd__dfrtp_2 _8559_ (.CLK(\clknet_leaf_61_u_dsync.out_clk ),
    .D(_1032_),
    .RESET_B(net863),
    .Q(\u_s1.u_sync_wbb.u_resp_if.wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_4 _8560_ (.CLK(\clknet_leaf_72_u_dsync.out_clk ),
    .D(_1033_),
    .RESET_B(net864),
    .Q(\u_s1.u_sync_wbb.u_resp_if.wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8561_ (.CLK(\clknet_leaf_61_u_dsync.out_clk ),
    .D(_1034_),
    .RESET_B(net879),
    .Q(\u_s1.u_sync_wbb.u_resp_if.wr_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_2 _8562_ (.CLK(\clknet_leaf_11_u_dsync.out_clk ),
    .D(_1035_),
    .RESET_B(net878),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_4 _8563_ (.CLK(\clknet_leaf_9_u_dsync.out_clk ),
    .D(_1036_),
    .RESET_B(net878),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_2 _8564_ (.CLK(\clknet_leaf_36_u_dsync.out_clk ),
    .D(_1037_),
    .RESET_B(net893),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8565_ (.CLK(\clknet_leaf_28_u_dsync.out_clk ),
    .D(_1038_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8566_ (.CLK(\clknet_leaf_32_u_dsync.out_clk ),
    .D(_1039_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8567_ (.CLK(\clknet_leaf_29_u_dsync.out_clk ),
    .D(_1040_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8568_ (.CLK(\clknet_leaf_29_u_dsync.out_clk ),
    .D(_1041_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8569_ (.CLK(\clknet_leaf_35_u_dsync.out_clk ),
    .D(_1042_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8570_ (.CLK(\clknet_leaf_28_u_dsync.out_clk ),
    .D(_1043_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8571_ (.CLK(\clknet_leaf_35_u_dsync.out_clk ),
    .D(_1044_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8572_ (.CLK(\clknet_leaf_34_u_dsync.out_clk ),
    .D(_1045_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8573_ (.CLK(\clknet_leaf_34_u_dsync.out_clk ),
    .D(_1046_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8574_ (.CLK(\clknet_leaf_45_u_dsync.out_clk ),
    .D(_1047_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8575_ (.CLK(\clknet_leaf_31_u_dsync.out_clk ),
    .D(_1048_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8576_ (.CLK(\clknet_leaf_31_u_dsync.out_clk ),
    .D(_1049_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8577_ (.CLK(\clknet_leaf_36_u_dsync.out_clk ),
    .D(_1050_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8578_ (.CLK(\clknet_leaf_42_u_dsync.out_clk ),
    .D(_1051_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8579_ (.CLK(\clknet_leaf_42_u_dsync.out_clk ),
    .D(_1052_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8580_ (.CLK(\clknet_leaf_46_u_dsync.out_clk ),
    .D(_1053_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8581_ (.CLK(\clknet_leaf_49_u_dsync.out_clk ),
    .D(_1054_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8582_ (.CLK(\clknet_leaf_47_u_dsync.out_clk ),
    .D(_1055_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8583_ (.CLK(\clknet_leaf_40_u_dsync.out_clk ),
    .D(_1056_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8584_ (.CLK(\clknet_leaf_41_u_dsync.out_clk ),
    .D(_1057_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8585_ (.CLK(\clknet_leaf_46_u_dsync.out_clk ),
    .D(_1058_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8586_ (.CLK(\clknet_leaf_41_u_dsync.out_clk ),
    .D(_1059_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8587_ (.CLK(\clknet_leaf_43_u_dsync.out_clk ),
    .D(_1060_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8588_ (.CLK(\clknet_leaf_47_u_dsync.out_clk ),
    .D(_1061_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8589_ (.CLK(\clknet_leaf_40_u_dsync.out_clk ),
    .D(_1062_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8590_ (.CLK(\clknet_leaf_44_u_dsync.out_clk ),
    .D(_1063_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8591_ (.CLK(\clknet_leaf_40_u_dsync.out_clk ),
    .D(_1064_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8592_ (.CLK(\clknet_leaf_47_u_dsync.out_clk ),
    .D(_1065_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _8593_ (.CLK(\clknet_leaf_43_u_dsync.out_clk ),
    .D(_1066_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _8594_ (.CLK(\clknet_leaf_45_u_dsync.out_clk ),
    .D(_1067_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _8595_ (.CLK(\clknet_leaf_44_u_dsync.out_clk ),
    .D(_1068_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _8596_ (.CLK(\clknet_leaf_46_u_dsync.out_clk ),
    .D(_1069_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _8597_ (.CLK(\clknet_leaf_31_u_dsync.out_clk ),
    .D(_1070_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _8598_ (.CLK(\clknet_leaf_40_u_dsync.out_clk ),
    .D(_1071_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _8599_ (.CLK(\clknet_leaf_41_u_dsync.out_clk ),
    .D(_1072_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _8600_ (.CLK(\clknet_leaf_40_u_dsync.out_clk ),
    .D(_1073_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _8601_ (.CLK(\clknet_leaf_39_u_dsync.out_clk ),
    .D(_1074_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _8602_ (.CLK(\clknet_leaf_40_u_dsync.out_clk ),
    .D(_1075_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _8603_ (.CLK(\clknet_leaf_44_u_dsync.out_clk ),
    .D(_1076_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _8604_ (.CLK(\clknet_leaf_46_u_dsync.out_clk ),
    .D(_1077_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _8605_ (.CLK(\clknet_leaf_32_u_dsync.out_clk ),
    .D(_1078_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _8606_ (.CLK(\clknet_leaf_36_u_dsync.out_clk ),
    .D(_1079_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _8607_ (.CLK(\clknet_leaf_37_u_dsync.out_clk ),
    .D(_1080_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][47] ));
 sky130_fd_sc_hd__dfxtp_1 _8608_ (.CLK(\clknet_leaf_32_u_dsync.out_clk ),
    .D(_1081_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][48] ));
 sky130_fd_sc_hd__dfxtp_1 _8609_ (.CLK(\clknet_leaf_36_u_dsync.out_clk ),
    .D(_1082_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][49] ));
 sky130_fd_sc_hd__dfxtp_1 _8610_ (.CLK(\clknet_leaf_32_u_dsync.out_clk ),
    .D(_1083_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][50] ));
 sky130_fd_sc_hd__dfxtp_1 _8611_ (.CLK(\clknet_leaf_36_u_dsync.out_clk ),
    .D(_1084_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][53] ));
 sky130_fd_sc_hd__dfxtp_1 _8612_ (.CLK(\clknet_leaf_34_u_dsync.out_clk ),
    .D(_1085_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][54] ));
 sky130_fd_sc_hd__dfxtp_1 _8613_ (.CLK(\clknet_leaf_33_u_dsync.out_clk ),
    .D(_1086_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][55] ));
 sky130_fd_sc_hd__dfxtp_1 _8614_ (.CLK(\clknet_leaf_33_u_dsync.out_clk ),
    .D(_1087_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][56] ));
 sky130_fd_sc_hd__dfxtp_1 _8615_ (.CLK(\clknet_leaf_34_u_dsync.out_clk ),
    .D(_1088_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][57] ));
 sky130_fd_sc_hd__dfxtp_1 _8616_ (.CLK(\clknet_leaf_35_u_dsync.out_clk ),
    .D(_1089_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][58] ));
 sky130_fd_sc_hd__dfxtp_1 _8617_ (.CLK(\clknet_leaf_33_u_dsync.out_clk ),
    .D(_1090_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][59] ));
 sky130_fd_sc_hd__dfxtp_1 _8618_ (.CLK(\clknet_leaf_36_u_dsync.out_clk ),
    .D(_1091_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][60] ));
 sky130_fd_sc_hd__dfxtp_1 _8619_ (.CLK(\clknet_leaf_11_u_dsync.out_clk ),
    .D(_1092_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[0][61] ));
 sky130_fd_sc_hd__dfrtp_1 _8620_ (.CLK(\clknet_leaf_9_u_dsync.out_clk ),
    .D(_1093_),
    .RESET_B(net872),
    .Q(\u_s1.u_sync_wbb.wbs_burst ));
 sky130_fd_sc_hd__dfrtp_1 _8621_ (.CLK(\clknet_leaf_67_u_dsync.out_clk ),
    .D(_1094_),
    .RESET_B(net863),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8622_ (.CLK(\clknet_leaf_9_u_dsync.out_clk ),
    .D(_1095_),
    .RESET_B(net872),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8623_ (.CLK(\clknet_leaf_37_u_dsync.out_clk ),
    .D(_1096_),
    .RESET_B(net885),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.rd_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8624_ (.CLK(\clknet_leaf_64_u_dsync.out_clk ),
    .D(_1097_),
    .RESET_B(net880),
    .Q(\u_s1.u_sync_wbb.u_resp_if.rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_4 _8625_ (.CLK(\clknet_leaf_64_u_dsync.out_clk ),
    .D(_1098_),
    .RESET_B(net880),
    .Q(\u_s1.u_sync_wbb.u_resp_if.rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_2 _8626_ (.CLK(\clknet_leaf_61_u_dsync.out_clk ),
    .D(_1099_),
    .RESET_B(net880),
    .Q(\u_s1.u_sync_wbb.u_resp_if.rd_ptr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8627_ (.CLK(\clknet_leaf_100_u_dsync.out_clk ),
    .D(_1100_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8628_ (.CLK(\clknet_leaf_105_u_dsync.out_clk ),
    .D(_1101_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8629_ (.CLK(\clknet_leaf_6_u_dsync.out_clk ),
    .D(_1102_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8630_ (.CLK(\clknet_leaf_97_u_dsync.out_clk ),
    .D(_1103_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8631_ (.CLK(\clknet_leaf_94_u_dsync.out_clk ),
    .D(_1104_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8632_ (.CLK(\clknet_leaf_98_u_dsync.out_clk ),
    .D(_1105_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8633_ (.CLK(\clknet_leaf_98_u_dsync.out_clk ),
    .D(_1106_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8634_ (.CLK(\clknet_leaf_97_u_dsync.out_clk ),
    .D(_1107_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8635_ (.CLK(\clknet_leaf_97_u_dsync.out_clk ),
    .D(_1108_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8636_ (.CLK(\clknet_leaf_98_u_dsync.out_clk ),
    .D(_1109_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8637_ (.CLK(\clknet_leaf_106_u_dsync.out_clk ),
    .D(_1110_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8638_ (.CLK(\clknet_leaf_102_u_dsync.out_clk ),
    .D(_1111_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8639_ (.CLK(\clknet_leaf_88_u_dsync.out_clk ),
    .D(_1112_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8640_ (.CLK(\clknet_leaf_90_u_dsync.out_clk ),
    .D(_1113_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8641_ (.CLK(\clknet_leaf_70_u_dsync.out_clk ),
    .D(_1114_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8642_ (.CLK(\clknet_leaf_70_u_dsync.out_clk ),
    .D(_1115_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8643_ (.CLK(\clknet_leaf_69_u_dsync.out_clk ),
    .D(_1116_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8644_ (.CLK(\clknet_leaf_93_u_dsync.out_clk ),
    .D(_1117_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8645_ (.CLK(\clknet_leaf_92_u_dsync.out_clk ),
    .D(_1118_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8646_ (.CLK(\clknet_leaf_93_u_dsync.out_clk ),
    .D(_1119_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8647_ (.CLK(\clknet_leaf_93_u_dsync.out_clk ),
    .D(_1120_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8648_ (.CLK(\clknet_leaf_86_u_dsync.out_clk ),
    .D(_1121_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8649_ (.CLK(\clknet_leaf_93_u_dsync.out_clk ),
    .D(_1122_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8650_ (.CLK(\clknet_leaf_93_u_dsync.out_clk ),
    .D(_1123_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8651_ (.CLK(\clknet_leaf_94_u_dsync.out_clk ),
    .D(_1124_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8652_ (.CLK(\clknet_leaf_94_u_dsync.out_clk ),
    .D(_1125_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8653_ (.CLK(\clknet_leaf_89_u_dsync.out_clk ),
    .D(_1126_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8654_ (.CLK(\clknet_leaf_87_u_dsync.out_clk ),
    .D(_1127_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8655_ (.CLK(\clknet_leaf_95_u_dsync.out_clk ),
    .D(_1128_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][32] ));
 sky130_fd_sc_hd__dfxtp_1 _8656_ (.CLK(\clknet_leaf_92_u_dsync.out_clk ),
    .D(_1129_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][33] ));
 sky130_fd_sc_hd__dfxtp_1 _8657_ (.CLK(\clknet_leaf_87_u_dsync.out_clk ),
    .D(_1130_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][34] ));
 sky130_fd_sc_hd__dfxtp_1 _8658_ (.CLK(\clknet_leaf_94_u_dsync.out_clk ),
    .D(_1131_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][35] ));
 sky130_fd_sc_hd__dfxtp_1 _8659_ (.CLK(\clknet_leaf_89_u_dsync.out_clk ),
    .D(_1132_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][36] ));
 sky130_fd_sc_hd__dfxtp_1 _8660_ (.CLK(\clknet_leaf_91_u_dsync.out_clk ),
    .D(_1133_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][37] ));
 sky130_fd_sc_hd__dfxtp_1 _8661_ (.CLK(\clknet_leaf_88_u_dsync.out_clk ),
    .D(_1134_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][38] ));
 sky130_fd_sc_hd__dfxtp_1 _8662_ (.CLK(\clknet_leaf_92_u_dsync.out_clk ),
    .D(_1135_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][39] ));
 sky130_fd_sc_hd__dfxtp_1 _8663_ (.CLK(\clknet_leaf_89_u_dsync.out_clk ),
    .D(_1136_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][40] ));
 sky130_fd_sc_hd__dfxtp_1 _8664_ (.CLK(\clknet_leaf_94_u_dsync.out_clk ),
    .D(_1137_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][41] ));
 sky130_fd_sc_hd__dfxtp_1 _8665_ (.CLK(\clknet_leaf_91_u_dsync.out_clk ),
    .D(_1138_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][42] ));
 sky130_fd_sc_hd__dfxtp_1 _8666_ (.CLK(\clknet_leaf_91_u_dsync.out_clk ),
    .D(_1139_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][43] ));
 sky130_fd_sc_hd__dfxtp_1 _8667_ (.CLK(\clknet_leaf_90_u_dsync.out_clk ),
    .D(_1140_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][44] ));
 sky130_fd_sc_hd__dfxtp_1 _8668_ (.CLK(\clknet_leaf_101_u_dsync.out_clk ),
    .D(_1141_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][45] ));
 sky130_fd_sc_hd__dfxtp_1 _8669_ (.CLK(\clknet_leaf_89_u_dsync.out_clk ),
    .D(_1142_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][46] ));
 sky130_fd_sc_hd__dfxtp_1 _8670_ (.CLK(\clknet_leaf_92_u_dsync.out_clk ),
    .D(_1143_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][47] ));
 sky130_fd_sc_hd__dfxtp_1 _8671_ (.CLK(\clknet_leaf_91_u_dsync.out_clk ),
    .D(_1144_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][48] ));
 sky130_fd_sc_hd__dfxtp_1 _8672_ (.CLK(\clknet_leaf_90_u_dsync.out_clk ),
    .D(_1145_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][49] ));
 sky130_fd_sc_hd__dfxtp_1 _8673_ (.CLK(\clknet_leaf_101_u_dsync.out_clk ),
    .D(_1146_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][50] ));
 sky130_fd_sc_hd__dfxtp_1 _8674_ (.CLK(\clknet_leaf_106_u_dsync.out_clk ),
    .D(_1147_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][53] ));
 sky130_fd_sc_hd__dfxtp_1 _8675_ (.CLK(\clknet_leaf_106_u_dsync.out_clk ),
    .D(_1148_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][54] ));
 sky130_fd_sc_hd__dfxtp_1 _8676_ (.CLK(\clknet_leaf_101_u_dsync.out_clk ),
    .D(_1149_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][55] ));
 sky130_fd_sc_hd__dfxtp_1 _8677_ (.CLK(\clknet_leaf_100_u_dsync.out_clk ),
    .D(_1150_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][56] ));
 sky130_fd_sc_hd__dfxtp_1 _8678_ (.CLK(\clknet_leaf_102_u_dsync.out_clk ),
    .D(_1151_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][57] ));
 sky130_fd_sc_hd__dfxtp_1 _8679_ (.CLK(\clknet_leaf_88_u_dsync.out_clk ),
    .D(_1152_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][58] ));
 sky130_fd_sc_hd__dfxtp_1 _8680_ (.CLK(\clknet_leaf_100_u_dsync.out_clk ),
    .D(_1153_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][59] ));
 sky130_fd_sc_hd__dfxtp_1 _8681_ (.CLK(\clknet_leaf_105_u_dsync.out_clk ),
    .D(_1154_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][60] ));
 sky130_fd_sc_hd__dfxtp_1 _8682_ (.CLK(\clknet_leaf_106_u_dsync.out_clk ),
    .D(_1155_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][61] ));
 sky130_fd_sc_hd__dfxtp_1 _8683_ (.CLK(\clknet_leaf_107_u_dsync.out_clk ),
    .D(_1156_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][62] ));
 sky130_fd_sc_hd__dfxtp_1 _8684_ (.CLK(\clknet_leaf_107_u_dsync.out_clk ),
    .D(_1157_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][63] ));
 sky130_fd_sc_hd__dfxtp_1 _8685_ (.CLK(\clknet_leaf_107_u_dsync.out_clk ),
    .D(_1158_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][64] ));
 sky130_fd_sc_hd__dfxtp_1 _8686_ (.CLK(\clknet_leaf_108_u_dsync.out_clk ),
    .D(_1159_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][65] ));
 sky130_fd_sc_hd__dfxtp_1 _8687_ (.CLK(\clknet_leaf_108_u_dsync.out_clk ),
    .D(_1160_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][66] ));
 sky130_fd_sc_hd__dfxtp_1 _8688_ (.CLK(\clknet_leaf_102_u_dsync.out_clk ),
    .D(_1161_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][67] ));
 sky130_fd_sc_hd__dfxtp_1 _8689_ (.CLK(\clknet_leaf_102_u_dsync.out_clk ),
    .D(_1162_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][68] ));
 sky130_fd_sc_hd__dfxtp_1 _8690_ (.CLK(\clknet_leaf_103_u_dsync.out_clk ),
    .D(_1163_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][69] ));
 sky130_fd_sc_hd__dfxtp_1 _8691_ (.CLK(\clknet_leaf_90_u_dsync.out_clk ),
    .D(_1164_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][70] ));
 sky130_fd_sc_hd__dfxtp_1 _8692_ (.CLK(\clknet_leaf_105_u_dsync.out_clk ),
    .D(_1165_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][71] ));
 sky130_fd_sc_hd__dfxtp_1 _8693_ (.CLK(\clknet_leaf_104_u_dsync.out_clk ),
    .D(_1166_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][72] ));
 sky130_fd_sc_hd__dfxtp_1 _8694_ (.CLK(\clknet_leaf_104_u_dsync.out_clk ),
    .D(_1167_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][73] ));
 sky130_fd_sc_hd__dfxtp_1 _8695_ (.CLK(\clknet_leaf_103_u_dsync.out_clk ),
    .D(_1168_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][74] ));
 sky130_fd_sc_hd__dfxtp_1 _8696_ (.CLK(\clknet_leaf_104_u_dsync.out_clk ),
    .D(_1169_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][75] ));
 sky130_fd_sc_hd__dfxtp_1 _8697_ (.CLK(\clknet_leaf_104_u_dsync.out_clk ),
    .D(_1170_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][76] ));
 sky130_fd_sc_hd__dfxtp_1 _8698_ (.CLK(\clknet_leaf_104_u_dsync.out_clk ),
    .D(_1171_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][77] ));
 sky130_fd_sc_hd__dfxtp_1 _8699_ (.CLK(\clknet_leaf_104_u_dsync.out_clk ),
    .D(_1172_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][78] ));
 sky130_fd_sc_hd__dfxtp_1 _8700_ (.CLK(\clknet_leaf_103_u_dsync.out_clk ),
    .D(_1173_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][79] ));
 sky130_fd_sc_hd__dfxtp_1 _8701_ (.CLK(\clknet_leaf_105_u_dsync.out_clk ),
    .D(_1174_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][80] ));
 sky130_fd_sc_hd__dfxtp_1 _8702_ (.CLK(\clknet_leaf_108_u_dsync.out_clk ),
    .D(_1175_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][81] ));
 sky130_fd_sc_hd__dfxtp_1 _8703_ (.CLK(\clknet_leaf_103_u_dsync.out_clk ),
    .D(_1176_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[3][82] ));
 sky130_fd_sc_hd__dfxtp_1 _8704_ (.CLK(\clknet_leaf_28_u_dsync.out_clk ),
    .D(_1177_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8705_ (.CLK(\clknet_leaf_28_u_dsync.out_clk ),
    .D(_1178_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8706_ (.CLK(\clknet_leaf_29_u_dsync.out_clk ),
    .D(_1179_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8707_ (.CLK(\clknet_leaf_25_u_dsync.out_clk ),
    .D(_1180_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8708_ (.CLK(\clknet_leaf_11_u_dsync.out_clk ),
    .D(_1181_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8709_ (.CLK(\clknet_leaf_28_u_dsync.out_clk ),
    .D(_1182_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8710_ (.CLK(\clknet_leaf_35_u_dsync.out_clk ),
    .D(_1183_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8711_ (.CLK(\clknet_leaf_34_u_dsync.out_clk ),
    .D(_1184_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8712_ (.CLK(\clknet_leaf_27_u_dsync.out_clk ),
    .D(_1185_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8713_ (.CLK(\clknet_leaf_31_u_dsync.out_clk ),
    .D(_1186_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8714_ (.CLK(\clknet_leaf_30_u_dsync.out_clk ),
    .D(_1187_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8715_ (.CLK(\clknet_leaf_32_u_dsync.out_clk ),
    .D(_1188_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8716_ (.CLK(\clknet_leaf_36_u_dsync.out_clk ),
    .D(_1189_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8717_ (.CLK(\clknet_leaf_43_u_dsync.out_clk ),
    .D(_1190_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8718_ (.CLK(\clknet_leaf_40_u_dsync.out_clk ),
    .D(_1191_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8719_ (.CLK(\clknet_leaf_46_u_dsync.out_clk ),
    .D(_1192_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8720_ (.CLK(\clknet_leaf_42_u_dsync.out_clk ),
    .D(_1193_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8721_ (.CLK(\clknet_leaf_46_u_dsync.out_clk ),
    .D(_1194_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8722_ (.CLK(\clknet_leaf_40_u_dsync.out_clk ),
    .D(_1195_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8723_ (.CLK(\clknet_leaf_43_u_dsync.out_clk ),
    .D(_1196_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8724_ (.CLK(\clknet_leaf_46_u_dsync.out_clk ),
    .D(_1197_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8725_ (.CLK(\clknet_leaf_41_u_dsync.out_clk ),
    .D(_1198_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8726_ (.CLK(\clknet_leaf_44_u_dsync.out_clk ),
    .D(_1199_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8727_ (.CLK(\clknet_leaf_45_u_dsync.out_clk ),
    .D(_1200_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8728_ (.CLK(\clknet_leaf_40_u_dsync.out_clk ),
    .D(_1201_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8729_ (.CLK(\clknet_leaf_44_u_dsync.out_clk ),
    .D(_1202_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8730_ (.CLK(\clknet_leaf_40_u_dsync.out_clk ),
    .D(_1203_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8731_ (.CLK(\clknet_leaf_44_u_dsync.out_clk ),
    .D(_1204_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _8732_ (.CLK(\clknet_leaf_44_u_dsync.out_clk ),
    .D(_1205_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _8733_ (.CLK(\clknet_leaf_45_u_dsync.out_clk ),
    .D(_1206_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _8734_ (.CLK(\clknet_leaf_32_u_dsync.out_clk ),
    .D(_1207_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _8735_ (.CLK(\clknet_leaf_45_u_dsync.out_clk ),
    .D(_1208_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _8736_ (.CLK(\clknet_leaf_31_u_dsync.out_clk ),
    .D(_1209_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _8737_ (.CLK(\clknet_leaf_40_u_dsync.out_clk ),
    .D(_1210_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _8738_ (.CLK(\clknet_leaf_41_u_dsync.out_clk ),
    .D(_1211_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _8739_ (.CLK(\clknet_leaf_44_u_dsync.out_clk ),
    .D(_1212_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _8740_ (.CLK(\clknet_leaf_39_u_dsync.out_clk ),
    .D(_1213_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _8741_ (.CLK(\clknet_leaf_36_u_dsync.out_clk ),
    .D(_1214_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _8742_ (.CLK(\clknet_leaf_33_u_dsync.out_clk ),
    .D(_1215_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _8743_ (.CLK(\clknet_leaf_46_u_dsync.out_clk ),
    .D(_1216_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _8744_ (.CLK(\clknet_leaf_31_u_dsync.out_clk ),
    .D(_1217_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _8745_ (.CLK(\clknet_leaf_36_u_dsync.out_clk ),
    .D(_1218_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _8746_ (.CLK(\clknet_leaf_36_u_dsync.out_clk ),
    .D(_1219_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][47] ));
 sky130_fd_sc_hd__dfxtp_1 _8747_ (.CLK(\clknet_leaf_33_u_dsync.out_clk ),
    .D(_1220_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][48] ));
 sky130_fd_sc_hd__dfxtp_1 _8748_ (.CLK(\clknet_leaf_36_u_dsync.out_clk ),
    .D(_1221_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][49] ));
 sky130_fd_sc_hd__dfxtp_1 _8749_ (.CLK(\clknet_leaf_31_u_dsync.out_clk ),
    .D(_1222_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][50] ));
 sky130_fd_sc_hd__dfxtp_1 _8750_ (.CLK(\clknet_leaf_33_u_dsync.out_clk ),
    .D(_1223_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][53] ));
 sky130_fd_sc_hd__dfxtp_1 _8751_ (.CLK(\clknet_leaf_34_u_dsync.out_clk ),
    .D(_1224_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][54] ));
 sky130_fd_sc_hd__dfxtp_1 _8752_ (.CLK(\clknet_leaf_36_u_dsync.out_clk ),
    .D(_1225_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][55] ));
 sky130_fd_sc_hd__dfxtp_1 _8753_ (.CLK(\clknet_leaf_36_u_dsync.out_clk ),
    .D(_1226_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][56] ));
 sky130_fd_sc_hd__dfxtp_1 _8754_ (.CLK(\clknet_leaf_34_u_dsync.out_clk ),
    .D(_1227_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][57] ));
 sky130_fd_sc_hd__dfxtp_1 _8755_ (.CLK(\clknet_leaf_35_u_dsync.out_clk ),
    .D(_1228_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][58] ));
 sky130_fd_sc_hd__dfxtp_1 _8756_ (.CLK(\clknet_leaf_33_u_dsync.out_clk ),
    .D(_1229_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][59] ));
 sky130_fd_sc_hd__dfxtp_1 _8757_ (.CLK(\clknet_leaf_35_u_dsync.out_clk ),
    .D(_1230_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][60] ));
 sky130_fd_sc_hd__dfxtp_1 _8758_ (.CLK(\clknet_leaf_35_u_dsync.out_clk ),
    .D(_1231_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[2][61] ));
 sky130_fd_sc_hd__dfstp_2 _8759_ (.CLK(\clknet_leaf_35_u_dsync.out_clk ),
    .D(_0006_),
    .SET_B(net890),
    .Q(\u_s2.u_sync_wbb.m_state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _8760_ (.CLK(\clknet_leaf_35_u_dsync.out_clk ),
    .D(_0007_),
    .RESET_B(net890),
    .Q(\u_s2.u_sync_wbb.m_state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _8761_ (.CLK(\clknet_leaf_35_u_dsync.out_clk ),
    .D(_0008_),
    .RESET_B(net890),
    .Q(\u_s2.u_sync_wbb.m_state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8762_ (.CLK(net1743),
    .D(net1731),
    .RESET_B(rst_n),
    .Q(\u_rst_sync.in_data_s ));
 sky130_fd_sc_hd__conb_1 _8762__1731 (.HI(net1731));
 sky130_fd_sc_hd__dfrtp_1 _8763_ (.CLK(\clknet_leaf_109_u_dsync.out_clk ),
    .D(\u_rst_sync.in_data_s ),
    .RESET_B(rst_n),
    .Q(\u_rst_sync.in_data_2s ));
 sky130_fd_sc_hd__dfxtp_1 _8764_ (.CLK(\clknet_leaf_7_u_dsync.out_clk ),
    .D(_1232_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8765_ (.CLK(\clknet_leaf_6_u_dsync.out_clk ),
    .D(_1233_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8766_ (.CLK(\clknet_leaf_7_u_dsync.out_clk ),
    .D(_1234_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8767_ (.CLK(\clknet_leaf_6_u_dsync.out_clk ),
    .D(_1235_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8768_ (.CLK(\clknet_leaf_10_u_dsync.out_clk ),
    .D(_1236_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8769_ (.CLK(\clknet_leaf_10_u_dsync.out_clk ),
    .D(_1237_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8770_ (.CLK(\clknet_leaf_6_u_dsync.out_clk ),
    .D(_1238_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8771_ (.CLK(\clknet_leaf_10_u_dsync.out_clk ),
    .D(_1239_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8772_ (.CLK(\clknet_leaf_6_u_dsync.out_clk ),
    .D(_1240_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8773_ (.CLK(\clknet_leaf_37_u_dsync.out_clk ),
    .D(_1241_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8774_ (.CLK(\clknet_leaf_8_u_dsync.out_clk ),
    .D(_1242_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8775_ (.CLK(\clknet_leaf_8_u_dsync.out_clk ),
    .D(_1243_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8776_ (.CLK(\clknet_leaf_9_u_dsync.out_clk ),
    .D(_1244_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8777_ (.CLK(\clknet_leaf_63_u_dsync.out_clk ),
    .D(_1245_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8778_ (.CLK(\clknet_leaf_65_u_dsync.out_clk ),
    .D(_1246_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8779_ (.CLK(\clknet_leaf_65_u_dsync.out_clk ),
    .D(_1247_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8780_ (.CLK(\clknet_leaf_66_u_dsync.out_clk ),
    .D(_1248_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8781_ (.CLK(\clknet_leaf_39_u_dsync.out_clk ),
    .D(_1249_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8782_ (.CLK(\clknet_leaf_65_u_dsync.out_clk ),
    .D(_1250_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8783_ (.CLK(\clknet_leaf_67_u_dsync.out_clk ),
    .D(_1251_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8784_ (.CLK(\clknet_leaf_39_u_dsync.out_clk ),
    .D(_1252_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8785_ (.CLK(\clknet_leaf_65_u_dsync.out_clk ),
    .D(_1253_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8786_ (.CLK(\clknet_leaf_63_u_dsync.out_clk ),
    .D(_1254_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8787_ (.CLK(\clknet_leaf_41_u_dsync.out_clk ),
    .D(_1255_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8788_ (.CLK(\clknet_leaf_39_u_dsync.out_clk ),
    .D(_1256_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8789_ (.CLK(\clknet_leaf_39_u_dsync.out_clk ),
    .D(_1257_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8790_ (.CLK(\clknet_leaf_66_u_dsync.out_clk ),
    .D(_1258_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8791_ (.CLK(\clknet_leaf_38_u_dsync.out_clk ),
    .D(_1259_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _8792_ (.CLK(\clknet_leaf_68_u_dsync.out_clk ),
    .D(_1260_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _8793_ (.CLK(\clknet_leaf_66_u_dsync.out_clk ),
    .D(_1261_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _8794_ (.CLK(\clknet_leaf_38_u_dsync.out_clk ),
    .D(_1262_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _8795_ (.CLK(\clknet_leaf_67_u_dsync.out_clk ),
    .D(_1263_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _8796_ (.CLK(\clknet_leaf_38_u_dsync.out_clk ),
    .D(_1264_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _8797_ (.CLK(\clknet_leaf_66_u_dsync.out_clk ),
    .D(_1265_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _8798_ (.CLK(\clknet_leaf_69_u_dsync.out_clk ),
    .D(_1266_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _8799_ (.CLK(\clknet_leaf_66_u_dsync.out_clk ),
    .D(_1267_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _8800_ (.CLK(\clknet_leaf_66_u_dsync.out_clk ),
    .D(_1268_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _8801_ (.CLK(\clknet_leaf_38_u_dsync.out_clk ),
    .D(_1269_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _8802_ (.CLK(\clknet_leaf_66_u_dsync.out_clk ),
    .D(_1270_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _8803_ (.CLK(\clknet_leaf_95_u_dsync.out_clk ),
    .D(_1271_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _8804_ (.CLK(\clknet_leaf_37_u_dsync.out_clk ),
    .D(_1272_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _8805_ (.CLK(\clknet_leaf_37_u_dsync.out_clk ),
    .D(_1273_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _8806_ (.CLK(\clknet_leaf_68_u_dsync.out_clk ),
    .D(_1274_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][47] ));
 sky130_fd_sc_hd__dfxtp_1 _8807_ (.CLK(\clknet_leaf_95_u_dsync.out_clk ),
    .D(_1275_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][48] ));
 sky130_fd_sc_hd__dfxtp_1 _8808_ (.CLK(\clknet_leaf_67_u_dsync.out_clk ),
    .D(_1276_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][49] ));
 sky130_fd_sc_hd__dfxtp_1 _8809_ (.CLK(\clknet_leaf_9_u_dsync.out_clk ),
    .D(_1277_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][50] ));
 sky130_fd_sc_hd__dfxtp_1 _8810_ (.CLK(\clknet_leaf_8_u_dsync.out_clk ),
    .D(_1278_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][53] ));
 sky130_fd_sc_hd__dfxtp_1 _8811_ (.CLK(\clknet_leaf_8_u_dsync.out_clk ),
    .D(_1279_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][54] ));
 sky130_fd_sc_hd__dfxtp_1 _8812_ (.CLK(\clknet_leaf_7_u_dsync.out_clk ),
    .D(_1280_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][55] ));
 sky130_fd_sc_hd__dfxtp_1 _8813_ (.CLK(\clknet_leaf_7_u_dsync.out_clk ),
    .D(_1281_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][56] ));
 sky130_fd_sc_hd__dfxtp_1 _8814_ (.CLK(\clknet_leaf_96_u_dsync.out_clk ),
    .D(_1282_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][57] ));
 sky130_fd_sc_hd__dfxtp_1 _8815_ (.CLK(\clknet_leaf_8_u_dsync.out_clk ),
    .D(_1283_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][58] ));
 sky130_fd_sc_hd__dfxtp_1 _8816_ (.CLK(\clknet_leaf_8_u_dsync.out_clk ),
    .D(_1284_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[2][59] ));
 sky130_fd_sc_hd__dfrtp_1 _8817_ (.CLK(\clknet_leaf_22_u_dsync.out_clk ),
    .D(_1285_),
    .RESET_B(net906),
    .Q(\u_reg.reg_7[24] ));
 sky130_fd_sc_hd__dfrtp_1 _8818_ (.CLK(\clknet_leaf_24_u_dsync.out_clk ),
    .D(_1286_),
    .RESET_B(net907),
    .Q(\u_reg.reg_7[25] ));
 sky130_fd_sc_hd__dfrtp_1 _8819_ (.CLK(\clknet_leaf_21_u_dsync.out_clk ),
    .D(_1287_),
    .RESET_B(net894),
    .Q(\u_reg.reg_7[26] ));
 sky130_fd_sc_hd__dfrtp_1 _8820_ (.CLK(\clknet_leaf_24_u_dsync.out_clk ),
    .D(_1288_),
    .RESET_B(net907),
    .Q(\u_reg.reg_7[27] ));
 sky130_fd_sc_hd__dfrtp_1 _8821_ (.CLK(\clknet_leaf_18_u_dsync.out_clk ),
    .D(_1289_),
    .RESET_B(net888),
    .Q(\u_reg.reg_7[28] ));
 sky130_fd_sc_hd__dfrtp_1 _8822_ (.CLK(\clknet_leaf_21_u_dsync.out_clk ),
    .D(_1290_),
    .RESET_B(net895),
    .Q(\u_reg.reg_7[29] ));
 sky130_fd_sc_hd__dfrtp_1 _8823_ (.CLK(\clknet_leaf_23_u_dsync.out_clk ),
    .D(_1291_),
    .RESET_B(net911),
    .Q(\u_reg.reg_7[30] ));
 sky130_fd_sc_hd__dfrtp_1 _8824_ (.CLK(\clknet_leaf_17_u_dsync.out_clk ),
    .D(_1292_),
    .RESET_B(net883),
    .Q(\u_reg.reg_7[31] ));
 sky130_fd_sc_hd__dfrtp_4 _8825_ (.CLK(\clknet_leaf_100_u_dsync.out_clk ),
    .D(_1293_),
    .RESET_B(net840),
    .Q(\u_s0.u_sync_wbb.wbm_ack_o ));
 sky130_fd_sc_hd__dfrtp_4 _8826_ (.CLK(\clknet_leaf_100_u_dsync.out_clk ),
    .D(_1294_),
    .RESET_B(net840),
    .Q(\u_s0.u_sync_wbb.wbm_lack_o ));
 sky130_fd_sc_hd__dfrtp_4 _8827_ (.CLK(\clknet_leaf_98_u_dsync.out_clk ),
    .D(_1295_),
    .RESET_B(net847),
    .Q(\u_s0.u_sync_wbb.m_cmd_wr_en ));
 sky130_fd_sc_hd__dfrtp_4 _8828_ (.CLK(\clknet_leaf_98_u_dsync.out_clk ),
    .D(_1296_),
    .RESET_B(net853),
    .Q(\u_s0.u_sync_wbb.m_resp_rd_en ));
 sky130_fd_sc_hd__dfrtp_4 _8829_ (.CLK(\clknet_leaf_13_u_dsync.out_clk ),
    .D(_1297_),
    .RESET_B(net877),
    .Q(\u_s1.u_sync_wbb.m_bl_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_2 _8830_ (.CLK(\clknet_leaf_12_u_dsync.out_clk ),
    .D(_1298_),
    .RESET_B(net881),
    .Q(\u_s1.u_sync_wbb.m_bl_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_4 _8831_ (.CLK(\clknet_leaf_12_u_dsync.out_clk ),
    .D(_1299_),
    .RESET_B(net890),
    .Q(\u_s1.u_sync_wbb.m_bl_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8832_ (.CLK(\clknet_leaf_12_u_dsync.out_clk ),
    .D(_1300_),
    .RESET_B(net885),
    .Q(\u_s1.u_sync_wbb.m_bl_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_2 _8833_ (.CLK(\clknet_leaf_11_u_dsync.out_clk ),
    .D(_1301_),
    .RESET_B(net885),
    .Q(\u_s1.u_sync_wbb.m_bl_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_2 _8834_ (.CLK(\clknet_leaf_11_u_dsync.out_clk ),
    .D(_1302_),
    .RESET_B(net885),
    .Q(\u_s1.u_sync_wbb.m_bl_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _8835_ (.CLK(\clknet_leaf_14_u_dsync.out_clk ),
    .D(_1303_),
    .RESET_B(net872),
    .Q(\u_s1.u_sync_wbb.m_bl_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _8836_ (.CLK(\clknet_leaf_5_u_dsync.out_clk ),
    .D(_1304_),
    .RESET_B(net855),
    .Q(\u_s1.u_sync_wbb.m_bl_cnt[7] ));
 sky130_fd_sc_hd__dfrtp_2 _8837_ (.CLK(\clknet_leaf_6_u_dsync.out_clk ),
    .D(_1305_),
    .RESET_B(net857),
    .Q(\u_s1.u_sync_wbb.m_bl_cnt[8] ));
 sky130_fd_sc_hd__dfrtp_1 _8838_ (.CLK(\clknet_leaf_5_u_dsync.out_clk ),
    .D(_1306_),
    .RESET_B(net858),
    .Q(\u_s1.u_sync_wbb.m_bl_cnt[9] ));
 sky130_fd_sc_hd__dfrtp_1 _8839_ (.CLK(\clknet_leaf_81_u_dsync.out_clk ),
    .D(s0_wbd_lack_i),
    .RESET_B(net836),
    .Q(\u_s0.u_sync_wbb.wbs_ack_f ));
 sky130_fd_sc_hd__dfrtp_1 _8840_ (.CLK(\clknet_leaf_81_u_dsync.out_clk ),
    .D(net342),
    .RESET_B(net835),
    .Q(\u_s0.u_sync_wbb.wbs_stb_l ));
 sky130_fd_sc_hd__dfrtp_4 _8841_ (.CLK(\clknet_leaf_78_u_dsync.out_clk ),
    .D(_1307_),
    .RESET_B(net844),
    .Q(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_2 _8842_ (.CLK(\clknet_leaf_77_u_dsync.out_clk ),
    .D(_1308_),
    .RESET_B(net851),
    .Q(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_2 _8843_ (.CLK(\clknet_leaf_70_u_dsync.out_clk ),
    .D(_1309_),
    .RESET_B(net853),
    .Q(\u_s0.u_sync_wbb.u_resp_if.wr_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_4 _8844_ (.CLK(\clknet_leaf_96_u_dsync.out_clk ),
    .D(_1310_),
    .RESET_B(net862),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_4 _8845_ (.CLK(\clknet_leaf_97_u_dsync.out_clk ),
    .D(_1311_),
    .RESET_B(net850),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_4 _8846_ (.CLK(\clknet_leaf_94_u_dsync.out_clk ),
    .D(_1312_),
    .RESET_B(net852),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.wr_ptr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8847_ (.CLK(\clknet_leaf_28_u_dsync.out_clk ),
    .D(_1313_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8848_ (.CLK(\clknet_leaf_28_u_dsync.out_clk ),
    .D(_1314_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8849_ (.CLK(\clknet_leaf_28_u_dsync.out_clk ),
    .D(_1315_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8850_ (.CLK(\clknet_leaf_29_u_dsync.out_clk ),
    .D(_1316_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8851_ (.CLK(\clknet_leaf_11_u_dsync.out_clk ),
    .D(_1317_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8852_ (.CLK(\clknet_leaf_28_u_dsync.out_clk ),
    .D(_1318_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8853_ (.CLK(\clknet_leaf_35_u_dsync.out_clk ),
    .D(_1319_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8854_ (.CLK(\clknet_leaf_34_u_dsync.out_clk ),
    .D(_1320_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8855_ (.CLK(\clknet_leaf_27_u_dsync.out_clk ),
    .D(_1321_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8856_ (.CLK(\clknet_leaf_31_u_dsync.out_clk ),
    .D(_1322_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8857_ (.CLK(\clknet_leaf_30_u_dsync.out_clk ),
    .D(_1323_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8858_ (.CLK(\clknet_leaf_32_u_dsync.out_clk ),
    .D(_1324_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8859_ (.CLK(\clknet_leaf_36_u_dsync.out_clk ),
    .D(_1325_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8860_ (.CLK(\clknet_leaf_42_u_dsync.out_clk ),
    .D(_1326_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8861_ (.CLK(\clknet_leaf_42_u_dsync.out_clk ),
    .D(_1327_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8862_ (.CLK(\clknet_leaf_46_u_dsync.out_clk ),
    .D(_1328_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8863_ (.CLK(\clknet_leaf_49_u_dsync.out_clk ),
    .D(_1329_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8864_ (.CLK(\clknet_leaf_47_u_dsync.out_clk ),
    .D(_1330_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8865_ (.CLK(\clknet_leaf_43_u_dsync.out_clk ),
    .D(_1331_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8866_ (.CLK(\clknet_leaf_43_u_dsync.out_clk ),
    .D(_1332_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8867_ (.CLK(\clknet_leaf_45_u_dsync.out_clk ),
    .D(_1333_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8868_ (.CLK(\clknet_leaf_41_u_dsync.out_clk ),
    .D(_1334_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8869_ (.CLK(\clknet_leaf_44_u_dsync.out_clk ),
    .D(_1335_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8870_ (.CLK(\clknet_leaf_45_u_dsync.out_clk ),
    .D(_1336_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8871_ (.CLK(\clknet_leaf_40_u_dsync.out_clk ),
    .D(_1337_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8872_ (.CLK(\clknet_leaf_44_u_dsync.out_clk ),
    .D(_1338_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8873_ (.CLK(\clknet_leaf_40_u_dsync.out_clk ),
    .D(_1339_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _8874_ (.CLK(\clknet_leaf_45_u_dsync.out_clk ),
    .D(_1340_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _8875_ (.CLK(\clknet_leaf_43_u_dsync.out_clk ),
    .D(_1341_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _8876_ (.CLK(\clknet_leaf_45_u_dsync.out_clk ),
    .D(_1342_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _8877_ (.CLK(\clknet_leaf_31_u_dsync.out_clk ),
    .D(_1343_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _8878_ (.CLK(\clknet_leaf_45_u_dsync.out_clk ),
    .D(_1344_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _8879_ (.CLK(\clknet_leaf_31_u_dsync.out_clk ),
    .D(_1345_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _8880_ (.CLK(\clknet_leaf_40_u_dsync.out_clk ),
    .D(_1346_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _8881_ (.CLK(\clknet_leaf_63_u_dsync.out_clk ),
    .D(_1347_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _8882_ (.CLK(\clknet_leaf_40_u_dsync.out_clk ),
    .D(_1348_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _8883_ (.CLK(\clknet_leaf_39_u_dsync.out_clk ),
    .D(_1349_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _8884_ (.CLK(\clknet_leaf_40_u_dsync.out_clk ),
    .D(_1350_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _8885_ (.CLK(\clknet_leaf_33_u_dsync.out_clk ),
    .D(_1351_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _8886_ (.CLK(\clknet_leaf_46_u_dsync.out_clk ),
    .D(_1352_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _8887_ (.CLK(\clknet_leaf_32_u_dsync.out_clk ),
    .D(_1353_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _8888_ (.CLK(\clknet_leaf_36_u_dsync.out_clk ),
    .D(_1354_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _8889_ (.CLK(\clknet_leaf_37_u_dsync.out_clk ),
    .D(_1355_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][47] ));
 sky130_fd_sc_hd__dfxtp_1 _8890_ (.CLK(\clknet_leaf_32_u_dsync.out_clk ),
    .D(_1356_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][48] ));
 sky130_fd_sc_hd__dfxtp_1 _8891_ (.CLK(\clknet_leaf_36_u_dsync.out_clk ),
    .D(_1357_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][49] ));
 sky130_fd_sc_hd__dfxtp_1 _8892_ (.CLK(\clknet_leaf_32_u_dsync.out_clk ),
    .D(_1358_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][50] ));
 sky130_fd_sc_hd__dfxtp_1 _8893_ (.CLK(\clknet_leaf_33_u_dsync.out_clk ),
    .D(_1359_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][53] ));
 sky130_fd_sc_hd__dfxtp_1 _8894_ (.CLK(\clknet_leaf_28_u_dsync.out_clk ),
    .D(_1360_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][54] ));
 sky130_fd_sc_hd__dfxtp_1 _8895_ (.CLK(\clknet_leaf_33_u_dsync.out_clk ),
    .D(_1361_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][55] ));
 sky130_fd_sc_hd__dfxtp_1 _8896_ (.CLK(\clknet_leaf_33_u_dsync.out_clk ),
    .D(_1362_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][56] ));
 sky130_fd_sc_hd__dfxtp_1 _8897_ (.CLK(\clknet_leaf_34_u_dsync.out_clk ),
    .D(_1363_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][57] ));
 sky130_fd_sc_hd__dfxtp_1 _8898_ (.CLK(\clknet_leaf_35_u_dsync.out_clk ),
    .D(_1364_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][58] ));
 sky130_fd_sc_hd__dfxtp_1 _8899_ (.CLK(\clknet_leaf_32_u_dsync.out_clk ),
    .D(_1365_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][59] ));
 sky130_fd_sc_hd__dfxtp_1 _8900_ (.CLK(\clknet_leaf_35_u_dsync.out_clk ),
    .D(_1366_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][60] ));
 sky130_fd_sc_hd__dfxtp_1 _8901_ (.CLK(\clknet_leaf_35_u_dsync.out_clk ),
    .D(_1367_),
    .Q(\u_s2.u_sync_wbb.u_cmd_if.mem[1][61] ));
 sky130_fd_sc_hd__dfrtp_1 _8902_ (.CLK(\clknet_leaf_82_u_dsync.out_clk ),
    .D(_1368_),
    .RESET_B(net838),
    .Q(\u_s0.u_sync_wbb.wbs_burst ));
 sky130_fd_sc_hd__dfrtp_1 _8903_ (.CLK(\clknet_leaf_86_u_dsync.out_clk ),
    .D(_1369_),
    .RESET_B(net842),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8904_ (.CLK(\clknet_leaf_94_u_dsync.out_clk ),
    .D(_1370_),
    .RESET_B(net851),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8905_ (.CLK(\clknet_leaf_94_u_dsync.out_clk ),
    .D(_1371_),
    .RESET_B(net851),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.rd_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8906_ (.CLK(\clknet_leaf_77_u_dsync.out_clk ),
    .D(_1372_),
    .RESET_B(net851),
    .Q(\u_s0.u_sync_wbb.u_resp_if.rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8907_ (.CLK(\clknet_leaf_77_u_dsync.out_clk ),
    .D(_1373_),
    .RESET_B(net851),
    .Q(\u_s0.u_sync_wbb.u_resp_if.rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_2 _8908_ (.CLK(\clknet_leaf_70_u_dsync.out_clk ),
    .D(_1374_),
    .RESET_B(net852),
    .Q(\u_s0.u_sync_wbb.u_resp_if.rd_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8909_ (.CLK(\clknet_leaf_5_u_dsync.out_clk ),
    .D(_1375_),
    .RESET_B(net849),
    .Q(\u_reg.reg_rdata[0] ));
 sky130_fd_sc_hd__dfrtp_4 _8910_ (.CLK(\clknet_leaf_107_u_dsync.out_clk ),
    .D(_1376_),
    .RESET_B(net841),
    .Q(\u_reg.reg_rdata[1] ));
 sky130_fd_sc_hd__dfrtp_4 _8911_ (.CLK(\clknet_leaf_0_u_dsync.out_clk ),
    .D(_1377_),
    .RESET_B(net840),
    .Q(\u_reg.reg_rdata[2] ));
 sky130_fd_sc_hd__dfrtp_4 _8912_ (.CLK(\clknet_leaf_1_u_dsync.out_clk ),
    .D(_1378_),
    .RESET_B(net846),
    .Q(\u_reg.reg_rdata[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8913_ (.CLK(\clknet_leaf_3_u_dsync.out_clk ),
    .D(_1379_),
    .RESET_B(net858),
    .Q(\u_reg.reg_rdata[4] ));
 sky130_fd_sc_hd__dfrtp_4 _8914_ (.CLK(\clknet_leaf_15_u_dsync.out_clk ),
    .D(_1380_),
    .RESET_B(net874),
    .Q(\u_reg.reg_rdata[5] ));
 sky130_fd_sc_hd__dfrtp_4 _8915_ (.CLK(\clknet_leaf_1_u_dsync.out_clk ),
    .D(_1381_),
    .RESET_B(net848),
    .Q(\u_reg.reg_rdata[6] ));
 sky130_fd_sc_hd__dfrtp_1 _8916_ (.CLK(\clknet_leaf_5_u_dsync.out_clk ),
    .D(_1382_),
    .RESET_B(net855),
    .Q(\u_reg.reg_rdata[7] ));
 sky130_fd_sc_hd__dfrtp_2 _8917_ (.CLK(\clknet_leaf_5_u_dsync.out_clk ),
    .D(_1383_),
    .RESET_B(net856),
    .Q(\u_reg.reg_rdata[8] ));
 sky130_fd_sc_hd__dfrtp_1 _8918_ (.CLK(\clknet_leaf_6_u_dsync.out_clk ),
    .D(_1384_),
    .RESET_B(net855),
    .Q(\u_reg.reg_rdata[9] ));
 sky130_fd_sc_hd__dfrtp_4 _8919_ (.CLK(\clknet_leaf_5_u_dsync.out_clk ),
    .D(_1385_),
    .RESET_B(net860),
    .Q(\u_reg.reg_rdata[10] ));
 sky130_fd_sc_hd__dfrtp_1 _8920_ (.CLK(\clknet_leaf_7_u_dsync.out_clk ),
    .D(_1386_),
    .RESET_B(net859),
    .Q(\u_reg.reg_rdata[11] ));
 sky130_fd_sc_hd__dfrtp_4 _8921_ (.CLK(\clknet_leaf_19_u_dsync.out_clk ),
    .D(_1387_),
    .RESET_B(net883),
    .Q(\u_reg.reg_rdata[12] ));
 sky130_fd_sc_hd__dfrtp_2 _8922_ (.CLK(\clknet_leaf_12_u_dsync.out_clk ),
    .D(_1388_),
    .RESET_B(net890),
    .Q(\u_reg.reg_rdata[13] ));
 sky130_fd_sc_hd__dfrtp_2 _8923_ (.CLK(\clknet_leaf_20_u_dsync.out_clk ),
    .D(_1389_),
    .RESET_B(net896),
    .Q(\u_reg.reg_rdata[14] ));
 sky130_fd_sc_hd__dfrtp_2 _8924_ (.CLK(\clknet_leaf_35_u_dsync.out_clk ),
    .D(_1390_),
    .RESET_B(net890),
    .Q(\u_reg.reg_rdata[15] ));
 sky130_fd_sc_hd__dfrtp_4 _8925_ (.CLK(\clknet_leaf_27_u_dsync.out_clk ),
    .D(_1391_),
    .RESET_B(net894),
    .Q(\u_reg.reg_rdata[16] ));
 sky130_fd_sc_hd__dfrtp_4 _8926_ (.CLK(\clknet_leaf_27_u_dsync.out_clk ),
    .D(_1392_),
    .RESET_B(net896),
    .Q(\u_reg.reg_rdata[17] ));
 sky130_fd_sc_hd__dfrtp_4 _8927_ (.CLK(\clknet_leaf_1_u_dsync.out_clk ),
    .D(_1393_),
    .RESET_B(net846),
    .Q(\u_reg.reg_rdata[18] ));
 sky130_fd_sc_hd__dfrtp_4 _8928_ (.CLK(\clknet_leaf_2_u_dsync.out_clk ),
    .D(_1394_),
    .RESET_B(net846),
    .Q(\u_reg.reg_rdata[19] ));
 sky130_fd_sc_hd__dfrtp_4 _8929_ (.CLK(\clknet_leaf_20_u_dsync.out_clk ),
    .D(_1395_),
    .RESET_B(net894),
    .Q(\u_reg.reg_rdata[20] ));
 sky130_fd_sc_hd__dfrtp_2 _8930_ (.CLK(\clknet_leaf_19_u_dsync.out_clk ),
    .D(_1396_),
    .RESET_B(net886),
    .Q(\u_reg.reg_rdata[21] ));
 sky130_fd_sc_hd__dfrtp_1 _8931_ (.CLK(\clknet_leaf_1_u_dsync.out_clk ),
    .D(_1397_),
    .RESET_B(net847),
    .Q(\u_reg.reg_rdata[22] ));
 sky130_fd_sc_hd__dfrtp_4 _8932_ (.CLK(\clknet_leaf_0_u_dsync.out_clk ),
    .D(_1398_),
    .RESET_B(net840),
    .Q(\u_reg.reg_rdata[23] ));
 sky130_fd_sc_hd__dfrtp_1 _8933_ (.CLK(\clknet_leaf_15_u_dsync.out_clk ),
    .D(_1399_),
    .RESET_B(net870),
    .Q(\u_reg.reg_rdata[24] ));
 sky130_fd_sc_hd__dfrtp_2 _8934_ (.CLK(\clknet_leaf_16_u_dsync.out_clk ),
    .D(_1400_),
    .RESET_B(net868),
    .Q(\u_reg.reg_rdata[25] ));
 sky130_fd_sc_hd__dfrtp_4 _8935_ (.CLK(\clknet_leaf_21_u_dsync.out_clk ),
    .D(_1401_),
    .RESET_B(net894),
    .Q(\u_reg.reg_rdata[26] ));
 sky130_fd_sc_hd__dfrtp_4 _8936_ (.CLK(\clknet_leaf_15_u_dsync.out_clk ),
    .D(_1402_),
    .RESET_B(net870),
    .Q(\u_reg.reg_rdata[27] ));
 sky130_fd_sc_hd__dfrtp_4 _8937_ (.CLK(\clknet_leaf_15_u_dsync.out_clk ),
    .D(_1403_),
    .RESET_B(net870),
    .Q(\u_reg.reg_rdata[28] ));
 sky130_fd_sc_hd__dfrtp_1 _8938_ (.CLK(\clknet_leaf_17_u_dsync.out_clk ),
    .D(_1404_),
    .RESET_B(net881),
    .Q(\u_reg.reg_rdata[29] ));
 sky130_fd_sc_hd__dfrtp_4 _8939_ (.CLK(\clknet_leaf_16_u_dsync.out_clk ),
    .D(_1405_),
    .RESET_B(net874),
    .Q(\u_reg.reg_rdata[30] ));
 sky130_fd_sc_hd__dfrtp_2 _8940_ (.CLK(\clknet_leaf_17_u_dsync.out_clk ),
    .D(_1406_),
    .RESET_B(net881),
    .Q(\u_reg.reg_rdata[31] ));
 sky130_fd_sc_hd__dfrtp_4 _8941_ (.CLK(\clknet_leaf_5_u_dsync.out_clk ),
    .D(_1407_),
    .RESET_B(net848),
    .Q(\u_dcg_s0.cfg_mode[0] ));
 sky130_fd_sc_hd__dfrtp_2 _8942_ (.CLK(\clknet_leaf_5_u_dsync.out_clk ),
    .D(_1408_),
    .RESET_B(net856),
    .Q(\u_dcg_s0.cfg_mode[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8943_ (.CLK(\clknet_leaf_5_u_dsync.out_clk ),
    .D(_1409_),
    .RESET_B(net849),
    .Q(\u_dcg_s1.cfg_mode[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8944_ (.CLK(\clknet_leaf_5_u_dsync.out_clk ),
    .D(_1410_),
    .RESET_B(net854),
    .Q(\u_dcg_s1.cfg_mode[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8945_ (.CLK(\clknet_leaf_3_u_dsync.out_clk ),
    .D(_1411_),
    .RESET_B(net860),
    .Q(\u_dcg_s2.cfg_mode[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8946_ (.CLK(\clknet_leaf_15_u_dsync.out_clk ),
    .D(_1412_),
    .RESET_B(net870),
    .Q(\u_dcg_s2.cfg_mode[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8947_ (.CLK(\clknet_leaf_3_u_dsync.out_clk ),
    .D(_1413_),
    .RESET_B(net860),
    .Q(\u_dcg_peri.cfg_mode[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8948_ (.CLK(\clknet_leaf_5_u_dsync.out_clk ),
    .D(_1414_),
    .RESET_B(net855),
    .Q(\u_dcg_peri.cfg_mode[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8949_ (.CLK(\clknet_leaf_1_u_dsync.out_clk ),
    .D(_1415_),
    .RESET_B(net848),
    .Q(\u_reg.reg_2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8950_ (.CLK(\clknet_leaf_1_u_dsync.out_clk ),
    .D(_1416_),
    .RESET_B(net847),
    .Q(\u_reg.reg_2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8951_ (.CLK(\clknet_leaf_1_u_dsync.out_clk ),
    .D(_1417_),
    .RESET_B(net848),
    .Q(\u_reg.reg_2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8952_ (.CLK(\clknet_leaf_1_u_dsync.out_clk ),
    .D(_1418_),
    .RESET_B(net847),
    .Q(\u_reg.reg_2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8953_ (.CLK(\clknet_leaf_17_u_dsync.out_clk ),
    .D(_1419_),
    .RESET_B(net881),
    .Q(\u_reg.reg_2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8954_ (.CLK(\clknet_leaf_15_u_dsync.out_clk ),
    .D(_1420_),
    .RESET_B(net874),
    .Q(\u_reg.reg_2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _8955_ (.CLK(\clknet_leaf_15_u_dsync.out_clk ),
    .D(_1421_),
    .RESET_B(net868),
    .Q(\u_reg.reg_2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _8956_ (.CLK(\clknet_leaf_15_u_dsync.out_clk ),
    .D(_1422_),
    .RESET_B(net874),
    .Q(\u_reg.reg_2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _8957_ (.CLK(\clknet_leaf_22_u_dsync.out_clk ),
    .D(_1423_),
    .RESET_B(net906),
    .Q(\u_reg.reg_3[16] ));
 sky130_fd_sc_hd__dfrtp_1 _8958_ (.CLK(\clknet_leaf_24_u_dsync.out_clk ),
    .D(_1424_),
    .RESET_B(net910),
    .Q(\u_reg.reg_3[17] ));
 sky130_fd_sc_hd__dfrtp_1 _8959_ (.CLK(\clknet_leaf_16_u_dsync.out_clk ),
    .D(_1425_),
    .RESET_B(net874),
    .Q(\u_reg.reg_3[18] ));
 sky130_fd_sc_hd__dfrtp_1 _8960_ (.CLK(\clknet_leaf_16_u_dsync.out_clk ),
    .D(_1426_),
    .RESET_B(net868),
    .Q(\u_reg.reg_3[19] ));
 sky130_fd_sc_hd__dfrtp_1 _8961_ (.CLK(\clknet_leaf_21_u_dsync.out_clk ),
    .D(_1427_),
    .RESET_B(net894),
    .Q(\u_reg.reg_3[20] ));
 sky130_fd_sc_hd__dfrtp_1 _8962_ (.CLK(\clknet_leaf_18_u_dsync.out_clk ),
    .D(_1428_),
    .RESET_B(net886),
    .Q(\u_reg.reg_3[21] ));
 sky130_fd_sc_hd__dfrtp_1 _8963_ (.CLK(\clknet_leaf_3_u_dsync.out_clk ),
    .D(_1429_),
    .RESET_B(net860),
    .Q(\u_reg.reg_3[22] ));
 sky130_fd_sc_hd__dfrtp_1 _8964_ (.CLK(\clknet_leaf_16_u_dsync.out_clk ),
    .D(_1430_),
    .RESET_B(net876),
    .Q(\u_reg.reg_3[23] ));
 sky130_fd_sc_hd__dfrtp_1 _8965_ (.CLK(\clknet_leaf_23_u_dsync.out_clk ),
    .D(_1431_),
    .RESET_B(net911),
    .Q(\u_reg.reg_4[24] ));
 sky130_fd_sc_hd__dfrtp_1 _8966_ (.CLK(\clknet_leaf_23_u_dsync.out_clk ),
    .D(_1432_),
    .RESET_B(net907),
    .Q(\u_reg.reg_4[25] ));
 sky130_fd_sc_hd__dfrtp_1 _8967_ (.CLK(\clknet_leaf_22_u_dsync.out_clk ),
    .D(_1433_),
    .RESET_B(net900),
    .Q(\u_reg.reg_4[26] ));
 sky130_fd_sc_hd__dfrtp_1 _8968_ (.CLK(\clknet_leaf_25_u_dsync.out_clk ),
    .D(_1434_),
    .RESET_B(net912),
    .Q(\u_reg.reg_4[27] ));
 sky130_fd_sc_hd__dfrtp_1 _8969_ (.CLK(\clknet_leaf_21_u_dsync.out_clk ),
    .D(_1435_),
    .RESET_B(net894),
    .Q(\u_reg.reg_4[28] ));
 sky130_fd_sc_hd__dfrtp_1 _8970_ (.CLK(\clknet_leaf_21_u_dsync.out_clk ),
    .D(_1436_),
    .RESET_B(net898),
    .Q(\u_reg.reg_4[29] ));
 sky130_fd_sc_hd__dfrtp_1 _8971_ (.CLK(\clknet_leaf_23_u_dsync.out_clk ),
    .D(_1437_),
    .RESET_B(net911),
    .Q(\u_reg.reg_4[30] ));
 sky130_fd_sc_hd__dfrtp_1 _8972_ (.CLK(\clknet_leaf_18_u_dsync.out_clk ),
    .D(_1438_),
    .RESET_B(net888),
    .Q(\u_reg.reg_4[31] ));
 sky130_fd_sc_hd__dfrtp_1 _8973_ (.CLK(\clknet_leaf_22_u_dsync.out_clk ),
    .D(_1439_),
    .RESET_B(net906),
    .Q(\u_reg.reg_5[24] ));
 sky130_fd_sc_hd__dfrtp_1 _8974_ (.CLK(\clknet_leaf_22_u_dsync.out_clk ),
    .D(_1440_),
    .RESET_B(net898),
    .Q(\u_reg.reg_5[25] ));
 sky130_fd_sc_hd__dfrtp_1 _8975_ (.CLK(\clknet_leaf_21_u_dsync.out_clk ),
    .D(_1441_),
    .RESET_B(net895),
    .Q(\u_reg.reg_5[26] ));
 sky130_fd_sc_hd__dfrtp_1 _8976_ (.CLK(\clknet_leaf_21_u_dsync.out_clk ),
    .D(_1442_),
    .RESET_B(net898),
    .Q(\u_reg.reg_5[27] ));
 sky130_fd_sc_hd__dfrtp_1 _8977_ (.CLK(\clknet_leaf_17_u_dsync.out_clk ),
    .D(_1443_),
    .RESET_B(net883),
    .Q(\u_reg.reg_5[28] ));
 sky130_fd_sc_hd__dfrtp_1 _8978_ (.CLK(\clknet_leaf_21_u_dsync.out_clk ),
    .D(_1444_),
    .RESET_B(net895),
    .Q(\u_reg.reg_5[29] ));
 sky130_fd_sc_hd__dfrtp_1 _8979_ (.CLK(\clknet_leaf_21_u_dsync.out_clk ),
    .D(_1445_),
    .RESET_B(net898),
    .Q(\u_reg.reg_5[30] ));
 sky130_fd_sc_hd__dfrtp_1 _8980_ (.CLK(\clknet_leaf_16_u_dsync.out_clk ),
    .D(_1446_),
    .RESET_B(net876),
    .Q(\u_reg.reg_5[31] ));
 sky130_fd_sc_hd__dfrtp_1 _8981_ (.CLK(\clknet_leaf_22_u_dsync.out_clk ),
    .D(_1447_),
    .RESET_B(net907),
    .Q(\u_reg.reg_6[24] ));
 sky130_fd_sc_hd__dfrtp_1 _8982_ (.CLK(\clknet_leaf_22_u_dsync.out_clk ),
    .D(_1448_),
    .RESET_B(net900),
    .Q(\u_reg.reg_6[25] ));
 sky130_fd_sc_hd__dfrtp_1 _8983_ (.CLK(\clknet_leaf_18_u_dsync.out_clk ),
    .D(_1449_),
    .RESET_B(net886),
    .Q(\u_reg.reg_6[26] ));
 sky130_fd_sc_hd__dfrtp_1 _8984_ (.CLK(\clknet_leaf_26_u_dsync.out_clk ),
    .D(_1450_),
    .RESET_B(net906),
    .Q(\u_reg.reg_6[27] ));
 sky130_fd_sc_hd__dfrtp_1 _8985_ (.CLK(\clknet_leaf_17_u_dsync.out_clk ),
    .D(_1451_),
    .RESET_B(net886),
    .Q(\u_reg.reg_6[28] ));
 sky130_fd_sc_hd__dfrtp_1 _8986_ (.CLK(\clknet_leaf_21_u_dsync.out_clk ),
    .D(_1452_),
    .RESET_B(net900),
    .Q(\u_reg.reg_6[29] ));
 sky130_fd_sc_hd__dfrtp_1 _8987_ (.CLK(\clknet_leaf_22_u_dsync.out_clk ),
    .D(_1453_),
    .RESET_B(net907),
    .Q(\u_reg.reg_6[30] ));
 sky130_fd_sc_hd__dfrtp_1 _8988_ (.CLK(\clknet_leaf_16_u_dsync.out_clk ),
    .D(_1454_),
    .RESET_B(net876),
    .Q(\u_reg.reg_6[31] ));
 sky130_fd_sc_hd__dfrtp_4 _8989_ (.CLK(\clknet_leaf_1_u_dsync.out_clk ),
    .D(net575),
    .RESET_B(net846),
    .Q(\u_reg.reg_ack ));
 sky130_fd_sc_hd__dfstp_1 _8990_ (.CLK(net1773),
    .D(_1455_),
    .SET_B(net892),
    .Q(\u_dcg_s0.hcnt[0] ));
 sky130_fd_sc_hd__dfstp_1 _8991_ (.CLK(net1773),
    .D(_1456_),
    .SET_B(net892),
    .Q(\u_dcg_s0.hcnt[1] ));
 sky130_fd_sc_hd__dfstp_1 _8992_ (.CLK(net1773),
    .D(_1457_),
    .SET_B(net892),
    .Q(\u_dcg_s0.hcnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8993_ (.CLK(net1773),
    .D(_1458_),
    .RESET_B(net902),
    .Q(\u_dcg_s0.hcnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8994_ (.CLK(\clknet_leaf_7_u_dsync.out_clk ),
    .D(_1459_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8995_ (.CLK(\clknet_leaf_6_u_dsync.out_clk ),
    .D(_1460_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8996_ (.CLK(\clknet_leaf_10_u_dsync.out_clk ),
    .D(_1461_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8997_ (.CLK(\clknet_leaf_7_u_dsync.out_clk ),
    .D(_1462_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8998_ (.CLK(\clknet_leaf_9_u_dsync.out_clk ),
    .D(_1463_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8999_ (.CLK(\clknet_leaf_10_u_dsync.out_clk ),
    .D(_1464_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _9000_ (.CLK(\clknet_leaf_6_u_dsync.out_clk ),
    .D(_1465_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _9001_ (.CLK(\clknet_leaf_10_u_dsync.out_clk ),
    .D(_1466_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _9002_ (.CLK(\clknet_leaf_99_u_dsync.out_clk ),
    .D(_1467_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _9003_ (.CLK(\clknet_leaf_37_u_dsync.out_clk ),
    .D(_1468_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _9004_ (.CLK(\clknet_leaf_9_u_dsync.out_clk ),
    .D(_1469_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _9005_ (.CLK(\clknet_leaf_9_u_dsync.out_clk ),
    .D(_1470_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _9006_ (.CLK(\clknet_leaf_37_u_dsync.out_clk ),
    .D(_1471_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _9007_ (.CLK(\clknet_leaf_63_u_dsync.out_clk ),
    .D(_1472_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _9008_ (.CLK(\clknet_leaf_64_u_dsync.out_clk ),
    .D(_1473_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _9009_ (.CLK(\clknet_leaf_64_u_dsync.out_clk ),
    .D(_1474_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _9010_ (.CLK(\clknet_leaf_65_u_dsync.out_clk ),
    .D(_1475_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _9011_ (.CLK(\clknet_leaf_65_u_dsync.out_clk ),
    .D(_1476_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _9012_ (.CLK(\clknet_leaf_64_u_dsync.out_clk ),
    .D(_1477_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _9013_ (.CLK(\clknet_leaf_68_u_dsync.out_clk ),
    .D(_1478_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _9014_ (.CLK(\clknet_leaf_39_u_dsync.out_clk ),
    .D(_1479_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _9015_ (.CLK(\clknet_leaf_65_u_dsync.out_clk ),
    .D(_1480_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _9016_ (.CLK(\clknet_leaf_64_u_dsync.out_clk ),
    .D(_1481_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _9017_ (.CLK(\clknet_leaf_41_u_dsync.out_clk ),
    .D(_1482_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _9018_ (.CLK(\clknet_leaf_39_u_dsync.out_clk ),
    .D(_1483_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _9019_ (.CLK(\clknet_leaf_39_u_dsync.out_clk ),
    .D(_1484_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _9020_ (.CLK(\clknet_leaf_67_u_dsync.out_clk ),
    .D(_1485_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _9021_ (.CLK(\clknet_leaf_38_u_dsync.out_clk ),
    .D(_1486_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _9022_ (.CLK(\clknet_leaf_68_u_dsync.out_clk ),
    .D(_1487_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _9023_ (.CLK(\clknet_leaf_39_u_dsync.out_clk ),
    .D(_1488_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _9024_ (.CLK(\clknet_leaf_38_u_dsync.out_clk ),
    .D(_1489_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _9025_ (.CLK(\clknet_leaf_68_u_dsync.out_clk ),
    .D(_1490_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _9026_ (.CLK(\clknet_leaf_38_u_dsync.out_clk ),
    .D(_1491_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _9027_ (.CLK(\clknet_leaf_65_u_dsync.out_clk ),
    .D(_1492_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _9028_ (.CLK(\clknet_leaf_69_u_dsync.out_clk ),
    .D(_1493_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _9029_ (.CLK(\clknet_leaf_66_u_dsync.out_clk ),
    .D(_1494_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _9030_ (.CLK(\clknet_leaf_66_u_dsync.out_clk ),
    .D(_1495_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _9031_ (.CLK(\clknet_leaf_38_u_dsync.out_clk ),
    .D(_1496_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _9032_ (.CLK(\clknet_leaf_67_u_dsync.out_clk ),
    .D(_1497_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _9033_ (.CLK(\clknet_leaf_95_u_dsync.out_clk ),
    .D(_1498_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _9034_ (.CLK(\clknet_leaf_38_u_dsync.out_clk ),
    .D(_1499_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _9035_ (.CLK(\clknet_leaf_37_u_dsync.out_clk ),
    .D(_1500_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _9036_ (.CLK(\clknet_leaf_68_u_dsync.out_clk ),
    .D(_1501_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][47] ));
 sky130_fd_sc_hd__dfxtp_1 _9037_ (.CLK(\clknet_leaf_95_u_dsync.out_clk ),
    .D(_1502_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][48] ));
 sky130_fd_sc_hd__dfxtp_1 _9038_ (.CLK(\clknet_leaf_67_u_dsync.out_clk ),
    .D(_1503_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][49] ));
 sky130_fd_sc_hd__dfxtp_1 _9039_ (.CLK(\clknet_leaf_38_u_dsync.out_clk ),
    .D(_1504_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][50] ));
 sky130_fd_sc_hd__dfxtp_1 _9040_ (.CLK(\clknet_leaf_8_u_dsync.out_clk ),
    .D(_1505_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][53] ));
 sky130_fd_sc_hd__dfxtp_1 _9041_ (.CLK(\clknet_leaf_96_u_dsync.out_clk ),
    .D(_1506_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][54] ));
 sky130_fd_sc_hd__dfxtp_1 _9042_ (.CLK(\clknet_leaf_7_u_dsync.out_clk ),
    .D(_1507_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][55] ));
 sky130_fd_sc_hd__dfxtp_1 _9043_ (.CLK(\clknet_leaf_7_u_dsync.out_clk ),
    .D(_1508_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][56] ));
 sky130_fd_sc_hd__dfxtp_1 _9044_ (.CLK(\clknet_leaf_96_u_dsync.out_clk ),
    .D(_1509_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][57] ));
 sky130_fd_sc_hd__dfxtp_1 _9045_ (.CLK(\clknet_leaf_8_u_dsync.out_clk ),
    .D(_1510_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][58] ));
 sky130_fd_sc_hd__dfxtp_1 _9046_ (.CLK(\clknet_leaf_8_u_dsync.out_clk ),
    .D(_1511_),
    .Q(\u_s1.u_sync_wbb.u_cmd_if.mem[0][59] ));
 sky130_fd_sc_hd__dfrtp_1 _9047_ (.CLK(net1766),
    .D(\u_dcg_s2.cfg_mode[0] ),
    .RESET_B(net869),
    .Q(\u_dcg_s2.u_dsync.in_data_s[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9048_ (.CLK(net1770),
    .D(\u_dcg_s2.cfg_mode[1] ),
    .RESET_B(net875),
    .Q(\u_dcg_s2.u_dsync.in_data_s[1] ));
 sky130_fd_sc_hd__dfrtp_1 _9049_ (.CLK(net1766),
    .D(\u_dcg_s2.u_dsync.in_data_s[0] ),
    .RESET_B(net869),
    .Q(\u_dcg_s2.u_dsync.in_data_2s[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9050_ (.CLK(net1770),
    .D(\u_dcg_s2.u_dsync.in_data_s[1] ),
    .RESET_B(net875),
    .Q(\u_dcg_s2.u_dsync.in_data_2s[1] ));
 sky130_fd_sc_hd__dfrtp_1 _9051_ (.CLK(net1770),
    .D(\u_dcg_s2.u_dsync.in_data_2s[0] ),
    .RESET_B(net871),
    .Q(\u_dcg_s2.cfg_mode_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9052_ (.CLK(net1770),
    .D(\u_dcg_s2.u_dsync.in_data_2s[1] ),
    .RESET_B(net870),
    .Q(\u_dcg_s2.cfg_mode_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _9053_ (.CLK(net1766),
    .D(\u_dcg_s1.cfg_mode[0] ),
    .RESET_B(net855),
    .Q(\u_dcg_s1.u_dsync.in_data_s[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9054_ (.CLK(clknet_2_1__leaf_mclk_raw),
    .D(\u_dcg_s1.cfg_mode[1] ),
    .RESET_B(net848),
    .Q(\u_dcg_s1.u_dsync.in_data_s[1] ));
 sky130_fd_sc_hd__dfrtp_1 _9055_ (.CLK(net1767),
    .D(\u_dcg_s1.u_dsync.in_data_s[0] ),
    .RESET_B(net854),
    .Q(\u_dcg_s1.u_dsync.in_data_2s[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9056_ (.CLK(clknet_2_1__leaf_mclk_raw),
    .D(net1961),
    .RESET_B(net848),
    .Q(\u_dcg_s1.u_dsync.in_data_2s[1] ));
 sky130_fd_sc_hd__dfrtp_1 _9057_ (.CLK(clknet_2_1__leaf_mclk_raw),
    .D(\u_dcg_s1.u_dsync.in_data_2s[0] ),
    .RESET_B(net854),
    .Q(\u_dcg_s1.cfg_mode_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9058_ (.CLK(clknet_2_1__leaf_mclk_raw),
    .D(net1963),
    .RESET_B(net850),
    .Q(\u_dcg_s1.cfg_mode_ss[1] ));
 sky130_fd_sc_hd__dfstp_2 _9059_ (.CLK(\clknet_leaf_100_u_dsync.out_clk ),
    .D(_0000_),
    .SET_B(net840),
    .Q(\u_s0.u_sync_wbb.m_state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _9060_ (.CLK(\clknet_leaf_100_u_dsync.out_clk ),
    .D(_0001_),
    .RESET_B(net841),
    .Q(\u_s0.u_sync_wbb.m_state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _9061_ (.CLK(\clknet_leaf_98_u_dsync.out_clk ),
    .D(_0002_),
    .RESET_B(net847),
    .Q(\u_s0.u_sync_wbb.m_state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _9062_ (.CLK(\clknet_leaf_100_u_dsync.out_clk ),
    .D(_1512_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _9063_ (.CLK(\clknet_leaf_105_u_dsync.out_clk ),
    .D(_1513_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _9064_ (.CLK(\clknet_leaf_6_u_dsync.out_clk ),
    .D(_1514_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _9065_ (.CLK(\clknet_leaf_97_u_dsync.out_clk ),
    .D(_1515_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _9066_ (.CLK(\clknet_leaf_94_u_dsync.out_clk ),
    .D(_1516_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _9067_ (.CLK(\clknet_leaf_98_u_dsync.out_clk ),
    .D(_1517_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _9068_ (.CLK(\clknet_leaf_97_u_dsync.out_clk ),
    .D(_1518_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _9069_ (.CLK(\clknet_leaf_97_u_dsync.out_clk ),
    .D(_1519_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _9070_ (.CLK(\clknet_leaf_98_u_dsync.out_clk ),
    .D(_1520_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _9071_ (.CLK(\clknet_leaf_101_u_dsync.out_clk ),
    .D(_1521_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _9072_ (.CLK(\clknet_leaf_100_u_dsync.out_clk ),
    .D(_1522_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _9073_ (.CLK(\clknet_leaf_102_u_dsync.out_clk ),
    .D(_1523_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _9074_ (.CLK(\clknet_leaf_88_u_dsync.out_clk ),
    .D(_1524_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _9075_ (.CLK(\clknet_leaf_89_u_dsync.out_clk ),
    .D(_1525_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _9076_ (.CLK(\clknet_leaf_70_u_dsync.out_clk ),
    .D(_1526_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _9077_ (.CLK(\clknet_leaf_70_u_dsync.out_clk ),
    .D(_1527_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _9078_ (.CLK(\clknet_leaf_69_u_dsync.out_clk ),
    .D(_1528_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _9079_ (.CLK(\clknet_leaf_93_u_dsync.out_clk ),
    .D(_1529_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _9080_ (.CLK(\clknet_leaf_86_u_dsync.out_clk ),
    .D(_1530_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _9081_ (.CLK(\clknet_leaf_93_u_dsync.out_clk ),
    .D(_1531_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _9082_ (.CLK(\clknet_leaf_70_u_dsync.out_clk ),
    .D(_1532_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _9083_ (.CLK(\clknet_leaf_86_u_dsync.out_clk ),
    .D(_1533_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _9084_ (.CLK(\clknet_leaf_86_u_dsync.out_clk ),
    .D(_1534_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _9085_ (.CLK(\clknet_leaf_93_u_dsync.out_clk ),
    .D(_1535_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _9086_ (.CLK(\clknet_leaf_94_u_dsync.out_clk ),
    .D(_1536_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _9087_ (.CLK(\clknet_leaf_69_u_dsync.out_clk ),
    .D(_1537_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _9088_ (.CLK(\clknet_leaf_88_u_dsync.out_clk ),
    .D(_1538_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _9089_ (.CLK(\clknet_leaf_87_u_dsync.out_clk ),
    .D(_1539_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _9090_ (.CLK(\clknet_leaf_95_u_dsync.out_clk ),
    .D(_1540_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _9091_ (.CLK(\clknet_leaf_92_u_dsync.out_clk ),
    .D(_1541_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _9092_ (.CLK(\clknet_leaf_87_u_dsync.out_clk ),
    .D(_1542_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _9093_ (.CLK(\clknet_leaf_94_u_dsync.out_clk ),
    .D(_1543_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _9094_ (.CLK(\clknet_leaf_89_u_dsync.out_clk ),
    .D(_1544_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _9095_ (.CLK(\clknet_leaf_92_u_dsync.out_clk ),
    .D(_1545_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _9096_ (.CLK(\clknet_leaf_87_u_dsync.out_clk ),
    .D(_1546_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _9097_ (.CLK(\clknet_leaf_92_u_dsync.out_clk ),
    .D(_1547_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _9098_ (.CLK(\clknet_leaf_87_u_dsync.out_clk ),
    .D(_1548_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _9099_ (.CLK(\clknet_leaf_94_u_dsync.out_clk ),
    .D(_1549_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _9100_ (.CLK(\clknet_leaf_92_u_dsync.out_clk ),
    .D(_1550_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _9101_ (.CLK(\clknet_leaf_91_u_dsync.out_clk ),
    .D(_1551_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _9102_ (.CLK(\clknet_leaf_90_u_dsync.out_clk ),
    .D(_1552_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _9103_ (.CLK(\clknet_leaf_101_u_dsync.out_clk ),
    .D(_1553_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _9104_ (.CLK(\clknet_leaf_89_u_dsync.out_clk ),
    .D(_1554_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _9105_ (.CLK(\clknet_leaf_86_u_dsync.out_clk ),
    .D(_1555_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][47] ));
 sky130_fd_sc_hd__dfxtp_1 _9106_ (.CLK(\clknet_leaf_91_u_dsync.out_clk ),
    .D(_1556_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][48] ));
 sky130_fd_sc_hd__dfxtp_1 _9107_ (.CLK(\clknet_leaf_90_u_dsync.out_clk ),
    .D(_1557_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][49] ));
 sky130_fd_sc_hd__dfxtp_1 _9108_ (.CLK(\clknet_leaf_101_u_dsync.out_clk ),
    .D(_1558_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][50] ));
 sky130_fd_sc_hd__dfxtp_1 _9109_ (.CLK(\clknet_leaf_106_u_dsync.out_clk ),
    .D(_1559_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][53] ));
 sky130_fd_sc_hd__dfxtp_1 _9110_ (.CLK(\clknet_leaf_106_u_dsync.out_clk ),
    .D(_1560_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][54] ));
 sky130_fd_sc_hd__dfxtp_1 _9111_ (.CLK(\clknet_leaf_101_u_dsync.out_clk ),
    .D(_1561_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][55] ));
 sky130_fd_sc_hd__dfxtp_1 _9112_ (.CLK(\clknet_leaf_100_u_dsync.out_clk ),
    .D(_1562_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][56] ));
 sky130_fd_sc_hd__dfxtp_1 _9113_ (.CLK(\clknet_leaf_103_u_dsync.out_clk ),
    .D(_1563_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][57] ));
 sky130_fd_sc_hd__dfxtp_1 _9114_ (.CLK(\clknet_leaf_88_u_dsync.out_clk ),
    .D(_1564_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][58] ));
 sky130_fd_sc_hd__dfxtp_1 _9115_ (.CLK(\clknet_leaf_101_u_dsync.out_clk ),
    .D(_1565_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][59] ));
 sky130_fd_sc_hd__dfxtp_1 _9116_ (.CLK(\clknet_leaf_105_u_dsync.out_clk ),
    .D(_1566_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][60] ));
 sky130_fd_sc_hd__dfxtp_1 _9117_ (.CLK(\clknet_leaf_106_u_dsync.out_clk ),
    .D(_1567_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][61] ));
 sky130_fd_sc_hd__dfxtp_1 _9118_ (.CLK(\clknet_leaf_107_u_dsync.out_clk ),
    .D(_1568_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][62] ));
 sky130_fd_sc_hd__dfxtp_1 _9119_ (.CLK(\clknet_leaf_107_u_dsync.out_clk ),
    .D(_1569_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][63] ));
 sky130_fd_sc_hd__dfxtp_1 _9120_ (.CLK(\clknet_leaf_107_u_dsync.out_clk ),
    .D(_1570_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][64] ));
 sky130_fd_sc_hd__dfxtp_1 _9121_ (.CLK(\clknet_leaf_108_u_dsync.out_clk ),
    .D(_1571_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][65] ));
 sky130_fd_sc_hd__dfxtp_1 _9122_ (.CLK(\clknet_leaf_108_u_dsync.out_clk ),
    .D(_1572_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][66] ));
 sky130_fd_sc_hd__dfxtp_1 _9123_ (.CLK(\clknet_leaf_102_u_dsync.out_clk ),
    .D(_1573_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][67] ));
 sky130_fd_sc_hd__dfxtp_1 _9124_ (.CLK(\clknet_leaf_102_u_dsync.out_clk ),
    .D(_1574_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][68] ));
 sky130_fd_sc_hd__dfxtp_1 _9125_ (.CLK(\clknet_leaf_103_u_dsync.out_clk ),
    .D(_1575_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][69] ));
 sky130_fd_sc_hd__dfxtp_1 _9126_ (.CLK(\clknet_leaf_90_u_dsync.out_clk ),
    .D(_1576_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][70] ));
 sky130_fd_sc_hd__dfxtp_1 _9127_ (.CLK(\clknet_leaf_106_u_dsync.out_clk ),
    .D(_1577_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][71] ));
 sky130_fd_sc_hd__dfxtp_1 _9128_ (.CLK(\clknet_leaf_103_u_dsync.out_clk ),
    .D(_1578_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][72] ));
 sky130_fd_sc_hd__dfxtp_1 _9129_ (.CLK(\clknet_leaf_102_u_dsync.out_clk ),
    .D(_1579_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][73] ));
 sky130_fd_sc_hd__dfxtp_1 _9130_ (.CLK(\clknet_leaf_103_u_dsync.out_clk ),
    .D(_1580_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][74] ));
 sky130_fd_sc_hd__dfxtp_1 _9131_ (.CLK(\clknet_leaf_104_u_dsync.out_clk ),
    .D(_1581_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][75] ));
 sky130_fd_sc_hd__dfxtp_1 _9132_ (.CLK(\clknet_leaf_104_u_dsync.out_clk ),
    .D(_1582_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][76] ));
 sky130_fd_sc_hd__dfxtp_1 _9133_ (.CLK(\clknet_leaf_103_u_dsync.out_clk ),
    .D(_1583_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][77] ));
 sky130_fd_sc_hd__dfxtp_1 _9134_ (.CLK(\clknet_leaf_104_u_dsync.out_clk ),
    .D(_1584_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][78] ));
 sky130_fd_sc_hd__dfxtp_1 _9135_ (.CLK(\clknet_leaf_102_u_dsync.out_clk ),
    .D(_1585_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][79] ));
 sky130_fd_sc_hd__dfxtp_1 _9136_ (.CLK(\clknet_leaf_105_u_dsync.out_clk ),
    .D(_1586_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][80] ));
 sky130_fd_sc_hd__dfxtp_1 _9137_ (.CLK(\clknet_leaf_105_u_dsync.out_clk ),
    .D(_1587_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][81] ));
 sky130_fd_sc_hd__dfxtp_1 _9138_ (.CLK(\clknet_leaf_103_u_dsync.out_clk ),
    .D(_1588_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[1][82] ));
 sky130_fd_sc_hd__dfxtp_1 _9139_ (.CLK(\clknet_leaf_100_u_dsync.out_clk ),
    .D(_1589_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _9140_ (.CLK(\clknet_leaf_105_u_dsync.out_clk ),
    .D(_1590_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _9141_ (.CLK(\clknet_leaf_99_u_dsync.out_clk ),
    .D(_1591_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _9142_ (.CLK(\clknet_leaf_97_u_dsync.out_clk ),
    .D(_1592_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _9143_ (.CLK(\clknet_leaf_98_u_dsync.out_clk ),
    .D(_1593_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _9144_ (.CLK(\clknet_leaf_98_u_dsync.out_clk ),
    .D(_1594_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _9145_ (.CLK(\clknet_leaf_98_u_dsync.out_clk ),
    .D(_1595_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _9146_ (.CLK(\clknet_leaf_97_u_dsync.out_clk ),
    .D(_1596_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _9147_ (.CLK(\clknet_leaf_99_u_dsync.out_clk ),
    .D(_1597_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _9148_ (.CLK(\clknet_leaf_101_u_dsync.out_clk ),
    .D(_1598_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _9149_ (.CLK(\clknet_leaf_106_u_dsync.out_clk ),
    .D(_1599_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _9150_ (.CLK(\clknet_leaf_102_u_dsync.out_clk ),
    .D(_1600_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _9151_ (.CLK(\clknet_leaf_88_u_dsync.out_clk ),
    .D(_1601_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _9152_ (.CLK(\clknet_leaf_90_u_dsync.out_clk ),
    .D(_1602_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _9153_ (.CLK(\clknet_leaf_70_u_dsync.out_clk ),
    .D(_1603_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _9154_ (.CLK(\clknet_leaf_70_u_dsync.out_clk ),
    .D(_1604_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _9155_ (.CLK(\clknet_leaf_69_u_dsync.out_clk ),
    .D(_1605_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _9156_ (.CLK(\clknet_leaf_93_u_dsync.out_clk ),
    .D(_1606_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _9157_ (.CLK(\clknet_leaf_92_u_dsync.out_clk ),
    .D(_1607_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _9158_ (.CLK(\clknet_leaf_93_u_dsync.out_clk ),
    .D(_1608_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _9159_ (.CLK(\clknet_leaf_93_u_dsync.out_clk ),
    .D(_1609_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _9160_ (.CLK(\clknet_leaf_86_u_dsync.out_clk ),
    .D(_1610_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _9161_ (.CLK(\clknet_leaf_93_u_dsync.out_clk ),
    .D(_1611_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _9162_ (.CLK(\clknet_leaf_93_u_dsync.out_clk ),
    .D(_1612_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _9163_ (.CLK(\clknet_leaf_94_u_dsync.out_clk ),
    .D(_1613_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _9164_ (.CLK(\clknet_leaf_94_u_dsync.out_clk ),
    .D(_1614_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _9165_ (.CLK(\clknet_leaf_89_u_dsync.out_clk ),
    .D(_1615_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _9166_ (.CLK(\clknet_leaf_86_u_dsync.out_clk ),
    .D(_1616_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _9167_ (.CLK(\clknet_leaf_95_u_dsync.out_clk ),
    .D(_1617_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _9168_ (.CLK(\clknet_leaf_92_u_dsync.out_clk ),
    .D(_1618_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _9169_ (.CLK(\clknet_leaf_92_u_dsync.out_clk ),
    .D(_1619_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _9170_ (.CLK(\clknet_leaf_94_u_dsync.out_clk ),
    .D(_1620_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _9171_ (.CLK(\clknet_leaf_89_u_dsync.out_clk ),
    .D(_1621_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _9172_ (.CLK(\clknet_leaf_91_u_dsync.out_clk ),
    .D(_1622_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _9173_ (.CLK(\clknet_leaf_88_u_dsync.out_clk ),
    .D(_1623_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _9174_ (.CLK(\clknet_leaf_92_u_dsync.out_clk ),
    .D(_1624_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _9175_ (.CLK(\clknet_leaf_89_u_dsync.out_clk ),
    .D(_1625_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _9176_ (.CLK(\clknet_leaf_94_u_dsync.out_clk ),
    .D(_1626_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _9177_ (.CLK(\clknet_leaf_91_u_dsync.out_clk ),
    .D(_1627_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _9178_ (.CLK(\clknet_leaf_91_u_dsync.out_clk ),
    .D(_1628_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _9179_ (.CLK(\clknet_leaf_90_u_dsync.out_clk ),
    .D(_1629_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _9180_ (.CLK(\clknet_leaf_101_u_dsync.out_clk ),
    .D(_1630_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _9181_ (.CLK(\clknet_leaf_89_u_dsync.out_clk ),
    .D(_1631_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _9182_ (.CLK(\clknet_leaf_92_u_dsync.out_clk ),
    .D(_1632_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][47] ));
 sky130_fd_sc_hd__dfxtp_1 _9183_ (.CLK(\clknet_leaf_91_u_dsync.out_clk ),
    .D(_1633_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][48] ));
 sky130_fd_sc_hd__dfxtp_1 _9184_ (.CLK(\clknet_leaf_90_u_dsync.out_clk ),
    .D(_1634_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][49] ));
 sky130_fd_sc_hd__dfxtp_1 _9185_ (.CLK(\clknet_leaf_98_u_dsync.out_clk ),
    .D(_1635_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][50] ));
 sky130_fd_sc_hd__dfxtp_1 _9186_ (.CLK(\clknet_leaf_106_u_dsync.out_clk ),
    .D(_1636_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][53] ));
 sky130_fd_sc_hd__dfxtp_1 _9187_ (.CLK(\clknet_leaf_106_u_dsync.out_clk ),
    .D(_1637_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][54] ));
 sky130_fd_sc_hd__dfxtp_1 _9188_ (.CLK(\clknet_leaf_101_u_dsync.out_clk ),
    .D(_1638_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][55] ));
 sky130_fd_sc_hd__dfxtp_1 _9189_ (.CLK(\clknet_leaf_100_u_dsync.out_clk ),
    .D(_1639_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][56] ));
 sky130_fd_sc_hd__dfxtp_1 _9190_ (.CLK(\clknet_leaf_102_u_dsync.out_clk ),
    .D(_1640_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][57] ));
 sky130_fd_sc_hd__dfxtp_1 _9191_ (.CLK(\clknet_leaf_88_u_dsync.out_clk ),
    .D(_1641_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][58] ));
 sky130_fd_sc_hd__dfxtp_1 _9192_ (.CLK(\clknet_leaf_100_u_dsync.out_clk ),
    .D(_1642_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][59] ));
 sky130_fd_sc_hd__dfxtp_1 _9193_ (.CLK(\clknet_leaf_105_u_dsync.out_clk ),
    .D(_1643_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][60] ));
 sky130_fd_sc_hd__dfxtp_1 _9194_ (.CLK(\clknet_leaf_106_u_dsync.out_clk ),
    .D(_1644_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][61] ));
 sky130_fd_sc_hd__dfxtp_1 _9195_ (.CLK(\clknet_leaf_107_u_dsync.out_clk ),
    .D(_1645_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][62] ));
 sky130_fd_sc_hd__dfxtp_1 _9196_ (.CLK(\clknet_leaf_107_u_dsync.out_clk ),
    .D(_1646_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][63] ));
 sky130_fd_sc_hd__dfxtp_1 _9197_ (.CLK(\clknet_leaf_108_u_dsync.out_clk ),
    .D(_1647_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][64] ));
 sky130_fd_sc_hd__dfxtp_1 _9198_ (.CLK(\clknet_leaf_108_u_dsync.out_clk ),
    .D(_1648_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][65] ));
 sky130_fd_sc_hd__dfxtp_1 _9199_ (.CLK(\clknet_leaf_108_u_dsync.out_clk ),
    .D(_1649_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][66] ));
 sky130_fd_sc_hd__dfxtp_1 _9200_ (.CLK(\clknet_leaf_102_u_dsync.out_clk ),
    .D(_1650_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][67] ));
 sky130_fd_sc_hd__dfxtp_1 _9201_ (.CLK(\clknet_leaf_102_u_dsync.out_clk ),
    .D(_1651_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][68] ));
 sky130_fd_sc_hd__dfxtp_1 _9202_ (.CLK(\clknet_leaf_103_u_dsync.out_clk ),
    .D(_1652_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][69] ));
 sky130_fd_sc_hd__dfxtp_1 _9203_ (.CLK(\clknet_leaf_103_u_dsync.out_clk ),
    .D(_1653_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][70] ));
 sky130_fd_sc_hd__dfxtp_1 _9204_ (.CLK(\clknet_leaf_106_u_dsync.out_clk ),
    .D(_1654_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][71] ));
 sky130_fd_sc_hd__dfxtp_1 _9205_ (.CLK(\clknet_leaf_104_u_dsync.out_clk ),
    .D(_1655_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][72] ));
 sky130_fd_sc_hd__dfxtp_1 _9206_ (.CLK(\clknet_leaf_106_u_dsync.out_clk ),
    .D(_1656_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][73] ));
 sky130_fd_sc_hd__dfxtp_1 _9207_ (.CLK(\clknet_leaf_103_u_dsync.out_clk ),
    .D(_1657_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][74] ));
 sky130_fd_sc_hd__dfxtp_1 _9208_ (.CLK(\clknet_leaf_104_u_dsync.out_clk ),
    .D(_1658_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][75] ));
 sky130_fd_sc_hd__dfxtp_1 _9209_ (.CLK(\clknet_leaf_104_u_dsync.out_clk ),
    .D(_1659_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][76] ));
 sky130_fd_sc_hd__dfxtp_1 _9210_ (.CLK(\clknet_leaf_104_u_dsync.out_clk ),
    .D(_1660_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][77] ));
 sky130_fd_sc_hd__dfxtp_1 _9211_ (.CLK(\clknet_leaf_104_u_dsync.out_clk ),
    .D(_1661_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][78] ));
 sky130_fd_sc_hd__dfxtp_1 _9212_ (.CLK(\clknet_leaf_103_u_dsync.out_clk ),
    .D(_1662_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][79] ));
 sky130_fd_sc_hd__dfxtp_1 _9213_ (.CLK(\clknet_leaf_105_u_dsync.out_clk ),
    .D(_1663_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][80] ));
 sky130_fd_sc_hd__dfxtp_1 _9214_ (.CLK(\clknet_leaf_108_u_dsync.out_clk ),
    .D(_1664_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][81] ));
 sky130_fd_sc_hd__dfxtp_1 _9215_ (.CLK(\clknet_leaf_103_u_dsync.out_clk ),
    .D(_1665_),
    .Q(\u_s0.u_sync_wbb.u_cmd_if.mem[2][82] ));
 sky130_fd_sc_hd__dfrtp_1 _9216_ (.CLK(net1770),
    .D(\u_dcg_s0.cfg_mode[0] ),
    .RESET_B(net881),
    .Q(\u_dcg_s0.u_dsync.in_data_s[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9217_ (.CLK(clknet_2_2__leaf_mclk_raw),
    .D(net1279),
    .RESET_B(net890),
    .Q(\u_dcg_s0.u_dsync.in_data_s[1] ));
 sky130_fd_sc_hd__dfrtp_4 _9218_ (.CLK(clknet_2_2__leaf_mclk_raw),
    .D(\u_dcg_s0.u_dsync.in_data_s[0] ),
    .RESET_B(net885),
    .Q(\u_dcg_s0.u_dsync.in_data_2s[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9219_ (.CLK(clknet_2_2__leaf_mclk_raw),
    .D(net1971),
    .RESET_B(net890),
    .Q(\u_dcg_s0.u_dsync.in_data_2s[1] ));
 sky130_fd_sc_hd__dfrtp_2 _9220_ (.CLK(net1773),
    .D(net1922),
    .RESET_B(net902),
    .Q(\u_dcg_s0.cfg_mode_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9221_ (.CLK(net1773),
    .D(net1849),
    .RESET_B(net891),
    .Q(\u_dcg_s0.cfg_mode_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _9222_ (.CLK(clknet_2_3__leaf_mclk_raw),
    .D(net1511),
    .RESET_B(net891),
    .Q(\u_dcg_s0.dst_idle_r ));
 sky130_fd_sc_hd__dfstp_1 _9223_ (.CLK(clknet_2_3__leaf_mclk_raw),
    .D(_1666_),
    .SET_B(net891),
    .Q(\u_dcg_s0.idle_his ));
 sky130_fd_sc_hd__dfrtp_1 _9224_ (.CLK(\clknet_leaf_0_u_dsync.out_clk ),
    .D(_1667_),
    .RESET_B(net841),
    .Q(\u_wbi_arb.gnt[0] ));
 sky130_fd_sc_hd__dfrtp_2 _9225_ (.CLK(\clknet_leaf_107_u_dsync.out_clk ),
    .D(_1668_),
    .RESET_B(net841),
    .Q(\u_wbi_arb.gnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _9226_ (.CLK(net1770),
    .D(\u_dcg_riscv.cfg_mode[0] ),
    .RESET_B(net875),
    .Q(\u_dcg_riscv.u_dsync.in_data_s[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9227_ (.CLK(net1771),
    .D(\u_dcg_riscv.cfg_mode[1] ),
    .RESET_B(net908),
    .Q(\u_dcg_riscv.u_dsync.in_data_s[1] ));
 sky130_fd_sc_hd__dfrtp_1 _9228_ (.CLK(net1770),
    .D(net1977),
    .RESET_B(net875),
    .Q(\u_dcg_riscv.u_dsync.in_data_2s[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9229_ (.CLK(net1771),
    .D(\u_dcg_riscv.u_dsync.in_data_s[1] ),
    .RESET_B(net907),
    .Q(\u_dcg_riscv.u_dsync.in_data_2s[1] ));
 sky130_fd_sc_hd__dfrtp_1 _9230_ (.CLK(net1770),
    .D(\u_dcg_riscv.u_dsync.in_data_2s[0] ),
    .RESET_B(net875),
    .Q(\u_dcg_riscv.cfg_mode_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9231_ (.CLK(net1771),
    .D(\u_dcg_riscv.u_dsync.in_data_2s[1] ),
    .RESET_B(net908),
    .Q(\u_dcg_riscv.cfg_mode_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _9232_ (.CLK(net1766),
    .D(\u_dcg_peri.cfg_mode[0] ),
    .RESET_B(net859),
    .Q(\u_dcg_peri.u_dsync.in_data_s[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9233_ (.CLK(net1766),
    .D(\u_dcg_peri.cfg_mode[1] ),
    .RESET_B(net861),
    .Q(\u_dcg_peri.u_dsync.in_data_s[1] ));
 sky130_fd_sc_hd__dfrtp_1 _9234_ (.CLK(net1766),
    .D(\u_dcg_peri.u_dsync.in_data_s[0] ),
    .RESET_B(net859),
    .Q(\u_dcg_peri.u_dsync.in_data_2s[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9235_ (.CLK(net1766),
    .D(\u_dcg_peri.u_dsync.in_data_s[1] ),
    .RESET_B(net859),
    .Q(\u_dcg_peri.u_dsync.in_data_2s[1] ));
 sky130_fd_sc_hd__dfrtp_1 _9236_ (.CLK(net1766),
    .D(\u_dcg_peri.u_dsync.in_data_2s[0] ),
    .RESET_B(net859),
    .Q(\u_dcg_peri.cfg_mode_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _9237_ (.CLK(net1766),
    .D(\u_dcg_peri.u_dsync.in_data_2s[1] ),
    .RESET_B(net860),
    .Q(\u_dcg_peri.cfg_mode_ss[1] ));
 sky130_fd_sc_hd__clkbuf_1 _9254_ (.A(ch_clk_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 _9255_ (.A(net1716),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 _9256_ (.A(net1715),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 _9257_ (.A(ch_data_in[0]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 _9258_ (.A(ch_data_in[1]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 _9259_ (.A(ch_data_in[2]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 _9260_ (.A(ch_data_in[3]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 _9261_ (.A(ch_data_in[4]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 _9262_ (.A(ch_data_in[5]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 _9263_ (.A(ch_data_in[6]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 _9264_ (.A(ch_data_in[7]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_4 _9265_ (.A(ch_data_in[8]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_4 _9266_ (.A(ch_data_in[9]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_4 _9267_ (.A(ch_data_in[10]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 _9268_ (.A(ch_data_in[11]),
    .X(net26));
 sky130_fd_sc_hd__buf_2 _9269_ (.A(net1689),
    .X(net37));
 sky130_fd_sc_hd__buf_2 _9270_ (.A(net1686),
    .X(net48));
 sky130_fd_sc_hd__buf_2 _9271_ (.A(net1680),
    .X(net59));
 sky130_fd_sc_hd__buf_2 _9272_ (.A(net1663),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 _9273_ (.A(ch_data_in[16]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 _9274_ (.A(ch_data_in[17]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 _9275_ (.A(ch_data_in[18]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 _9276_ (.A(ch_data_in[19]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 _9277_ (.A(ch_data_in[20]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 _9278_ (.A(ch_data_in[21]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _9279_ (.A(ch_data_in[22]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _9280_ (.A(ch_data_in[23]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 _9281_ (.A(net1662),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 _9282_ (.A(net1661),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _9283_ (.A(net1660),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _9284_ (.A(net1659),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 _9285_ (.A(net1658),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 _9286_ (.A(net1657),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 _9287_ (.A(net1656),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 _9288_ (.A(net1655),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 _9289_ (.A(net1654),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 _9290_ (.A(net1653),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 _9291_ (.A(net1652),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 _9292_ (.A(net1651),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 _9293_ (.A(net1650),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 _9294_ (.A(net1649),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 _9295_ (.A(net1648),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 _9296_ (.A(net1647),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 _9297_ (.A(net1646),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 _9298_ (.A(net1645),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 _9299_ (.A(net1644),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 _9300_ (.A(net1643),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_2 _9301_ (.A(ch_data_in[44]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 _9302_ (.A(ch_data_in[45]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 _9303_ (.A(ch_data_in[46]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 _9304_ (.A(ch_data_in[47]),
    .X(net103));
 sky130_fd_sc_hd__buf_2 _9305_ (.A(ch_data_in[48]),
    .X(net104));
 sky130_fd_sc_hd__buf_2 _9306_ (.A(ch_data_in[49]),
    .X(net105));
 sky130_fd_sc_hd__buf_2 _9307_ (.A(ch_data_in[50]),
    .X(net107));
 sky130_fd_sc_hd__buf_2 _9308_ (.A(ch_data_in[51]),
    .X(net108));
 sky130_fd_sc_hd__buf_2 _9309_ (.A(ch_data_in[52]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 _9310_ (.A(ch_data_in[53]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 _9311_ (.A(ch_data_in[54]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 _9312_ (.A(ch_data_in[55]),
    .X(net112));
 sky130_fd_sc_hd__buf_2 _9313_ (.A(ch_data_in[56]),
    .X(net113));
 sky130_fd_sc_hd__buf_2 _9314_ (.A(ch_data_in[57]),
    .X(net114));
 sky130_fd_sc_hd__buf_2 _9315_ (.A(ch_data_in[58]),
    .X(net115));
 sky130_fd_sc_hd__buf_2 _9316_ (.A(ch_data_in[59]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 _9317_ (.A(ch_data_in[60]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 _9318_ (.A(ch_data_in[61]),
    .X(net119));
 sky130_fd_sc_hd__buf_2 _9319_ (.A(ch_data_in[62]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 _9320_ (.A(ch_data_in[63]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 _9321_ (.A(ch_data_in[64]),
    .X(net122));
 sky130_fd_sc_hd__buf_2 _9322_ (.A(ch_data_in[65]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 _9323_ (.A(ch_data_in[66]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 _9324_ (.A(ch_data_in[67]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 _9325_ (.A(ch_data_in[68]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 _9326_ (.A(ch_data_in[69]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 _9327_ (.A(ch_data_in[70]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_2 _9328_ (.A(ch_data_in[71]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 _9329_ (.A(ch_data_in[72]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_2 _9330_ (.A(ch_data_in[73]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 _9331_ (.A(ch_data_in[74]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 _9332_ (.A(ch_data_in[75]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 _9333_ (.A(ch_data_in[76]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 _9334_ (.A(net1641),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 _9335_ (.A(net1639),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 _9336_ (.A(net1637),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 _9337_ (.A(net1635),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 _9338_ (.A(net1633),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 _9339_ (.A(net1631),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 _9340_ (.A(net1629),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 _9341_ (.A(net1627),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 _9342_ (.A(net1625),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 _9343_ (.A(net1623),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 _9344_ (.A(net1621),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 _9345_ (.A(net1619),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 _9346_ (.A(net1617),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 _9347_ (.A(net1615),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 _9348_ (.A(net1613),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 _9349_ (.A(net1611),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 _9350_ (.A(net1609),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 _9351_ (.A(net1607),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_2 _9352_ (.A(net1605),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 _9353_ (.A(net1603),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_2 _9354_ (.A(net1601),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_2 _9355_ (.A(net1600),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_2 _9356_ (.A(net1599),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_2 _9357_ (.A(net1713),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 _9358_ (.A(net1711),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 _9359_ (.A(net1709),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 _9360_ (.A(net1707),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 _9361_ (.A(net1705),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 _9362_ (.A(net1703),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 _9363_ (.A(net1701),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 _9364_ (.A(net1699),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 _9365_ (.A(net1697),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 _9366_ (.A(net1695),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 _9367_ (.A(net1693),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 _9368_ (.A(net1691),
    .X(net17));
 sky130_fd_sc_hd__buf_6 _9369_ (.A(ch_data_in[112]),
    .X(net18));
 sky130_fd_sc_hd__buf_6 _9370_ (.A(ch_data_in[113]),
    .X(net19));
 sky130_fd_sc_hd__buf_6 _9371_ (.A(ch_data_in[114]),
    .X(net20));
 sky130_fd_sc_hd__buf_6 _9372_ (.A(ch_data_in[115]),
    .X(net21));
 sky130_fd_sc_hd__buf_6 _9373_ (.A(ch_data_in[116]),
    .X(net22));
 sky130_fd_sc_hd__buf_6 _9374_ (.A(ch_data_in[117]),
    .X(net23));
 sky130_fd_sc_hd__buf_6 _9375_ (.A(ch_data_in[118]),
    .X(net24));
 sky130_fd_sc_hd__buf_6 _9376_ (.A(ch_data_in[119]),
    .X(net25));
 sky130_fd_sc_hd__buf_6 _9377_ (.A(ch_data_in[120]),
    .X(net27));
 sky130_fd_sc_hd__buf_6 _9378_ (.A(ch_data_in[121]),
    .X(net28));
 sky130_fd_sc_hd__buf_6 _9379_ (.A(ch_data_in[122]),
    .X(net29));
 sky130_fd_sc_hd__buf_6 _9380_ (.A(ch_data_in[123]),
    .X(net30));
 sky130_fd_sc_hd__buf_6 _9381_ (.A(ch_data_in[124]),
    .X(net31));
 sky130_fd_sc_hd__buf_6 _9382_ (.A(ch_data_in[125]),
    .X(net32));
 sky130_fd_sc_hd__buf_6 _9383_ (.A(ch_data_in[126]),
    .X(net33));
 sky130_fd_sc_hd__buf_6 _9384_ (.A(ch_data_in[127]),
    .X(net34));
 sky130_fd_sc_hd__buf_6 _9385_ (.A(ch_data_in[128]),
    .X(net35));
 sky130_fd_sc_hd__buf_6 _9386_ (.A(ch_data_in[129]),
    .X(net36));
 sky130_fd_sc_hd__buf_6 _9387_ (.A(ch_data_in[130]),
    .X(net38));
 sky130_fd_sc_hd__buf_6 _9388_ (.A(ch_data_in[131]),
    .X(net39));
 sky130_fd_sc_hd__buf_6 _9389_ (.A(ch_data_in[132]),
    .X(net40));
 sky130_fd_sc_hd__buf_6 _9390_ (.A(ch_data_in[133]),
    .X(net41));
 sky130_fd_sc_hd__buf_6 _9391_ (.A(ch_data_in[134]),
    .X(net42));
 sky130_fd_sc_hd__buf_6 _9392_ (.A(ch_data_in[135]),
    .X(net43));
 sky130_fd_sc_hd__buf_6 _9393_ (.A(ch_data_in[136]),
    .X(net44));
 sky130_fd_sc_hd__buf_6 _9394_ (.A(ch_data_in[137]),
    .X(net45));
 sky130_fd_sc_hd__buf_4 _9395_ (.A(ch_data_in[138]),
    .X(net46));
 sky130_fd_sc_hd__buf_2 _9396_ (.A(net1688),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 _9397_ (.A(net1685),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 _9398_ (.A(net1684),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 _9399_ (.A(net1683),
    .X(net51));
 sky130_fd_sc_hd__buf_2 _9400_ (.A(net1682),
    .X(net52));
 sky130_fd_sc_hd__buf_6 _9401_ (.A(ch_data_in[144]),
    .X(net53));
 sky130_fd_sc_hd__buf_4 _9402_ (.A(ch_data_in[145]),
    .X(net54));
 sky130_fd_sc_hd__buf_6 _9403_ (.A(ch_data_in[146]),
    .X(net55));
 sky130_fd_sc_hd__buf_6 _9404_ (.A(ch_data_in[147]),
    .X(net56));
 sky130_fd_sc_hd__buf_6 _9405_ (.A(ch_data_in[148]),
    .X(net57));
 sky130_fd_sc_hd__buf_6 _9406_ (.A(ch_data_in[149]),
    .X(net58));
 sky130_fd_sc_hd__buf_2 _9407_ (.A(net1677),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_4 _9408_ (.A(net1674),
    .X(net61));
 sky130_fd_sc_hd__buf_6 _9409_ (.A(ch_data_in[152]),
    .X(net62));
 sky130_fd_sc_hd__buf_6 _9410_ (.A(ch_data_in[153]),
    .X(net63));
 sky130_fd_sc_hd__buf_6 _9411_ (.A(ch_data_in[154]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 _9412_ (.A(net1671),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 _9413_ (.A(net1668),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 _9414_ (.A(net1665),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 _9415_ (.A(net342),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_1 _9416_ (.A(net389),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_1 _9417_ (.A(net438),
    .X(net475));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_mclk_raw (.A(net1761),
    .X(clknet_0_mclk_raw));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_dsync.out_clk  (.A(net1733),
    .X(\clknet_0_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0_0_mclk_raw (.A(net1764),
    .X(clknet_1_0_0_mclk_raw));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0_0_u_dsync.out_clk  (.A(net1737),
    .X(\clknet_1_0_0_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1_0_mclk_raw (.A(net1765),
    .X(clknet_1_1_0_mclk_raw));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1_0_u_dsync.out_clk  (.A(net1736),
    .X(\clknet_1_1_0_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_mclk_raw (.A(clknet_1_0_0_mclk_raw),
    .X(clknet_2_0__leaf_mclk_raw));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_mclk_raw (.A(clknet_1_0_0_mclk_raw),
    .X(clknet_2_1__leaf_mclk_raw));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_mclk_raw (.A(clknet_1_1_0_mclk_raw),
    .X(clknet_2_2__leaf_mclk_raw));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_mclk_raw (.A(clknet_1_1_0_mclk_raw),
    .X(clknet_2_3__leaf_mclk_raw));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_0__f_u_dsync.out_clk  (.A(net1738),
    .X(\clknet_3_0__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_1__f_u_dsync.out_clk  (.A(net1739),
    .X(\clknet_3_1__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_2__f_u_dsync.out_clk  (.A(net1738),
    .X(\clknet_3_2__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_3__f_u_dsync.out_clk  (.A(net1739),
    .X(\clknet_3_3__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_4__f_u_dsync.out_clk  (.A(\clknet_1_1_0_u_dsync.out_clk ),
    .X(\clknet_3_4__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_5__f_u_dsync.out_clk  (.A(net1740),
    .X(\clknet_3_5__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_6__f_u_dsync.out_clk  (.A(net1741),
    .X(\clknet_3_6__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_7__f_u_dsync.out_clk  (.A(net1740),
    .X(\clknet_3_7__leaf_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_0_u_dsync.out_clk  (.A(net1742),
    .X(\clknet_leaf_0_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_100_u_dsync.out_clk  (.A(net1742),
    .X(\clknet_leaf_100_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_101_u_dsync.out_clk  (.A(net1742),
    .X(\clknet_leaf_101_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_102_u_dsync.out_clk  (.A(\clknet_3_0__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_102_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_103_u_dsync.out_clk  (.A(net1743),
    .X(\clknet_leaf_103_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_104_u_dsync.out_clk  (.A(net1744),
    .X(\clknet_leaf_104_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_105_u_dsync.out_clk  (.A(net1744),
    .X(\clknet_leaf_105_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_106_u_dsync.out_clk  (.A(\clknet_3_0__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_106_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_107_u_dsync.out_clk  (.A(\clknet_3_0__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_107_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_108_u_dsync.out_clk  (.A(net1743),
    .X(\clknet_leaf_108_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_109_u_dsync.out_clk  (.A(net1744),
    .X(\clknet_leaf_109_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_10_u_dsync.out_clk  (.A(net1753),
    .X(\clknet_leaf_10_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_11_u_dsync.out_clk  (.A(net1754),
    .X(\clknet_leaf_11_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_12_u_dsync.out_clk  (.A(\clknet_3_4__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_12_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_13_u_dsync.out_clk  (.A(net1754),
    .X(\clknet_leaf_13_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_14_u_dsync.out_clk  (.A(net1753),
    .X(\clknet_leaf_14_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_15_u_dsync.out_clk  (.A(net1753),
    .X(\clknet_leaf_15_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_16_u_dsync.out_clk  (.A(net1753),
    .X(\clknet_leaf_16_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_17_u_dsync.out_clk  (.A(net1754),
    .X(\clknet_leaf_17_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_18_u_dsync.out_clk  (.A(net1752),
    .X(\clknet_leaf_18_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_19_u_dsync.out_clk  (.A(net1752),
    .X(\clknet_leaf_19_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_1_u_dsync.out_clk  (.A(net1746),
    .X(\clknet_leaf_1_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_20_u_dsync.out_clk  (.A(net1752),
    .X(\clknet_leaf_20_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_21_u_dsync.out_clk  (.A(net1755),
    .X(\clknet_leaf_21_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_22_u_dsync.out_clk  (.A(\clknet_3_5__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_22_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_23_u_dsync.out_clk  (.A(net1757),
    .X(\clknet_leaf_23_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_24_u_dsync.out_clk  (.A(net1757),
    .X(\clknet_leaf_24_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_25_u_dsync.out_clk  (.A(net1757),
    .X(\clknet_leaf_25_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_26_u_dsync.out_clk  (.A(net1755),
    .X(\clknet_leaf_26_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_27_u_dsync.out_clk  (.A(net1755),
    .X(\clknet_leaf_27_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_28_u_dsync.out_clk  (.A(net1757),
    .X(\clknet_leaf_28_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_29_u_dsync.out_clk  (.A(net1756),
    .X(\clknet_leaf_29_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_2_u_dsync.out_clk  (.A(\clknet_3_1__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_2_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_30_u_dsync.out_clk  (.A(net1756),
    .X(\clknet_leaf_30_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_31_u_dsync.out_clk  (.A(net1756),
    .X(\clknet_leaf_31_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_32_u_dsync.out_clk  (.A(net1758),
    .X(\clknet_leaf_32_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_33_u_dsync.out_clk  (.A(net1755),
    .X(\clknet_leaf_33_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_34_u_dsync.out_clk  (.A(net1755),
    .X(\clknet_leaf_34_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_35_u_dsync.out_clk  (.A(\clknet_3_4__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_35_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_36_u_dsync.out_clk  (.A(net1759),
    .X(\clknet_leaf_36_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_37_u_dsync.out_clk  (.A(\clknet_3_6__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_37_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_38_u_dsync.out_clk  (.A(\clknet_3_6__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_38_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_39_u_dsync.out_clk  (.A(\clknet_3_6__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_39_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_3_u_dsync.out_clk  (.A(net1745),
    .X(\clknet_leaf_3_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_40_u_dsync.out_clk  (.A(net1759),
    .X(\clknet_leaf_40_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_41_u_dsync.out_clk  (.A(\clknet_3_6__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_41_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_42_u_dsync.out_clk  (.A(net1759),
    .X(\clknet_leaf_42_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_43_u_dsync.out_clk  (.A(net1758),
    .X(\clknet_leaf_43_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_44_u_dsync.out_clk  (.A(net1758),
    .X(\clknet_leaf_44_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_45_u_dsync.out_clk  (.A(net1757),
    .X(\clknet_leaf_45_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_46_u_dsync.out_clk  (.A(net1756),
    .X(\clknet_leaf_46_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_47_u_dsync.out_clk  (.A(net1756),
    .X(\clknet_leaf_47_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_48_u_dsync.out_clk  (.A(net1760),
    .X(\clknet_leaf_48_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_49_u_dsync.out_clk  (.A(\clknet_3_7__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_49_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_4_u_dsync.out_clk  (.A(net1745),
    .X(\clknet_leaf_4_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_50_u_dsync.out_clk  (.A(\clknet_3_7__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_50_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_51_u_dsync.out_clk  (.A(net1760),
    .X(\clknet_leaf_51_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_52_u_dsync.out_clk  (.A(net1760),
    .X(\clknet_leaf_52_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_53_u_dsync.out_clk  (.A(\clknet_3_7__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_53_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_54_u_dsync.out_clk  (.A(\clknet_3_7__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_54_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_55_u_dsync.out_clk  (.A(net1759),
    .X(\clknet_leaf_55_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_56_u_dsync.out_clk  (.A(\clknet_3_6__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_56_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_57_u_dsync.out_clk  (.A(\clknet_3_6__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_57_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_58_u_dsync.out_clk  (.A(\clknet_3_6__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_58_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_59_u_dsync.out_clk  (.A(\clknet_3_6__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_59_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_5_u_dsync.out_clk  (.A(\clknet_3_1__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_5_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_60_u_dsync.out_clk  (.A(\clknet_3_6__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_60_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_61_u_dsync.out_clk  (.A(\clknet_3_6__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_61_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_62_u_dsync.out_clk  (.A(\clknet_3_6__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_62_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_63_u_dsync.out_clk  (.A(\clknet_3_6__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_63_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_64_u_dsync.out_clk  (.A(\clknet_3_6__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_64_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_65_u_dsync.out_clk  (.A(\clknet_3_6__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_65_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_66_u_dsync.out_clk  (.A(net1750),
    .X(\clknet_leaf_66_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_67_u_dsync.out_clk  (.A(net1750),
    .X(\clknet_leaf_67_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_68_u_dsync.out_clk  (.A(net1750),
    .X(\clknet_leaf_68_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_69_u_dsync.out_clk  (.A(\clknet_3_3__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_69_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_6_u_dsync.out_clk  (.A(\clknet_3_1__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_6_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_70_u_dsync.out_clk  (.A(net1749),
    .X(\clknet_leaf_70_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_71_u_dsync.out_clk  (.A(net1751),
    .X(\clknet_leaf_71_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_72_u_dsync.out_clk  (.A(net1751),
    .X(\clknet_leaf_72_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_73_u_dsync.out_clk  (.A(net1751),
    .X(\clknet_leaf_73_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_74_u_dsync.out_clk  (.A(net1751),
    .X(\clknet_leaf_74_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_75_u_dsync.out_clk  (.A(\clknet_3_3__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_75_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_76_u_dsync.out_clk  (.A(net1749),
    .X(\clknet_leaf_76_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_77_u_dsync.out_clk  (.A(net1749),
    .X(\clknet_leaf_77_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_78_u_dsync.out_clk  (.A(net1748),
    .X(\clknet_leaf_78_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_79_u_dsync.out_clk  (.A(net1748),
    .X(\clknet_leaf_79_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_7_u_dsync.out_clk  (.A(net1745),
    .X(\clknet_leaf_7_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_80_u_dsync.out_clk  (.A(\clknet_3_2__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_80_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_81_u_dsync.out_clk  (.A(net1747),
    .X(\clknet_leaf_81_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_82_u_dsync.out_clk  (.A(net1747),
    .X(\clknet_leaf_82_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_83_u_dsync.out_clk  (.A(net1747),
    .X(\clknet_leaf_83_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_84_u_dsync.out_clk  (.A(net1747),
    .X(\clknet_leaf_84_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_85_u_dsync.out_clk  (.A(\clknet_3_2__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_85_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_86_u_dsync.out_clk  (.A(net1748),
    .X(\clknet_leaf_86_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_87_u_dsync.out_clk  (.A(\clknet_3_2__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_87_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_88_u_dsync.out_clk  (.A(net1747),
    .X(\clknet_leaf_88_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_89_u_dsync.out_clk  (.A(net1744),
    .X(\clknet_leaf_89_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_8_u_dsync.out_clk  (.A(net1745),
    .X(\clknet_leaf_8_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_90_u_dsync.out_clk  (.A(net1744),
    .X(\clknet_leaf_90_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_91_u_dsync.out_clk  (.A(net1742),
    .X(\clknet_leaf_91_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_92_u_dsync.out_clk  (.A(net1742),
    .X(\clknet_leaf_92_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_93_u_dsync.out_clk  (.A(net1749),
    .X(\clknet_leaf_93_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_94_u_dsync.out_clk  (.A(net1749),
    .X(\clknet_leaf_94_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_95_u_dsync.out_clk  (.A(\clknet_3_3__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_95_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_96_u_dsync.out_clk  (.A(net1745),
    .X(\clknet_leaf_96_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_97_u_dsync.out_clk  (.A(\clknet_3_1__leaf_u_dsync.out_clk ),
    .X(\clknet_leaf_97_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_98_u_dsync.out_clk  (.A(net1746),
    .X(\clknet_leaf_98_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_99_u_dsync.out_clk  (.A(net1746),
    .X(\clknet_leaf_99_u_dsync.out_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_9_u_dsync.out_clk  (.A(net1753),
    .X(\clknet_leaf_9_u_dsync.out_clk ));
 sky130_fd_sc_hd__buf_4 fanout1000 (.A(_2800_),
    .X(net1000));
 sky130_fd_sc_hd__clkbuf_4 fanout1001 (.A(_2800_),
    .X(net1001));
 sky130_fd_sc_hd__buf_4 fanout1002 (.A(net1004),
    .X(net1002));
 sky130_fd_sc_hd__clkbuf_4 fanout1003 (.A(net1004),
    .X(net1003));
 sky130_fd_sc_hd__buf_6 fanout1004 (.A(net1953),
    .X(net1004));
 sky130_fd_sc_hd__clkbuf_4 fanout1005 (.A(_2590_),
    .X(net1005));
 sky130_fd_sc_hd__clkbuf_2 fanout1006 (.A(_2590_),
    .X(net1006));
 sky130_fd_sc_hd__buf_2 fanout1143 (.A(net1144),
    .X(net1143));
 sky130_fd_sc_hd__buf_2 fanout1144 (.A(_2021_),
    .X(net1144));
 sky130_fd_sc_hd__clkbuf_4 fanout1145 (.A(net1147),
    .X(net1145));
 sky130_fd_sc_hd__clkbuf_2 fanout1146 (.A(net1147),
    .X(net1146));
 sky130_fd_sc_hd__clkbuf_2 fanout1147 (.A(_2021_),
    .X(net1147));
 sky130_fd_sc_hd__clkbuf_8 fanout1148 (.A(net1152),
    .X(net1148));
 sky130_fd_sc_hd__buf_4 fanout1149 (.A(net1151),
    .X(net1149));
 sky130_fd_sc_hd__buf_2 fanout1150 (.A(net1151),
    .X(net1150));
 sky130_fd_sc_hd__buf_4 fanout1151 (.A(net1152),
    .X(net1151));
 sky130_fd_sc_hd__buf_4 fanout1152 (.A(_2020_),
    .X(net1152));
 sky130_fd_sc_hd__clkbuf_4 fanout1153 (.A(net1156),
    .X(net1153));
 sky130_fd_sc_hd__clkbuf_2 fanout1154 (.A(net1156),
    .X(net1154));
 sky130_fd_sc_hd__clkbuf_4 fanout1155 (.A(net1156),
    .X(net1155));
 sky130_fd_sc_hd__buf_2 fanout1156 (.A(net1157),
    .X(net1156));
 sky130_fd_sc_hd__clkbuf_4 fanout1157 (.A(_2014_),
    .X(net1157));
 sky130_fd_sc_hd__buf_2 fanout1158 (.A(net1160),
    .X(net1158));
 sky130_fd_sc_hd__buf_2 fanout1159 (.A(net1160),
    .X(net1159));
 sky130_fd_sc_hd__buf_2 fanout1160 (.A(_2011_),
    .X(net1160));
 sky130_fd_sc_hd__clkbuf_4 fanout1161 (.A(_2011_),
    .X(net1161));
 sky130_fd_sc_hd__clkbuf_4 fanout1162 (.A(net1163),
    .X(net1162));
 sky130_fd_sc_hd__clkbuf_4 fanout1163 (.A(_2008_),
    .X(net1163));
 sky130_fd_sc_hd__clkbuf_4 fanout1164 (.A(_2008_),
    .X(net1164));
 sky130_fd_sc_hd__clkbuf_2 fanout1165 (.A(_2008_),
    .X(net1165));
 sky130_fd_sc_hd__buf_6 fanout1166 (.A(net1167),
    .X(net1166));
 sky130_fd_sc_hd__buf_6 fanout1167 (.A(net1171),
    .X(net1167));
 sky130_fd_sc_hd__clkbuf_4 fanout1168 (.A(net1169),
    .X(net1168));
 sky130_fd_sc_hd__clkbuf_4 fanout1169 (.A(net1170),
    .X(net1169));
 sky130_fd_sc_hd__clkbuf_4 fanout1170 (.A(net1171),
    .X(net1170));
 sky130_fd_sc_hd__buf_4 fanout1171 (.A(_1936_),
    .X(net1171));
 sky130_fd_sc_hd__clkbuf_4 fanout1172 (.A(net1173),
    .X(net1172));
 sky130_fd_sc_hd__buf_4 fanout1173 (.A(_1935_),
    .X(net1173));
 sky130_fd_sc_hd__buf_4 fanout1174 (.A(net1176),
    .X(net1174));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1175 (.A(net1176),
    .X(net1175));
 sky130_fd_sc_hd__buf_4 fanout1176 (.A(_1920_),
    .X(net1176));
 sky130_fd_sc_hd__clkbuf_4 fanout1177 (.A(net1178),
    .X(net1177));
 sky130_fd_sc_hd__buf_2 fanout1178 (.A(net1179),
    .X(net1178));
 sky130_fd_sc_hd__clkbuf_4 fanout1179 (.A(_1917_),
    .X(net1179));
 sky130_fd_sc_hd__buf_4 fanout1180 (.A(_1915_),
    .X(net1180));
 sky130_fd_sc_hd__buf_4 fanout1182 (.A(_1851_),
    .X(net1182));
 sky130_fd_sc_hd__clkbuf_4 fanout1183 (.A(_1833_),
    .X(net1183));
 sky130_fd_sc_hd__clkbuf_2 fanout1184 (.A(_1833_),
    .X(net1184));
 sky130_fd_sc_hd__clkbuf_4 fanout1185 (.A(net1186),
    .X(net1185));
 sky130_fd_sc_hd__clkbuf_8 fanout1186 (.A(_1832_),
    .X(net1186));
 sky130_fd_sc_hd__buf_6 fanout1187 (.A(net1188),
    .X(net1187));
 sky130_fd_sc_hd__buf_6 fanout1188 (.A(_1831_),
    .X(net1188));
 sky130_fd_sc_hd__buf_2 fanout1189 (.A(net1190),
    .X(net1189));
 sky130_fd_sc_hd__buf_2 fanout1190 (.A(net1191),
    .X(net1190));
 sky130_fd_sc_hd__clkbuf_4 fanout1191 (.A(_1831_),
    .X(net1191));
 sky130_fd_sc_hd__clkbuf_4 fanout1192 (.A(_1830_),
    .X(net1192));
 sky130_fd_sc_hd__buf_4 fanout1193 (.A(_1731_),
    .X(net1193));
 sky130_fd_sc_hd__clkbuf_4 fanout1194 (.A(net1196),
    .X(net1194));
 sky130_fd_sc_hd__clkbuf_2 fanout1195 (.A(net1196),
    .X(net1195));
 sky130_fd_sc_hd__clkbuf_4 fanout1196 (.A(net1198),
    .X(net1196));
 sky130_fd_sc_hd__clkbuf_4 fanout1197 (.A(net1198),
    .X(net1197));
 sky130_fd_sc_hd__clkbuf_4 fanout1198 (.A(_1730_),
    .X(net1198));
 sky130_fd_sc_hd__clkbuf_4 fanout1199 (.A(net1200),
    .X(net1199));
 sky130_fd_sc_hd__clkbuf_4 fanout1200 (.A(net1201),
    .X(net1200));
 sky130_fd_sc_hd__buf_4 fanout1201 (.A(_1730_),
    .X(net1201));
 sky130_fd_sc_hd__buf_2 fanout1202 (.A(net1203),
    .X(net1202));
 sky130_fd_sc_hd__buf_4 fanout1203 (.A(_1729_),
    .X(net1203));
 sky130_fd_sc_hd__clkbuf_4 fanout1204 (.A(net1205),
    .X(net1204));
 sky130_fd_sc_hd__buf_4 fanout1205 (.A(_1729_),
    .X(net1205));
 sky130_fd_sc_hd__buf_4 fanout1206 (.A(net1209),
    .X(net1206));
 sky130_fd_sc_hd__clkbuf_4 fanout1207 (.A(net1208),
    .X(net1207));
 sky130_fd_sc_hd__buf_4 fanout1208 (.A(net1209),
    .X(net1208));
 sky130_fd_sc_hd__buf_4 fanout1209 (.A(_1727_),
    .X(net1209));
 sky130_fd_sc_hd__clkbuf_4 fanout1210 (.A(net1218),
    .X(net1210));
 sky130_fd_sc_hd__buf_4 fanout1211 (.A(net1218),
    .X(net1211));
 sky130_fd_sc_hd__buf_2 fanout1212 (.A(net1218),
    .X(net1212));
 sky130_fd_sc_hd__clkbuf_4 fanout1213 (.A(net1214),
    .X(net1213));
 sky130_fd_sc_hd__clkbuf_2 fanout1214 (.A(net1217),
    .X(net1214));
 sky130_fd_sc_hd__clkbuf_4 fanout1215 (.A(net1217),
    .X(net1215));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1216 (.A(net1217),
    .X(net1216));
 sky130_fd_sc_hd__clkbuf_2 fanout1217 (.A(net1218),
    .X(net1217));
 sky130_fd_sc_hd__buf_4 fanout1218 (.A(_1708_),
    .X(net1218));
 sky130_fd_sc_hd__clkbuf_4 fanout1219 (.A(net1223),
    .X(net1219));
 sky130_fd_sc_hd__clkbuf_4 fanout1220 (.A(net1223),
    .X(net1220));
 sky130_fd_sc_hd__clkbuf_4 fanout1221 (.A(net1223),
    .X(net1221));
 sky130_fd_sc_hd__clkbuf_4 fanout1222 (.A(net1223),
    .X(net1222));
 sky130_fd_sc_hd__buf_6 fanout1223 (.A(_1707_),
    .X(net1223));
 sky130_fd_sc_hd__buf_4 fanout1224 (.A(_1677_),
    .X(net1224));
 sky130_fd_sc_hd__clkbuf_4 fanout1225 (.A(_1677_),
    .X(net1225));
 sky130_fd_sc_hd__clkbuf_4 fanout1226 (.A(net1231),
    .X(net1226));
 sky130_fd_sc_hd__clkbuf_2 fanout1227 (.A(net1231),
    .X(net1227));
 sky130_fd_sc_hd__clkbuf_4 fanout1228 (.A(net1231),
    .X(net1228));
 sky130_fd_sc_hd__clkbuf_4 fanout1229 (.A(net1230),
    .X(net1229));
 sky130_fd_sc_hd__clkbuf_4 fanout1230 (.A(net1231),
    .X(net1230));
 sky130_fd_sc_hd__buf_2 fanout1231 (.A(_1677_),
    .X(net1231));
 sky130_fd_sc_hd__buf_4 fanout1232 (.A(net1233),
    .X(net1232));
 sky130_fd_sc_hd__buf_4 fanout1233 (.A(net1238),
    .X(net1233));
 sky130_fd_sc_hd__buf_2 fanout1234 (.A(net1235),
    .X(net1234));
 sky130_fd_sc_hd__clkbuf_2 fanout1235 (.A(net1236),
    .X(net1235));
 sky130_fd_sc_hd__buf_2 fanout1236 (.A(net1237),
    .X(net1236));
 sky130_fd_sc_hd__clkbuf_4 fanout1237 (.A(net1238),
    .X(net1237));
 sky130_fd_sc_hd__buf_4 fanout1238 (.A(_1676_),
    .X(net1238));
 sky130_fd_sc_hd__buf_4 fanout1239 (.A(net1240),
    .X(net1239));
 sky130_fd_sc_hd__buf_4 fanout1240 (.A(_1673_),
    .X(net1240));
 sky130_fd_sc_hd__buf_2 fanout1241 (.A(net1242),
    .X(net1241));
 sky130_fd_sc_hd__clkbuf_2 fanout1242 (.A(net1243),
    .X(net1242));
 sky130_fd_sc_hd__clkbuf_4 fanout1243 (.A(_1673_),
    .X(net1243));
 sky130_fd_sc_hd__clkbuf_4 fanout1244 (.A(_1673_),
    .X(net1244));
 sky130_fd_sc_hd__buf_4 fanout1245 (.A(net1246),
    .X(net1245));
 sky130_fd_sc_hd__buf_4 fanout1246 (.A(net1252),
    .X(net1246));
 sky130_fd_sc_hd__buf_2 fanout1247 (.A(net1252),
    .X(net1247));
 sky130_fd_sc_hd__clkbuf_2 fanout1248 (.A(net1252),
    .X(net1248));
 sky130_fd_sc_hd__clkbuf_4 fanout1249 (.A(net1250),
    .X(net1249));
 sky130_fd_sc_hd__buf_2 fanout1250 (.A(net1251),
    .X(net1250));
 sky130_fd_sc_hd__buf_2 fanout1251 (.A(net1252),
    .X(net1251));
 sky130_fd_sc_hd__buf_4 fanout1252 (.A(_1672_),
    .X(net1252));
 sky130_fd_sc_hd__buf_2 fanout1253 (.A(net1254),
    .X(net1253));
 sky130_fd_sc_hd__buf_2 fanout1254 (.A(_1670_),
    .X(net1254));
 sky130_fd_sc_hd__buf_2 fanout1255 (.A(net1256),
    .X(net1255));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1256 (.A(net1257),
    .X(net1256));
 sky130_fd_sc_hd__clkbuf_2 fanout1257 (.A(net1258),
    .X(net1257));
 sky130_fd_sc_hd__clkbuf_4 fanout1258 (.A(_1670_),
    .X(net1258));
 sky130_fd_sc_hd__clkbuf_4 fanout1259 (.A(net1263),
    .X(net1259));
 sky130_fd_sc_hd__clkbuf_4 fanout1260 (.A(net1263),
    .X(net1260));
 sky130_fd_sc_hd__clkbuf_4 fanout1261 (.A(net1263),
    .X(net1261));
 sky130_fd_sc_hd__buf_4 fanout1262 (.A(net1263),
    .X(net1262));
 sky130_fd_sc_hd__clkbuf_4 fanout1263 (.A(_1670_),
    .X(net1263));
 sky130_fd_sc_hd__clkbuf_4 fanout1264 (.A(net1268),
    .X(net1264));
 sky130_fd_sc_hd__buf_2 fanout1265 (.A(net1266),
    .X(net1265));
 sky130_fd_sc_hd__clkbuf_2 fanout1266 (.A(net1267),
    .X(net1266));
 sky130_fd_sc_hd__clkbuf_2 fanout1267 (.A(net1268),
    .X(net1267));
 sky130_fd_sc_hd__clkbuf_4 fanout1268 (.A(_1669_),
    .X(net1268));
 sky130_fd_sc_hd__clkbuf_4 fanout1269 (.A(net1271),
    .X(net1269));
 sky130_fd_sc_hd__buf_2 fanout1270 (.A(net1271),
    .X(net1270));
 sky130_fd_sc_hd__buf_2 fanout1271 (.A(_1669_),
    .X(net1271));
 sky130_fd_sc_hd__buf_2 fanout1272 (.A(net1273),
    .X(net1272));
 sky130_fd_sc_hd__clkbuf_2 fanout1273 (.A(_1669_),
    .X(net1273));
 sky130_fd_sc_hd__clkbuf_4 fanout1274 (.A(net1275),
    .X(net1274));
 sky130_fd_sc_hd__buf_4 fanout1275 (.A(\u_wbi_arb.gnt[1] ),
    .X(net1275));
 sky130_fd_sc_hd__clkbuf_4 fanout1276 (.A(net1277),
    .X(net1276));
 sky130_fd_sc_hd__buf_2 fanout1277 (.A(net1278),
    .X(net1277));
 sky130_fd_sc_hd__clkbuf_4 fanout1278 (.A(\u_wbi_arb.gnt[0] ),
    .X(net1278));
 sky130_fd_sc_hd__buf_4 fanout1313 (.A(net1317),
    .X(net1313));
 sky130_fd_sc_hd__buf_2 fanout1314 (.A(net1317),
    .X(net1314));
 sky130_fd_sc_hd__buf_4 fanout1315 (.A(net1316),
    .X(net1315));
 sky130_fd_sc_hd__buf_4 fanout1316 (.A(net1317),
    .X(net1316));
 sky130_fd_sc_hd__clkbuf_4 fanout1317 (.A(\u_s0.u_sync_wbb.u_resp_if.rd_ptr[1] ),
    .X(net1317));
 sky130_fd_sc_hd__buf_6 fanout1318 (.A(net1322),
    .X(net1318));
 sky130_fd_sc_hd__clkbuf_4 fanout1319 (.A(net1322),
    .X(net1319));
 sky130_fd_sc_hd__buf_4 fanout1320 (.A(net1321),
    .X(net1320));
 sky130_fd_sc_hd__buf_6 fanout1321 (.A(net1322),
    .X(net1321));
 sky130_fd_sc_hd__buf_4 fanout1322 (.A(\u_s0.u_sync_wbb.u_resp_if.rd_ptr[0] ),
    .X(net1322));
 sky130_fd_sc_hd__buf_4 fanout1323 (.A(net1325),
    .X(net1323));
 sky130_fd_sc_hd__buf_4 fanout1324 (.A(net1325),
    .X(net1324));
 sky130_fd_sc_hd__clkbuf_4 fanout1325 (.A(net1332),
    .X(net1325));
 sky130_fd_sc_hd__buf_4 fanout1326 (.A(net1327),
    .X(net1326));
 sky130_fd_sc_hd__buf_4 fanout1327 (.A(net1332),
    .X(net1327));
 sky130_fd_sc_hd__buf_4 fanout1328 (.A(net1332),
    .X(net1328));
 sky130_fd_sc_hd__clkbuf_4 fanout1329 (.A(net1332),
    .X(net1329));
 sky130_fd_sc_hd__buf_4 fanout1330 (.A(net1332),
    .X(net1330));
 sky130_fd_sc_hd__clkbuf_4 fanout1331 (.A(net1332),
    .X(net1331));
 sky130_fd_sc_hd__buf_6 fanout1332 (.A(\u_s0.u_sync_wbb.u_cmd_if.rd_ptr[1] ),
    .X(net1332));
 sky130_fd_sc_hd__buf_6 fanout1333 (.A(net1335),
    .X(net1333));
 sky130_fd_sc_hd__buf_6 fanout1334 (.A(net1335),
    .X(net1334));
 sky130_fd_sc_hd__buf_4 fanout1335 (.A(net1342),
    .X(net1335));
 sky130_fd_sc_hd__buf_6 fanout1336 (.A(net1337),
    .X(net1336));
 sky130_fd_sc_hd__buf_6 fanout1337 (.A(net1342),
    .X(net1337));
 sky130_fd_sc_hd__buf_6 fanout1338 (.A(net1342),
    .X(net1338));
 sky130_fd_sc_hd__buf_4 fanout1339 (.A(net1342),
    .X(net1339));
 sky130_fd_sc_hd__buf_6 fanout1340 (.A(net1342),
    .X(net1340));
 sky130_fd_sc_hd__buf_4 fanout1341 (.A(net1342),
    .X(net1341));
 sky130_fd_sc_hd__buf_6 fanout1342 (.A(\u_s0.u_sync_wbb.u_cmd_if.rd_ptr[0] ),
    .X(net1342));
 sky130_fd_sc_hd__buf_4 fanout1343 (.A(net1344),
    .X(net1343));
 sky130_fd_sc_hd__buf_6 fanout1344 (.A(\u_s1.u_sync_wbb.u_resp_if.rd_ptr[1] ),
    .X(net1344));
 sky130_fd_sc_hd__buf_4 fanout1345 (.A(\u_s1.u_sync_wbb.u_resp_if.rd_ptr[1] ),
    .X(net1345));
 sky130_fd_sc_hd__buf_2 fanout1346 (.A(\u_s1.u_sync_wbb.u_resp_if.rd_ptr[1] ),
    .X(net1346));
 sky130_fd_sc_hd__buf_6 fanout1347 (.A(net1348),
    .X(net1347));
 sky130_fd_sc_hd__buf_6 fanout1348 (.A(net1351),
    .X(net1348));
 sky130_fd_sc_hd__buf_6 fanout1349 (.A(net1351),
    .X(net1349));
 sky130_fd_sc_hd__clkbuf_4 fanout1350 (.A(net1351),
    .X(net1350));
 sky130_fd_sc_hd__clkbuf_4 fanout1351 (.A(\u_s1.u_sync_wbb.u_resp_if.rd_ptr[0] ),
    .X(net1351));
 sky130_fd_sc_hd__buf_4 fanout1352 (.A(net1354),
    .X(net1352));
 sky130_fd_sc_hd__buf_4 fanout1353 (.A(net1354),
    .X(net1353));
 sky130_fd_sc_hd__clkbuf_4 fanout1354 (.A(\u_s1.u_sync_wbb.u_cmd_if.rd_ptr[1] ),
    .X(net1354));
 sky130_fd_sc_hd__buf_4 fanout1355 (.A(net1358),
    .X(net1355));
 sky130_fd_sc_hd__clkbuf_4 fanout1356 (.A(net1358),
    .X(net1356));
 sky130_fd_sc_hd__buf_4 fanout1357 (.A(net1358),
    .X(net1357));
 sky130_fd_sc_hd__clkbuf_4 fanout1358 (.A(\u_s1.u_sync_wbb.u_cmd_if.rd_ptr[1] ),
    .X(net1358));
 sky130_fd_sc_hd__buf_6 fanout1359 (.A(net1361),
    .X(net1359));
 sky130_fd_sc_hd__buf_6 fanout1360 (.A(net1361),
    .X(net1360));
 sky130_fd_sc_hd__clkbuf_8 fanout1361 (.A(\u_s1.u_sync_wbb.u_cmd_if.rd_ptr[0] ),
    .X(net1361));
 sky130_fd_sc_hd__clkbuf_8 fanout1362 (.A(net1365),
    .X(net1362));
 sky130_fd_sc_hd__clkbuf_8 fanout1363 (.A(net1365),
    .X(net1363));
 sky130_fd_sc_hd__buf_6 fanout1364 (.A(net1365),
    .X(net1364));
 sky130_fd_sc_hd__buf_4 fanout1365 (.A(\u_s1.u_sync_wbb.u_cmd_if.rd_ptr[0] ),
    .X(net1365));
 sky130_fd_sc_hd__buf_2 fanout1368 (.A(net1370),
    .X(net1368));
 sky130_fd_sc_hd__clkbuf_2 fanout1369 (.A(net1370),
    .X(net1369));
 sky130_fd_sc_hd__clkbuf_2 fanout1370 (.A(net1371),
    .X(net1370));
 sky130_fd_sc_hd__clkbuf_4 fanout1371 (.A(\u_s0.gnt[1] ),
    .X(net1371));
 sky130_fd_sc_hd__buf_2 fanout1372 (.A(net1374),
    .X(net1372));
 sky130_fd_sc_hd__clkbuf_1 fanout1373 (.A(net1374),
    .X(net1373));
 sky130_fd_sc_hd__clkbuf_2 fanout1374 (.A(\u_s0.gnt[0] ),
    .X(net1374));
 sky130_fd_sc_hd__buf_2 fanout1375 (.A(\u_s0.gnt[0] ),
    .X(net1375));
 sky130_fd_sc_hd__buf_6 fanout1376 (.A(\u_s2.u_sync_wbb.u_resp_if.rd_ptr[1] ),
    .X(net1376));
 sky130_fd_sc_hd__clkbuf_4 fanout1377 (.A(\u_s2.u_sync_wbb.u_resp_if.rd_ptr[1] ),
    .X(net1377));
 sky130_fd_sc_hd__buf_4 fanout1378 (.A(net1379),
    .X(net1378));
 sky130_fd_sc_hd__buf_6 fanout1379 (.A(\u_s2.u_sync_wbb.u_resp_if.rd_ptr[1] ),
    .X(net1379));
 sky130_fd_sc_hd__buf_8 fanout1380 (.A(net1384),
    .X(net1380));
 sky130_fd_sc_hd__buf_4 fanout1381 (.A(net1384),
    .X(net1381));
 sky130_fd_sc_hd__buf_6 fanout1382 (.A(net1383),
    .X(net1382));
 sky130_fd_sc_hd__buf_8 fanout1383 (.A(net1384),
    .X(net1383));
 sky130_fd_sc_hd__buf_4 fanout1384 (.A(\u_s2.u_sync_wbb.u_resp_if.rd_ptr[0] ),
    .X(net1384));
 sky130_fd_sc_hd__buf_4 fanout1385 (.A(\u_s2.u_sync_wbb.u_cmd_if.rd_ptr[1] ),
    .X(net1385));
 sky130_fd_sc_hd__clkbuf_4 fanout1386 (.A(\u_s2.u_sync_wbb.u_cmd_if.rd_ptr[1] ),
    .X(net1386));
 sky130_fd_sc_hd__buf_4 fanout1387 (.A(net1388),
    .X(net1387));
 sky130_fd_sc_hd__clkbuf_4 fanout1388 (.A(\u_s2.u_sync_wbb.u_cmd_if.rd_ptr[1] ),
    .X(net1388));
 sky130_fd_sc_hd__buf_4 fanout1389 (.A(net1391),
    .X(net1389));
 sky130_fd_sc_hd__buf_4 fanout1390 (.A(net1391),
    .X(net1390));
 sky130_fd_sc_hd__buf_4 fanout1391 (.A(\u_s2.u_sync_wbb.u_cmd_if.rd_ptr[1] ),
    .X(net1391));
 sky130_fd_sc_hd__buf_6 fanout1392 (.A(net1399),
    .X(net1392));
 sky130_fd_sc_hd__buf_4 fanout1393 (.A(net1399),
    .X(net1393));
 sky130_fd_sc_hd__buf_6 fanout1394 (.A(net1395),
    .X(net1394));
 sky130_fd_sc_hd__buf_4 fanout1395 (.A(net1399),
    .X(net1395));
 sky130_fd_sc_hd__buf_6 fanout1396 (.A(net1399),
    .X(net1396));
 sky130_fd_sc_hd__buf_6 fanout1397 (.A(net1399),
    .X(net1397));
 sky130_fd_sc_hd__clkbuf_4 fanout1398 (.A(net1399),
    .X(net1398));
 sky130_fd_sc_hd__buf_6 fanout1399 (.A(\u_s2.u_sync_wbb.u_cmd_if.rd_ptr[0] ),
    .X(net1399));
 sky130_fd_sc_hd__buf_8 fanout1400 (.A(\u_s2.u_sync_wbb.wbm_lack_o ),
    .X(net1400));
 sky130_fd_sc_hd__clkbuf_4 fanout1404 (.A(\u_s1.gnt[1] ),
    .X(net1404));
 sky130_fd_sc_hd__buf_4 fanout1405 (.A(\u_s1.gnt[0] ),
    .X(net1405));
 sky130_fd_sc_hd__clkbuf_2 fanout1406 (.A(\u_s1.gnt[0] ),
    .X(net1406));
 sky130_fd_sc_hd__buf_2 fanout1407 (.A(net1408),
    .X(net1407));
 sky130_fd_sc_hd__buf_4 fanout1408 (.A(\u_s2.gnt[1] ),
    .X(net1408));
 sky130_fd_sc_hd__clkbuf_4 fanout1409 (.A(net1410),
    .X(net1409));
 sky130_fd_sc_hd__clkbuf_4 fanout1410 (.A(\u_s2.gnt[0] ),
    .X(net1410));
 sky130_fd_sc_hd__buf_6 fanout1495 (.A(net1498),
    .X(net1495));
 sky130_fd_sc_hd__buf_4 fanout1496 (.A(net1498),
    .X(net1496));
 sky130_fd_sc_hd__buf_2 fanout1497 (.A(net1498),
    .X(net1497));
 sky130_fd_sc_hd__buf_4 fanout1498 (.A(net1784),
    .X(net1498));
 sky130_fd_sc_hd__clkbuf_8 fanout1499 (.A(net1784),
    .X(net1499));
 sky130_fd_sc_hd__buf_4 fanout1500 (.A(net1784),
    .X(net1500));
 sky130_fd_sc_hd__buf_4 fanout1501 (.A(net1502),
    .X(net1501));
 sky130_fd_sc_hd__clkbuf_4 fanout1502 (.A(net1784),
    .X(net1502));
 sky130_fd_sc_hd__buf_4 fanout1503 (.A(net1504),
    .X(net1503));
 sky130_fd_sc_hd__buf_2 fanout1504 (.A(net1510),
    .X(net1504));
 sky130_fd_sc_hd__buf_4 fanout1505 (.A(net1510),
    .X(net1505));
 sky130_fd_sc_hd__buf_2 fanout1506 (.A(net1510),
    .X(net1506));
 sky130_fd_sc_hd__buf_4 fanout1507 (.A(net1508),
    .X(net1507));
 sky130_fd_sc_hd__buf_4 fanout1508 (.A(net1509),
    .X(net1508));
 sky130_fd_sc_hd__buf_6 fanout1509 (.A(net1510),
    .X(net1509));
 sky130_fd_sc_hd__clkbuf_4 fanout1510 (.A(net2047),
    .X(net1510));
 sky130_fd_sc_hd__buf_6 fanout481 (.A(_2789_),
    .X(net481));
 sky130_fd_sc_hd__clkbuf_4 fanout482 (.A(_2789_),
    .X(net482));
 sky130_fd_sc_hd__buf_4 fanout483 (.A(_2789_),
    .X(net483));
 sky130_fd_sc_hd__clkbuf_4 fanout484 (.A(_2789_),
    .X(net484));
 sky130_fd_sc_hd__clkbuf_8 fanout486 (.A(_3362_),
    .X(net486));
 sky130_fd_sc_hd__clkbuf_2 fanout487 (.A(_3362_),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_4 fanout488 (.A(net489),
    .X(net488));
 sky130_fd_sc_hd__buf_4 fanout489 (.A(_3278_),
    .X(net489));
 sky130_fd_sc_hd__buf_4 fanout490 (.A(net493),
    .X(net490));
 sky130_fd_sc_hd__buf_4 fanout491 (.A(net493),
    .X(net491));
 sky130_fd_sc_hd__buf_6 fanout492 (.A(net493),
    .X(net492));
 sky130_fd_sc_hd__buf_4 fanout493 (.A(_3251_),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_8 fanout494 (.A(_3131_),
    .X(net494));
 sky130_fd_sc_hd__buf_2 fanout495 (.A(_3131_),
    .X(net495));
 sky130_fd_sc_hd__buf_4 fanout496 (.A(net497),
    .X(net496));
 sky130_fd_sc_hd__buf_6 fanout497 (.A(_3131_),
    .X(net497));
 sky130_fd_sc_hd__clkbuf_8 fanout498 (.A(_2788_),
    .X(net498));
 sky130_fd_sc_hd__buf_2 fanout499 (.A(_2788_),
    .X(net499));
 sky130_fd_sc_hd__buf_6 fanout500 (.A(_2788_),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_4 fanout501 (.A(_2788_),
    .X(net501));
 sky130_fd_sc_hd__buf_4 fanout502 (.A(net503),
    .X(net502));
 sky130_fd_sc_hd__buf_4 fanout503 (.A(_2787_),
    .X(net503));
 sky130_fd_sc_hd__buf_6 fanout504 (.A(_2787_),
    .X(net504));
 sky130_fd_sc_hd__buf_2 fanout505 (.A(_2787_),
    .X(net505));
 sky130_fd_sc_hd__buf_6 fanout506 (.A(net509),
    .X(net506));
 sky130_fd_sc_hd__buf_6 fanout507 (.A(net509),
    .X(net507));
 sky130_fd_sc_hd__clkbuf_4 fanout508 (.A(net509),
    .X(net508));
 sky130_fd_sc_hd__buf_4 fanout509 (.A(_2785_),
    .X(net509));
 sky130_fd_sc_hd__clkbuf_4 fanout513 (.A(_2593_),
    .X(net513));
 sky130_fd_sc_hd__clkbuf_2 fanout514 (.A(_2593_),
    .X(net514));
 sky130_fd_sc_hd__buf_6 fanout518 (.A(_3432_),
    .X(net518));
 sky130_fd_sc_hd__buf_4 fanout521 (.A(net524),
    .X(net521));
 sky130_fd_sc_hd__buf_4 fanout522 (.A(net524),
    .X(net522));
 sky130_fd_sc_hd__clkbuf_8 fanout523 (.A(net524),
    .X(net523));
 sky130_fd_sc_hd__buf_4 fanout524 (.A(_3254_),
    .X(net524));
 sky130_fd_sc_hd__buf_4 fanout525 (.A(net528),
    .X(net525));
 sky130_fd_sc_hd__buf_4 fanout526 (.A(net528),
    .X(net526));
 sky130_fd_sc_hd__clkbuf_8 fanout527 (.A(net528),
    .X(net527));
 sky130_fd_sc_hd__clkbuf_4 fanout528 (.A(_3253_),
    .X(net528));
 sky130_fd_sc_hd__buf_4 fanout529 (.A(net530),
    .X(net529));
 sky130_fd_sc_hd__buf_4 fanout530 (.A(net532),
    .X(net530));
 sky130_fd_sc_hd__buf_6 fanout531 (.A(net532),
    .X(net531));
 sky130_fd_sc_hd__buf_4 fanout532 (.A(_3252_),
    .X(net532));
 sky130_fd_sc_hd__clkbuf_8 fanout533 (.A(net536),
    .X(net533));
 sky130_fd_sc_hd__buf_4 fanout534 (.A(net536),
    .X(net534));
 sky130_fd_sc_hd__buf_4 fanout535 (.A(net536),
    .X(net535));
 sky130_fd_sc_hd__buf_4 fanout536 (.A(_3130_),
    .X(net536));
 sky130_fd_sc_hd__buf_4 fanout537 (.A(net540),
    .X(net537));
 sky130_fd_sc_hd__buf_4 fanout538 (.A(net539),
    .X(net538));
 sky130_fd_sc_hd__buf_4 fanout539 (.A(net540),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_4 fanout540 (.A(_3129_),
    .X(net540));
 sky130_fd_sc_hd__clkbuf_8 fanout541 (.A(_3128_),
    .X(net541));
 sky130_fd_sc_hd__buf_2 fanout542 (.A(_3128_),
    .X(net542));
 sky130_fd_sc_hd__buf_6 fanout543 (.A(_3128_),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_4 fanout544 (.A(_3128_),
    .X(net544));
 sky130_fd_sc_hd__clkbuf_4 fanout545 (.A(_2780_),
    .X(net545));
 sky130_fd_sc_hd__buf_2 fanout546 (.A(net549),
    .X(net546));
 sky130_fd_sc_hd__buf_4 fanout547 (.A(net548),
    .X(net547));
 sky130_fd_sc_hd__buf_4 fanout548 (.A(net549),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_4 fanout562 (.A(net563),
    .X(net562));
 sky130_fd_sc_hd__buf_4 fanout563 (.A(net564),
    .X(net563));
 sky130_fd_sc_hd__buf_2 fanout564 (.A(net566),
    .X(net564));
 sky130_fd_sc_hd__clkbuf_4 fanout565 (.A(net566),
    .X(net565));
 sky130_fd_sc_hd__buf_2 fanout566 (.A(net571),
    .X(net566));
 sky130_fd_sc_hd__buf_4 fanout567 (.A(net568),
    .X(net567));
 sky130_fd_sc_hd__buf_4 fanout568 (.A(net571),
    .X(net568));
 sky130_fd_sc_hd__buf_4 fanout569 (.A(net571),
    .X(net569));
 sky130_fd_sc_hd__buf_4 fanout570 (.A(net571),
    .X(net570));
 sky130_fd_sc_hd__clkbuf_8 fanout571 (.A(_2418_),
    .X(net571));
 sky130_fd_sc_hd__buf_6 fanout574 (.A(net579),
    .X(net574));
 sky130_fd_sc_hd__buf_6 fanout576 (.A(net578),
    .X(net576));
 sky130_fd_sc_hd__clkbuf_4 fanout577 (.A(net578),
    .X(net577));
 sky130_fd_sc_hd__buf_6 fanout578 (.A(_0009_),
    .X(net578));
 sky130_fd_sc_hd__clkbuf_4 fanout580 (.A(net581),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_4 fanout581 (.A(_1998_),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_4 fanout582 (.A(net583),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_2 fanout583 (.A(net584),
    .X(net583));
 sky130_fd_sc_hd__clkbuf_2 fanout584 (.A(_1992_),
    .X(net584));
 sky130_fd_sc_hd__buf_4 fanout586 (.A(net587),
    .X(net586));
 sky130_fd_sc_hd__clkbuf_8 fanout587 (.A(_2775_),
    .X(net587));
 sky130_fd_sc_hd__buf_4 fanout588 (.A(net589),
    .X(net588));
 sky130_fd_sc_hd__buf_6 fanout589 (.A(net591),
    .X(net589));
 sky130_fd_sc_hd__buf_4 fanout593 (.A(_2748_),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_4 fanout594 (.A(net597),
    .X(net594));
 sky130_fd_sc_hd__buf_4 fanout595 (.A(net596),
    .X(net595));
 sky130_fd_sc_hd__buf_6 fanout596 (.A(net597),
    .X(net596));
 sky130_fd_sc_hd__clkbuf_8 fanout598 (.A(_2744_),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_4 fanout599 (.A(net602),
    .X(net599));
 sky130_fd_sc_hd__buf_6 fanout600 (.A(net602),
    .X(net600));
 sky130_fd_sc_hd__buf_4 fanout601 (.A(net602),
    .X(net601));
 sky130_fd_sc_hd__buf_6 fanout603 (.A(net608),
    .X(net603));
 sky130_fd_sc_hd__buf_4 fanout604 (.A(net606),
    .X(net604));
 sky130_fd_sc_hd__buf_4 fanout605 (.A(net607),
    .X(net605));
 sky130_fd_sc_hd__clkbuf_1 fanout606 (.A(net608),
    .X(net606));
 sky130_fd_sc_hd__buf_4 fanout608 (.A(_2738_),
    .X(net608));
 sky130_fd_sc_hd__buf_6 fanout610 (.A(net614),
    .X(net610));
 sky130_fd_sc_hd__buf_4 fanout611 (.A(net612),
    .X(net611));
 sky130_fd_sc_hd__buf_6 fanout612 (.A(net616),
    .X(net612));
 sky130_fd_sc_hd__buf_6 fanout614 (.A(_2691_),
    .X(net614));
 sky130_fd_sc_hd__buf_2 fanout618 (.A(net620),
    .X(net618));
 sky130_fd_sc_hd__clkbuf_4 fanout619 (.A(net620),
    .X(net619));
 sky130_fd_sc_hd__clkbuf_4 fanout620 (.A(_2665_),
    .X(net620));
 sky130_fd_sc_hd__buf_4 fanout621 (.A(_2663_),
    .X(net621));
 sky130_fd_sc_hd__clkbuf_4 fanout622 (.A(net625),
    .X(net622));
 sky130_fd_sc_hd__buf_4 fanout623 (.A(net624),
    .X(net623));
 sky130_fd_sc_hd__buf_6 fanout624 (.A(net625),
    .X(net624));
 sky130_fd_sc_hd__buf_4 fanout626 (.A(_2024_),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_2 fanout627 (.A(net628),
    .X(net627));
 sky130_fd_sc_hd__buf_4 fanout713 (.A(net718),
    .X(net713));
 sky130_fd_sc_hd__buf_4 fanout714 (.A(net715),
    .X(net714));
 sky130_fd_sc_hd__clkbuf_4 fanout715 (.A(net718),
    .X(net715));
 sky130_fd_sc_hd__buf_6 fanout716 (.A(net717),
    .X(net716));
 sky130_fd_sc_hd__buf_8 fanout717 (.A(net718),
    .X(net717));
 sky130_fd_sc_hd__buf_6 fanout718 (.A(_2003_),
    .X(net718));
 sky130_fd_sc_hd__clkbuf_4 fanout721 (.A(_1960_),
    .X(net721));
 sky130_fd_sc_hd__clkbuf_2 fanout722 (.A(_1960_),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_4 fanout723 (.A(_1960_),
    .X(net723));
 sky130_fd_sc_hd__clkbuf_2 fanout724 (.A(_1960_),
    .X(net724));
 sky130_fd_sc_hd__buf_2 fanout733 (.A(net734),
    .X(net733));
 sky130_fd_sc_hd__buf_2 fanout734 (.A(_1769_),
    .X(net734));
 sky130_fd_sc_hd__clkbuf_4 fanout735 (.A(_1769_),
    .X(net735));
 sky130_fd_sc_hd__buf_2 fanout736 (.A(_1769_),
    .X(net736));
 sky130_fd_sc_hd__buf_4 fanout739 (.A(net741),
    .X(net739));
 sky130_fd_sc_hd__buf_4 fanout740 (.A(net741),
    .X(net740));
 sky130_fd_sc_hd__buf_4 fanout741 (.A(net748),
    .X(net741));
 sky130_fd_sc_hd__buf_4 fanout742 (.A(net743),
    .X(net742));
 sky130_fd_sc_hd__buf_4 fanout743 (.A(net748),
    .X(net743));
 sky130_fd_sc_hd__buf_4 fanout744 (.A(net748),
    .X(net744));
 sky130_fd_sc_hd__buf_2 fanout745 (.A(net748),
    .X(net745));
 sky130_fd_sc_hd__buf_4 fanout746 (.A(net747),
    .X(net746));
 sky130_fd_sc_hd__buf_4 fanout747 (.A(net748),
    .X(net747));
 sky130_fd_sc_hd__buf_4 fanout748 (.A(_3420_),
    .X(net748));
 sky130_fd_sc_hd__buf_4 fanout749 (.A(net750),
    .X(net749));
 sky130_fd_sc_hd__buf_4 fanout750 (.A(net751),
    .X(net750));
 sky130_fd_sc_hd__buf_4 fanout751 (.A(_2944_),
    .X(net751));
 sky130_fd_sc_hd__buf_4 fanout752 (.A(net755),
    .X(net752));
 sky130_fd_sc_hd__buf_2 fanout753 (.A(net755),
    .X(net753));
 sky130_fd_sc_hd__buf_4 fanout754 (.A(net755),
    .X(net754));
 sky130_fd_sc_hd__clkbuf_4 fanout755 (.A(_2944_),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_4 fanout756 (.A(net759),
    .X(net756));
 sky130_fd_sc_hd__buf_2 fanout757 (.A(net758),
    .X(net757));
 sky130_fd_sc_hd__clkbuf_4 fanout758 (.A(net759),
    .X(net758));
 sky130_fd_sc_hd__buf_2 fanout759 (.A(_2501_),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_4 fanout760 (.A(net763),
    .X(net760));
 sky130_fd_sc_hd__buf_2 fanout761 (.A(net762),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_4 fanout762 (.A(net763),
    .X(net762));
 sky130_fd_sc_hd__clkbuf_4 fanout763 (.A(_2495_),
    .X(net763));
 sky130_fd_sc_hd__clkbuf_4 fanout764 (.A(net765),
    .X(net764));
 sky130_fd_sc_hd__clkbuf_4 fanout765 (.A(_2259_),
    .X(net765));
 sky130_fd_sc_hd__clkbuf_4 fanout766 (.A(net1776),
    .X(net766));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout767 (.A(net1776),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_4 fanout768 (.A(_2189_),
    .X(net768));
 sky130_fd_sc_hd__clkbuf_2 fanout769 (.A(_2189_),
    .X(net769));
 sky130_fd_sc_hd__clkbuf_4 fanout770 (.A(_2189_),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_2 fanout771 (.A(_2189_),
    .X(net771));
 sky130_fd_sc_hd__buf_4 fanout772 (.A(net773),
    .X(net772));
 sky130_fd_sc_hd__buf_2 fanout773 (.A(net778),
    .X(net773));
 sky130_fd_sc_hd__buf_4 fanout774 (.A(net778),
    .X(net774));
 sky130_fd_sc_hd__buf_4 fanout775 (.A(net777),
    .X(net775));
 sky130_fd_sc_hd__buf_2 fanout776 (.A(net777),
    .X(net776));
 sky130_fd_sc_hd__buf_4 fanout777 (.A(net778),
    .X(net777));
 sky130_fd_sc_hd__buf_4 fanout778 (.A(_2005_),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_4 fanout779 (.A(net780),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_4 fanout780 (.A(_1956_),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_4 fanout781 (.A(net1775),
    .X(net781));
 sky130_fd_sc_hd__clkbuf_2 fanout782 (.A(net1775),
    .X(net782));
 sky130_fd_sc_hd__clkbuf_4 fanout799 (.A(net800),
    .X(net799));
 sky130_fd_sc_hd__buf_2 fanout800 (.A(_1855_),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_4 fanout801 (.A(net1774),
    .X(net801));
 sky130_fd_sc_hd__clkbuf_2 fanout802 (.A(net1774),
    .X(net802));
 sky130_fd_sc_hd__clkbuf_4 fanout803 (.A(_1852_),
    .X(net803));
 sky130_fd_sc_hd__clkbuf_2 fanout804 (.A(_1852_),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_4 fanout805 (.A(_1852_),
    .X(net805));
 sky130_fd_sc_hd__clkbuf_2 fanout806 (.A(_1852_),
    .X(net806));
 sky130_fd_sc_hd__buf_2 fanout808 (.A(_1800_),
    .X(net808));
 sky130_fd_sc_hd__buf_2 fanout809 (.A(net810),
    .X(net809));
 sky130_fd_sc_hd__buf_2 fanout810 (.A(_1780_),
    .X(net810));
 sky130_fd_sc_hd__clkbuf_4 fanout811 (.A(net812),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_4 fanout812 (.A(_1780_),
    .X(net812));
 sky130_fd_sc_hd__buf_8 fanout813 (.A(net814),
    .X(net813));
 sky130_fd_sc_hd__buf_6 fanout814 (.A(_1757_),
    .X(net814));
 sky130_fd_sc_hd__clkbuf_4 fanout815 (.A(_1757_),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_2 fanout816 (.A(_1757_),
    .X(net816));
 sky130_fd_sc_hd__buf_2 fanout817 (.A(net818),
    .X(net817));
 sky130_fd_sc_hd__buf_2 fanout818 (.A(net820),
    .X(net818));
 sky130_fd_sc_hd__clkbuf_4 fanout819 (.A(net820),
    .X(net819));
 sky130_fd_sc_hd__buf_2 fanout820 (.A(_1747_),
    .X(net820));
 sky130_fd_sc_hd__buf_2 fanout821 (.A(net822),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_4 fanout822 (.A(net823),
    .X(net822));
 sky130_fd_sc_hd__buf_4 fanout823 (.A(_1724_),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_4 fanout824 (.A(net825),
    .X(net824));
 sky130_fd_sc_hd__buf_4 fanout825 (.A(net826),
    .X(net825));
 sky130_fd_sc_hd__buf_2 fanout826 (.A(net833),
    .X(net826));
 sky130_fd_sc_hd__buf_4 fanout827 (.A(net828),
    .X(net827));
 sky130_fd_sc_hd__clkbuf_2 fanout828 (.A(net833),
    .X(net828));
 sky130_fd_sc_hd__buf_4 fanout829 (.A(net830),
    .X(net829));
 sky130_fd_sc_hd__buf_4 fanout830 (.A(net833),
    .X(net830));
 sky130_fd_sc_hd__buf_4 fanout831 (.A(net832),
    .X(net831));
 sky130_fd_sc_hd__buf_6 fanout832 (.A(net833),
    .X(net832));
 sky130_fd_sc_hd__buf_4 fanout833 (.A(_1718_),
    .X(net833));
 sky130_fd_sc_hd__buf_4 fanout834 (.A(net836),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_2 fanout835 (.A(net836),
    .X(net835));
 sky130_fd_sc_hd__buf_4 fanout836 (.A(net837),
    .X(net836));
 sky130_fd_sc_hd__buf_4 fanout837 (.A(net845),
    .X(net837));
 sky130_fd_sc_hd__buf_4 fanout838 (.A(net839),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_2 fanout839 (.A(net845),
    .X(net839));
 sky130_fd_sc_hd__buf_4 fanout840 (.A(net841),
    .X(net840));
 sky130_fd_sc_hd__buf_4 fanout841 (.A(net845),
    .X(net841));
 sky130_fd_sc_hd__buf_4 fanout842 (.A(net843),
    .X(net842));
 sky130_fd_sc_hd__clkbuf_4 fanout843 (.A(net844),
    .X(net843));
 sky130_fd_sc_hd__clkbuf_4 fanout844 (.A(net845),
    .X(net844));
 sky130_fd_sc_hd__buf_4 fanout845 (.A(net866),
    .X(net845));
 sky130_fd_sc_hd__buf_4 fanout846 (.A(net847),
    .X(net846));
 sky130_fd_sc_hd__buf_4 fanout847 (.A(net853),
    .X(net847));
 sky130_fd_sc_hd__buf_4 fanout848 (.A(net850),
    .X(net848));
 sky130_fd_sc_hd__buf_2 fanout849 (.A(net850),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_4 fanout850 (.A(net853),
    .X(net850));
 sky130_fd_sc_hd__buf_4 fanout851 (.A(net853),
    .X(net851));
 sky130_fd_sc_hd__buf_4 fanout852 (.A(net853),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_8 fanout853 (.A(net867),
    .X(net853));
 sky130_fd_sc_hd__buf_4 fanout854 (.A(net856),
    .X(net854));
 sky130_fd_sc_hd__buf_4 fanout855 (.A(net856),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_4 fanout856 (.A(net857),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_4 fanout857 (.A(net867),
    .X(net857));
 sky130_fd_sc_hd__buf_4 fanout858 (.A(net860),
    .X(net858));
 sky130_fd_sc_hd__clkbuf_2 fanout859 (.A(net860),
    .X(net859));
 sky130_fd_sc_hd__buf_4 fanout860 (.A(net861),
    .X(net860));
 sky130_fd_sc_hd__clkbuf_4 fanout861 (.A(net867),
    .X(net861));
 sky130_fd_sc_hd__buf_4 fanout862 (.A(net865),
    .X(net862));
 sky130_fd_sc_hd__buf_4 fanout863 (.A(net865),
    .X(net863));
 sky130_fd_sc_hd__clkbuf_2 fanout864 (.A(net865),
    .X(net864));
 sky130_fd_sc_hd__buf_4 fanout865 (.A(net867),
    .X(net865));
 sky130_fd_sc_hd__buf_6 fanout866 (.A(\u_dcg_peri.reset_n ),
    .X(net866));
 sky130_fd_sc_hd__buf_4 fanout868 (.A(net871),
    .X(net868));
 sky130_fd_sc_hd__clkbuf_2 fanout869 (.A(net871),
    .X(net869));
 sky130_fd_sc_hd__buf_4 fanout870 (.A(net871),
    .X(net870));
 sky130_fd_sc_hd__clkbuf_4 fanout871 (.A(net873),
    .X(net871));
 sky130_fd_sc_hd__buf_4 fanout872 (.A(net873),
    .X(net872));
 sky130_fd_sc_hd__buf_2 fanout873 (.A(net919),
    .X(net873));
 sky130_fd_sc_hd__clkbuf_4 fanout874 (.A(net877),
    .X(net874));
 sky130_fd_sc_hd__clkbuf_4 fanout875 (.A(net877),
    .X(net875));
 sky130_fd_sc_hd__clkbuf_4 fanout876 (.A(net877),
    .X(net876));
 sky130_fd_sc_hd__buf_2 fanout877 (.A(net878),
    .X(net877));
 sky130_fd_sc_hd__buf_4 fanout878 (.A(net919),
    .X(net878));
 sky130_fd_sc_hd__buf_4 fanout879 (.A(net880),
    .X(net879));
 sky130_fd_sc_hd__buf_4 fanout880 (.A(net919),
    .X(net880));
 sky130_fd_sc_hd__buf_4 fanout881 (.A(net884),
    .X(net881));
 sky130_fd_sc_hd__buf_2 fanout882 (.A(net884),
    .X(net882));
 sky130_fd_sc_hd__buf_4 fanout883 (.A(net884),
    .X(net883));
 sky130_fd_sc_hd__clkbuf_4 fanout884 (.A(net885),
    .X(net884));
 sky130_fd_sc_hd__clkbuf_4 fanout885 (.A(net893),
    .X(net885));
 sky130_fd_sc_hd__buf_4 fanout886 (.A(net889),
    .X(net886));
 sky130_fd_sc_hd__buf_2 fanout887 (.A(net889),
    .X(net887));
 sky130_fd_sc_hd__buf_4 fanout888 (.A(net889),
    .X(net888));
 sky130_fd_sc_hd__buf_2 fanout889 (.A(net893),
    .X(net889));
 sky130_fd_sc_hd__buf_4 fanout890 (.A(net893),
    .X(net890));
 sky130_fd_sc_hd__buf_6 fanout891 (.A(net893),
    .X(net891));
 sky130_fd_sc_hd__clkbuf_2 fanout892 (.A(net893),
    .X(net892));
 sky130_fd_sc_hd__buf_4 fanout893 (.A(net919),
    .X(net893));
 sky130_fd_sc_hd__clkbuf_4 fanout894 (.A(net896),
    .X(net894));
 sky130_fd_sc_hd__buf_4 fanout895 (.A(net896),
    .X(net895));
 sky130_fd_sc_hd__buf_2 fanout896 (.A(net897),
    .X(net896));
 sky130_fd_sc_hd__buf_2 fanout897 (.A(net918),
    .X(net897));
 sky130_fd_sc_hd__buf_4 fanout898 (.A(net901),
    .X(net898));
 sky130_fd_sc_hd__clkbuf_2 fanout899 (.A(net901),
    .X(net899));
 sky130_fd_sc_hd__buf_4 fanout900 (.A(net901),
    .X(net900));
 sky130_fd_sc_hd__buf_2 fanout901 (.A(net918),
    .X(net901));
 sky130_fd_sc_hd__buf_4 fanout902 (.A(net903),
    .X(net902));
 sky130_fd_sc_hd__clkbuf_4 fanout903 (.A(net905),
    .X(net903));
 sky130_fd_sc_hd__buf_4 fanout904 (.A(net905),
    .X(net904));
 sky130_fd_sc_hd__clkbuf_4 fanout905 (.A(net918),
    .X(net905));
 sky130_fd_sc_hd__clkbuf_4 fanout906 (.A(net908),
    .X(net906));
 sky130_fd_sc_hd__clkbuf_4 fanout907 (.A(net908),
    .X(net907));
 sky130_fd_sc_hd__buf_2 fanout908 (.A(net917),
    .X(net908));
 sky130_fd_sc_hd__buf_4 fanout909 (.A(net917),
    .X(net909));
 sky130_fd_sc_hd__buf_4 fanout910 (.A(net912),
    .X(net910));
 sky130_fd_sc_hd__buf_4 fanout911 (.A(net912),
    .X(net911));
 sky130_fd_sc_hd__clkbuf_4 fanout912 (.A(net914),
    .X(net912));
 sky130_fd_sc_hd__buf_4 fanout913 (.A(net914),
    .X(net913));
 sky130_fd_sc_hd__clkbuf_4 fanout914 (.A(net917),
    .X(net914));
 sky130_fd_sc_hd__clkbuf_8 fanout915 (.A(net917),
    .X(net915));
 sky130_fd_sc_hd__buf_2 fanout916 (.A(net917),
    .X(net916));
 sky130_fd_sc_hd__buf_4 fanout917 (.A(net918),
    .X(net917));
 sky130_fd_sc_hd__clkbuf_4 fanout918 (.A(net919),
    .X(net918));
 sky130_fd_sc_hd__buf_6 fanout919 (.A(net920),
    .X(net919));
 sky130_fd_sc_hd__buf_4 fanout921 (.A(net924),
    .X(net921));
 sky130_fd_sc_hd__buf_2 fanout922 (.A(net924),
    .X(net922));
 sky130_fd_sc_hd__buf_4 fanout923 (.A(net924),
    .X(net923));
 sky130_fd_sc_hd__buf_2 fanout924 (.A(_3594_),
    .X(net924));
 sky130_fd_sc_hd__buf_4 fanout925 (.A(net926),
    .X(net925));
 sky130_fd_sc_hd__buf_6 fanout926 (.A(_3594_),
    .X(net926));
 sky130_fd_sc_hd__buf_6 fanout927 (.A(net930),
    .X(net927));
 sky130_fd_sc_hd__buf_4 fanout928 (.A(net930),
    .X(net928));
 sky130_fd_sc_hd__buf_2 fanout929 (.A(net930),
    .X(net929));
 sky130_fd_sc_hd__buf_4 fanout930 (.A(_3594_),
    .X(net930));
 sky130_fd_sc_hd__buf_4 fanout931 (.A(net933),
    .X(net931));
 sky130_fd_sc_hd__buf_4 fanout932 (.A(net933),
    .X(net932));
 sky130_fd_sc_hd__buf_4 fanout933 (.A(_3593_),
    .X(net933));
 sky130_fd_sc_hd__clkbuf_8 fanout934 (.A(net936),
    .X(net934));
 sky130_fd_sc_hd__buf_4 fanout935 (.A(net936),
    .X(net935));
 sky130_fd_sc_hd__buf_6 fanout936 (.A(_3593_),
    .X(net936));
 sky130_fd_sc_hd__buf_4 fanout937 (.A(net940),
    .X(net937));
 sky130_fd_sc_hd__buf_2 fanout938 (.A(net940),
    .X(net938));
 sky130_fd_sc_hd__buf_4 fanout939 (.A(net940),
    .X(net939));
 sky130_fd_sc_hd__clkbuf_4 fanout940 (.A(_3421_),
    .X(net940));
 sky130_fd_sc_hd__buf_4 fanout941 (.A(net943),
    .X(net941));
 sky130_fd_sc_hd__buf_4 fanout942 (.A(net943),
    .X(net942));
 sky130_fd_sc_hd__buf_4 fanout943 (.A(_3421_),
    .X(net943));
 sky130_fd_sc_hd__buf_6 fanout944 (.A(net946),
    .X(net944));
 sky130_fd_sc_hd__buf_4 fanout945 (.A(net946),
    .X(net945));
 sky130_fd_sc_hd__clkbuf_8 fanout946 (.A(_3350_),
    .X(net946));
 sky130_fd_sc_hd__buf_6 fanout947 (.A(net950),
    .X(net947));
 sky130_fd_sc_hd__buf_4 fanout948 (.A(net950),
    .X(net948));
 sky130_fd_sc_hd__buf_2 fanout949 (.A(net950),
    .X(net949));
 sky130_fd_sc_hd__clkbuf_4 fanout950 (.A(_3350_),
    .X(net950));
 sky130_fd_sc_hd__clkbuf_8 fanout951 (.A(net954),
    .X(net951));
 sky130_fd_sc_hd__buf_4 fanout952 (.A(net954),
    .X(net952));
 sky130_fd_sc_hd__buf_4 fanout953 (.A(net954),
    .X(net953));
 sky130_fd_sc_hd__clkbuf_4 fanout954 (.A(net957),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_8 fanout955 (.A(net956),
    .X(net955));
 sky130_fd_sc_hd__buf_6 fanout956 (.A(net957),
    .X(net956));
 sky130_fd_sc_hd__buf_4 fanout957 (.A(_3349_),
    .X(net957));
 sky130_fd_sc_hd__buf_4 fanout958 (.A(net961),
    .X(net958));
 sky130_fd_sc_hd__buf_2 fanout959 (.A(net961),
    .X(net959));
 sky130_fd_sc_hd__buf_4 fanout960 (.A(net961),
    .X(net960));
 sky130_fd_sc_hd__buf_2 fanout961 (.A(net968),
    .X(net961));
 sky130_fd_sc_hd__buf_4 fanout962 (.A(net963),
    .X(net962));
 sky130_fd_sc_hd__buf_4 fanout963 (.A(net968),
    .X(net963));
 sky130_fd_sc_hd__buf_6 fanout964 (.A(net967),
    .X(net964));
 sky130_fd_sc_hd__buf_4 fanout965 (.A(net967),
    .X(net965));
 sky130_fd_sc_hd__buf_4 fanout966 (.A(net967),
    .X(net966));
 sky130_fd_sc_hd__buf_2 fanout967 (.A(net968),
    .X(net967));
 sky130_fd_sc_hd__buf_4 fanout968 (.A(_3348_),
    .X(net968));
 sky130_fd_sc_hd__clkbuf_8 fanout969 (.A(net972),
    .X(net969));
 sky130_fd_sc_hd__clkbuf_4 fanout970 (.A(net972),
    .X(net970));
 sky130_fd_sc_hd__buf_4 fanout971 (.A(net972),
    .X(net971));
 sky130_fd_sc_hd__clkbuf_4 fanout972 (.A(_3336_),
    .X(net972));
 sky130_fd_sc_hd__clkbuf_8 fanout973 (.A(net975),
    .X(net973));
 sky130_fd_sc_hd__buf_2 fanout974 (.A(net975),
    .X(net974));
 sky130_fd_sc_hd__buf_6 fanout975 (.A(_3336_),
    .X(net975));
 sky130_fd_sc_hd__clkbuf_4 fanout976 (.A(net977),
    .X(net976));
 sky130_fd_sc_hd__clkbuf_4 fanout977 (.A(_3266_),
    .X(net977));
 sky130_fd_sc_hd__buf_4 fanout978 (.A(_3265_),
    .X(net978));
 sky130_fd_sc_hd__buf_4 fanout979 (.A(net981),
    .X(net979));
 sky130_fd_sc_hd__buf_4 fanout980 (.A(net981),
    .X(net980));
 sky130_fd_sc_hd__clkbuf_4 fanout981 (.A(net988),
    .X(net981));
 sky130_fd_sc_hd__buf_4 fanout982 (.A(net983),
    .X(net982));
 sky130_fd_sc_hd__buf_4 fanout983 (.A(net988),
    .X(net983));
 sky130_fd_sc_hd__buf_4 fanout984 (.A(net985),
    .X(net984));
 sky130_fd_sc_hd__buf_2 fanout985 (.A(net988),
    .X(net985));
 sky130_fd_sc_hd__clkbuf_8 fanout986 (.A(net987),
    .X(net986));
 sky130_fd_sc_hd__buf_4 fanout987 (.A(net988),
    .X(net987));
 sky130_fd_sc_hd__buf_4 fanout988 (.A(_2945_),
    .X(net988));
 sky130_fd_sc_hd__buf_4 fanout989 (.A(net992),
    .X(net989));
 sky130_fd_sc_hd__buf_4 fanout990 (.A(net992),
    .X(net990));
 sky130_fd_sc_hd__clkbuf_4 fanout991 (.A(net992),
    .X(net991));
 sky130_fd_sc_hd__clkbuf_4 fanout992 (.A(_2934_),
    .X(net992));
 sky130_fd_sc_hd__buf_4 fanout993 (.A(net994),
    .X(net993));
 sky130_fd_sc_hd__buf_4 fanout994 (.A(net995),
    .X(net994));
 sky130_fd_sc_hd__buf_6 fanout995 (.A(_2934_),
    .X(net995));
 sky130_fd_sc_hd__buf_4 fanout996 (.A(_2921_),
    .X(net996));
 sky130_fd_sc_hd__buf_4 fanout997 (.A(net1799),
    .X(net997));
 sky130_fd_sc_hd__buf_4 fanout998 (.A(net999),
    .X(net998));
 sky130_fd_sc_hd__buf_4 fanout999 (.A(_2800_),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(s2_wbd_dat_i[10]),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(s1_wbd_dat_i[27]),
    .X(net1873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\u_s2.u_sync_wbb.u_resp_if.wr_ptr[0] ),
    .X(net1874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(s1_wbd_dat_i[24]),
    .X(net1875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(s1_wbd_dat_i[10]),
    .X(net1876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(s1_wbd_dat_i[19]),
    .X(net1877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\u_rst_sync.in_data_2s ),
    .X(net1878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(s0_wbd_dat_i[17]),
    .X(net1879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(s0_wbd_dat_i[6]),
    .X(net1880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(s0_wbd_dat_i[15]),
    .X(net1881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(s0_wbd_dat_i[2]),
    .X(net1882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net2089),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(m1_wbd_adr_i[2]),
    .X(net1883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_3223_),
    .X(net1884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_3224_),
    .X(net1885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(s0_wbd_dat_i[7]),
    .X(net1886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(m2_wbd_adr_i[5]),
    .X(net1887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_3233_),
    .X(net1888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(s0_wbd_dat_i[18]),
    .X(net1889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(s0_wbd_dat_i[4]),
    .X(net1890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(s0_wbd_dat_i[26]),
    .X(net1891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(s0_wbd_dat_i[9]),
    .X(net1892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\u_s2.u_sync_wbb.u_cmd_if.mem[3][61] ),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(s0_wbd_dat_i[24]),
    .X(net1893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(m0_wbd_adr_i[21]),
    .X(net1894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(m2_wbd_dat_i[28]),
    .X(net1895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_2764_),
    .X(net1896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(s0_wbd_dat_i[13]),
    .X(net1897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(s0_wbd_dat_i[10]),
    .X(net1898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(s0_wbd_dat_i[31]),
    .X(net1899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(m0_wbd_adr_i[28]),
    .X(net1900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_3116_),
    .X(net1901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(s0_wbd_dat_i[1]),
    .X(net1902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_2373_),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(s0_wbd_dat_i[3]),
    .X(net1903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(s0_wbd_dat_i[8]),
    .X(net1904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(s1_wbd_dat_i[12]),
    .X(net1905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(s1_wbd_dat_i[7]),
    .X(net1906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(s0_wbd_dat_i[25]),
    .X(net1907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(m0_wbd_adr_i[13]),
    .X(net1908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_3071_),
    .X(net1909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(s1_wbd_dat_i[9]),
    .X(net1910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(s1_wbd_dat_i[4]),
    .X(net1911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(s0_wbd_dat_i[21]),
    .X(net1912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0064_),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(s1_wbd_dat_i[0]),
    .X(net1913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(s1_wbd_dat_i[14]),
    .X(net1914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(m0_wbd_sel_i[1]),
    .X(net1915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(_3137_),
    .X(net1916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(m2_wbd_adr_i[4]),
    .X(net1917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_3229_),
    .X(net1918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_3230_),
    .X(net1919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(s1_wbd_dat_i[15]),
    .X(net1920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(s1_wbd_dat_i[16]),
    .X(net1921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\u_dcg_s0.u_dsync.in_data_2s[0] ),
    .X(net1922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\u_s2.u_sync_wbb.u_cmd_if.mem[2][60] ),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(s1_wbd_dat_i[18]),
    .X(net1923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(s1_wbd_dat_i[1]),
    .X(net1924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\u_s1.u_sync_wbb.m_state[0] ),
    .X(net1925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_0004_),
    .X(net1926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(s2_wbd_dat_i[24]),
    .X(net1927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(m2_wbd_dat_i[18]),
    .X(net1928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(s1_wbd_dat_i[2]),
    .X(net1929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(s2_wbd_dat_i[28]),
    .X(net1930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(m2_wbd_adr_i[3]),
    .X(net1931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_3226_),
    .X(net1932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_2372_),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_3227_),
    .X(net1933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(m2_wbd_dat_i[25]),
    .X(net1934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_3206_),
    .X(net1935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(s1_wbd_dat_i[5]),
    .X(net1936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(s2_wbd_dat_i[26]),
    .X(net1937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(s1_wbd_dat_i[8]),
    .X(net1938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(s2_wbd_dat_i[30]),
    .X(net1939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\u_dsync.in_data_2s[3] ),
    .X(net1940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(s2_wbd_dat_i[25]),
    .X(net1941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(s1_wbd_dat_i[6]),
    .X(net1942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(s2_wbd_dat_i[6]),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(s2_wbd_dat_i[31]),
    .X(net1943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\u_dsync.in_data_2s[4] ),
    .X(net1944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(m1_wbd_dat_i[27]),
    .X(net1945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(m0_wbd_adr_i[8]),
    .X(net1946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(m2_wbd_dat_i[11]),
    .X(net1947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(_2727_),
    .X(net1948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(m1_wbd_dat_i[17]),
    .X(net1949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(m2_wbd_dat_i[20]),
    .X(net1950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\u_s1.u_sync_wbb.u_cmd_if.mem[3][47] ),
    .X(net1951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\u_s1.u_sync_wbb.u_cmd_if.wr_ptr[0] ),
    .X(net1952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(s2_wbd_dat_i[12]),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(_2800_),
    .X(net1953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(m0_wbd_adr_i[9]),
    .X(net1954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(m2_wbd_dat_i[26]),
    .X(net1955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\u_dsync.in_data_s[7] ),
    .X(net1956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\u_s0.u_sync_wbb.u_cmd_if.mem[0][29] ),
    .X(net1957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(_2442_),
    .X(net1958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\u_dsync.in_data_s[5] ),
    .X(net1959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\u_dsync.in_data_s[3] ),
    .X(net1960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\u_dcg_s1.u_dsync.in_data_s[1] ),
    .X(net1961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\u_s1.u_sync_wbb.m_bl_cnt[3] ),
    .X(net1962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(s2_wbd_dat_i[18]),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\u_dcg_s1.u_dsync.in_data_2s[1] ),
    .X(net1963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(m2_wbd_dat_i[30]),
    .X(net1964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\u_dsync.in_data_2s[2] ),
    .X(net1965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\u_dsync.in_data_2s[6] ),
    .X(net1966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(m0_wbd_dat_i[7]),
    .X(net1967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(_3162_),
    .X(net1968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\u_dsync.in_data_s[1] ),
    .X(net1969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(m0_wbd_sel_i[3]),
    .X(net1970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\u_dcg_s0.u_dsync.in_data_s[1] ),
    .X(net1971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\u_dsync.in_data_s[6] ),
    .X(net1972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(s0_wbd_dat_i[12]),
    .X(net1980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\u_reg.reg_5[17] ),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(m2_wbd_dat_i[4]),
    .X(net1973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(m0_wbd_sel_i[2]),
    .X(net1974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\u_dsync.in_data_2s[0] ),
    .X(net1975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(m0_wbd_dat_i[19]),
    .X(net1976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\u_dcg_riscv.u_dsync.in_data_s[0] ),
    .X(net1977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(s0_wbd_dat_i[20]),
    .X(net1978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(s0_wbd_dat_i[28]),
    .X(net1979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(s0_wbd_dat_i[0]),
    .X(net1984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(m0_wbd_dat_i[30]),
    .X(net1985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(_2769_),
    .X(net1986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_3524_),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(s0_wbd_dat_i[14]),
    .X(net1987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(s0_wbd_dat_i[26]),
    .X(net1988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(s0_wbd_dat_i[23]),
    .X(net1989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(m0_wbd_adr_i[24]),
    .X(net1990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(m1_wbd_adr_i[23]),
    .X(net1991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_3100_),
    .X(net1992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(s0_wbd_dat_i[19]),
    .X(net1993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(m0_wbd_adr_i[29]),
    .X(net1994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(m1_wbd_adr_i[19]),
    .X(net1995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(s0_wbd_dat_i[11]),
    .X(net1996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(s2_wbd_dat_i[3]),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(m2_wbd_adr_i[14]),
    .X(net1997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_3074_),
    .X(net1998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(s0_wbd_dat_i[10]),
    .X(net1999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(m1_wbd_adr_i[21]),
    .X(net2000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_3094_),
    .X(net2001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(s0_wbd_dat_i[25]),
    .X(net2002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(s0_wbd_dat_i[13]),
    .X(net2003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(m1_wbd_adr_i[18]),
    .X(net2004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(_3085_),
    .X(net2005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(m1_wbd_dat_i[4]),
    .X(net2006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(s2_wbd_dat_i[5]),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_2969_),
    .X(net2007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(m1_wbd_dat_i[19]),
    .X(net2008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_3007_),
    .X(net2009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(m0_wbd_dat_i[27]),
    .X(net2010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(_2761_),
    .X(net2011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(m0_wbd_adr_i[25]),
    .X(net2012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(m2_wbd_dat_i[28]),
    .X(net2013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(_3214_),
    .X(net2014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(m0_wbd_adr_i[20]),
    .X(net2015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(m1_wbd_dat_i[24]),
    .X(net2016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(s2_wbd_dat_i[2]),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_3019_),
    .X(net2017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(m0_wbd_dat_i[26]),
    .X(net2018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(m2_wbd_dat_i[17]),
    .X(net2019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(_3188_),
    .X(net2020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(m0_wbd_adr_i[8]),
    .X(net2021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_3056_),
    .X(net2022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(m1_wbd_dat_i[29]),
    .X(net2023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(_2767_),
    .X(net2024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(m2_wbd_adr_i[8]),
    .X(net2025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(_3242_),
    .X(net2026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\u_s2.u_sync_wbb.m_state[2] ),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(m0_wbd_sel_i[3]),
    .X(net2027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(m0_wbd_dat_i[29]),
    .X(net2028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(_3216_),
    .X(net2029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(m0_wbd_sel_i[1]),
    .X(net2030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(m0_wbd_adr_i[9]),
    .X(net2031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(m1_wbd_adr_i[9]),
    .X(net2032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(s1_wbd_dat_i[22]),
    .X(net2033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(m0_wbd_adr_i[22]),
    .X(net2034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(m0_wbd_adr_i[6]),
    .X(net2035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(m2_wbd_dat_i[15]),
    .X(net2036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_2920_),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(m1_wbd_dat_i[25]),
    .X(net2037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(_3022_),
    .X(net2038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(m1_wbd_dat_i[16]),
    .X(net2039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(_2998_),
    .X(net2040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(m2_wbd_dat_i[27]),
    .X(net2041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(s1_wbd_dat_i[19]),
    .X(net2042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(m1_wbd_dat_i[27]),
    .X(net2043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(s1_wbd_dat_i[10]),
    .X(net2044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(s1_wbd_dat_i[24]),
    .X(net2045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(m0_wbd_sel_i[2]),
    .X(net2046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_1022_),
    .X(net1800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(s1_wbd_ack_i),
    .X(net2047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(s1_wbd_dat_i[26]),
    .X(net2048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(s0_wbd_ack_i),
    .X(net2049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(m2_wbd_dat_i[0]),
    .X(net2050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(m2_wbd_dat_i[22]),
    .X(net2051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(m1_wbd_dat_i[2]),
    .X(net2052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(_3150_),
    .X(net2053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(m2_wbd_dat_i[19]),
    .X(net2054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(m1_wbd_dat_i[12]),
    .X(net2055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(m2_wbd_dat_i[18]),
    .X(net2056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(s2_wbd_dat_i[15]),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(m0_wbd_dat_i[31]),
    .X(net2057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(_3035_),
    .X(net2058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(m1_wbd_sel_i[3]),
    .X(net2059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(s0_wbd_dat_i[2]),
    .X(net2060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(m2_wbd_dat_i[29]),
    .X(net2061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(m0_wbd_dat_i[4]),
    .X(net2062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(s0_wbd_dat_i[4]),
    .X(net2063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(m1_wbd_dat_i[20]),
    .X(net2064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(s0_wbd_dat_i[5]),
    .X(net2065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(m2_wbd_dat_i[13]),
    .X(net2066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(s2_wbd_dat_i[0]),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(m2_wbd_dat_i[26]),
    .X(net2067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(m1_wbd_dat_i[10]),
    .X(net2068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(_3170_),
    .X(net2069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(s2_wbd_dat_i[29]),
    .X(net2070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(m1_wbd_dat_i[30]),
    .X(net2071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(m2_wbd_dat_i[14]),
    .X(net2072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(_3179_),
    .X(net2073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(m2_wbd_adr_i[9]),
    .X(net2074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(m0_wbd_dat_i[20]),
    .X(net2075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(m2_wbd_dat_i[16]),
    .X(net2076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(m0_wbd_adr_i[27]),
    .X(net1981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\u_s2.u_sync_wbb.u_cmd_if.mem[2][7] ),
    .X(net1803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(m1_wbd_dat_i[8]),
    .X(net2077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(m2_wbd_dat_i[1]),
    .X(net2078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(m2_wbd_dat_i[25]),
    .X(net2079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(_2873_),
    .X(net2080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(s2_wbd_dat_i[7]),
    .X(net2081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(m2_wbd_sel_i[0]),
    .X(net2082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(_3134_),
    .X(net2083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(m1_wbd_dat_i[7]),
    .X(net2084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(m1_wbd_sel_i[0]),
    .X(net2085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(m1_wbd_adr_i[30]),
    .X(net2086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_2574_),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(m2_wbd_sel_i[3]),
    .X(net2087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(m2_wbd_dat_i[3]),
    .X(net2088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(s2_wbd_ack_i),
    .X(net2089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(m1_wbd_adr_i[26]),
    .X(net2090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(m1_wbd_dat_i[28]),
    .X(net2091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(m2_wbd_adr_i[5]),
    .X(net2092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(m0_wbd_adr_i[3]),
    .X(net2093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(s2_wbd_dat_i[1]),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(s2_wbd_dat_i[17]),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(s2_wbd_dat_i[22]),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(s2_wbd_dat_i[16]),
    .X(net1808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(s2_wbd_dat_i[19]),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(s2_wbd_dat_i[27]),
    .X(net1810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(s2_wbd_dat_i[14]),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(s2_wbd_dat_i[21]),
    .X(net1812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(s0_wbd_dat_i[27]),
    .X(net1982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(s2_wbd_dat_i[11]),
    .X(net1813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(s2_wbd_dat_i[13]),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\u_s2.u_sync_wbb.u_cmd_if.mem[0][5] ),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_2572_),
    .X(net1816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\u_s2.u_sync_wbb.m_state[1] ),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_2929_),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0483_),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\u_reg.cfg_dcg_ctrl[26] ),
    .X(net1820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_3558_),
    .X(net1821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_3561_),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(m1_wbd_adr_i[6]),
    .X(net1983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\u_dsync.in_data_2s[7] ),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\u_reg.cfg_dcg_ctrl[16] ),
    .X(net1824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_3520_),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\u_s2.u_sync_wbb.m_state[0] ),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_1972_),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(s2_wbd_dat_i[23]),
    .X(net1828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(s2_wbd_dat_i[20]),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(s2_wbd_dat_i[9]),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(s2_wbd_dat_i[8]),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(m0_wbd_adr_i[6]),
    .X(net1832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(s2_wbd_dat_i[4]),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_3236_),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(s0_wbd_dat_i[12]),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(s0_wbd_dat_i[20]),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(s0_wbd_dat_i[27]),
    .X(net1836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(s0_wbd_dat_i[28]),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(s0_wbd_dat_i[30]),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(m2_wbd_dat_i[24]),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_3204_),
    .X(net1840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(s0_wbd_dat_i[14]),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(m0_wbd_adr_i[23]),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(_0313_),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(m0_wbd_adr_i[19]),
    .X(net1843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(s0_wbd_dat_i[22]),
    .X(net1844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(s0_wbd_dat_i[29]),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(s0_wbd_dat_i[23]),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(m0_wbd_adr_i[26]),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_3110_),
    .X(net1848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\u_dcg_s0.u_dsync.in_data_2s[1] ),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(s1_wbd_dat_i[3]),
    .X(net1850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(s0_wbd_dat_i[16]),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(m0_wbd_adr_i[31]),
    .X(net1852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net1783),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_3125_),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(m0_wbd_adr_i[18]),
    .X(net1854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(m2_wbd_dat_i[2]),
    .X(net1855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(s1_wbd_dat_i[13]),
    .X(net1856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(s1_wbd_dat_i[20]),
    .X(net1857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(m0_wbd_adr_i[14]),
    .X(net1858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(s1_wbd_dat_i[29]),
    .X(net1859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(s1_wbd_dat_i[17]),
    .X(net1860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(s1_wbd_dat_i[28]),
    .X(net1861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(s1_wbd_dat_i[21]),
    .X(net1862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0351_),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(s1_wbd_dat_i[31]),
    .X(net1863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(s1_wbd_dat_i[11]),
    .X(net1864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(s1_wbd_dat_i[25]),
    .X(net1865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(m0_wbd_adr_i[30]),
    .X(net1866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_3122_),
    .X(net1867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(m0_wbd_adr_i[15]),
    .X(net1868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_3077_),
    .X(net1869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(s1_wbd_dat_i[23]),
    .X(net1870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(s1_wbd_dat_i[22]),
    .X(net1871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(s1_wbd_dat_i[30]),
    .X(net1872));
 sky130_fd_sc_hd__buf_4 max_length1036 (.A(_2152_),
    .X(net1036));
 sky130_fd_sc_hd__buf_4 max_length1050 (.A(_2134_),
    .X(net1050));
 sky130_fd_sc_hd__buf_6 max_length1097 (.A(_2081_),
    .X(net1097));
 sky130_fd_sc_hd__buf_4 max_length11 (.A(net1744),
    .X(net1743));
 sky130_fd_sc_hd__buf_6 max_length1101 (.A(_2076_),
    .X(net1101));
 sky130_fd_sc_hd__buf_4 max_length1119 (.A(_2056_),
    .X(net1119));
 sky130_fd_sc_hd__buf_6 max_length12 (.A(\clknet_3_0__leaf_u_dsync.out_clk ),
    .X(net1744));
 sky130_fd_sc_hd__buf_6 max_length14 (.A(\clknet_3_1__leaf_u_dsync.out_clk ),
    .X(net1746));
 sky130_fd_sc_hd__buf_4 max_length1403 (.A(\u_s2.u_sync_wbb.wbm_ack_o ),
    .X(net1403));
 sky130_fd_sc_hd__buf_6 max_length15 (.A(\clknet_3_2__leaf_u_dsync.out_clk ),
    .X(net1747));
 sky130_fd_sc_hd__buf_4 max_length1518 (.A(net1973),
    .X(net1518));
 sky130_fd_sc_hd__buf_4 max_length1521 (.A(m2_wbd_dat_i[29]),
    .X(net1521));
 sky130_fd_sc_hd__buf_4 max_length1530 (.A(m2_wbd_dat_i[15]),
    .X(net1530));
 sky130_fd_sc_hd__buf_6 max_length16 (.A(\clknet_3_2__leaf_u_dsync.out_clk ),
    .X(net1748));
 sky130_fd_sc_hd__buf_6 max_length17 (.A(\clknet_3_3__leaf_u_dsync.out_clk ),
    .X(net1749));
 sky130_fd_sc_hd__buf_6 max_length18 (.A(net1751),
    .X(net1750));
 sky130_fd_sc_hd__buf_6 max_length19 (.A(\clknet_3_3__leaf_u_dsync.out_clk ),
    .X(net1751));
 sky130_fd_sc_hd__buf_4 max_length20 (.A(\clknet_3_4__leaf_u_dsync.out_clk ),
    .X(net1752));
 sky130_fd_sc_hd__buf_6 max_length22 (.A(\clknet_3_4__leaf_u_dsync.out_clk ),
    .X(net1754));
 sky130_fd_sc_hd__buf_4 max_length26 (.A(\clknet_3_5__leaf_u_dsync.out_clk ),
    .X(net1758));
 sky130_fd_sc_hd__clkbuf_2 max_length37 (.A(clknet_2_1__leaf_mclk_raw),
    .X(net1769));
 sky130_fd_sc_hd__buf_6 max_length520 (.A(_3351_),
    .X(net520));
 sky130_fd_sc_hd__clkbuf_8 max_length554 (.A(_2746_),
    .X(net554));
 sky130_fd_sc_hd__clkbuf_4 max_length7 (.A(\clknet_1_0_0_u_dsync.out_clk ),
    .X(net1739));
 sky130_fd_sc_hd__buf_4 max_length704 (.A(_2690_),
    .X(net704));
 sky130_fd_sc_hd__buf_2 max_length9 (.A(\clknet_1_1_0_u_dsync.out_clk ),
    .X(net1741));
 sky130_fd_sc_hd__buf_2 output1 (.A(net1),
    .X(ch_clk_out[0]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(ch_data_out[105]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(ch_data_out[44]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(ch_data_out[45]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(ch_data_out[46]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(ch_data_out[47]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(ch_data_out[48]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(ch_data_out[49]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(ch_data_out[4]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(ch_data_out[50]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(ch_data_out[51]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(ch_data_out[52]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(ch_data_out[106]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(ch_data_out[53]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(ch_data_out[54]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(ch_data_out[55]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(ch_data_out[56]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(ch_data_out[57]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(ch_data_out[58]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(ch_data_out[59]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(ch_data_out[5]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(ch_data_out[60]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net119),
    .X(ch_data_out[61]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(ch_data_out[107]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(ch_data_out[62]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(ch_data_out[63]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(ch_data_out[64]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(ch_data_out[65]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(ch_data_out[66]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(ch_data_out[67]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(ch_data_out[68]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(ch_data_out[69]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(ch_data_out[6]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(ch_data_out[70]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(ch_data_out[108]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(ch_data_out[71]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(ch_data_out[72]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(ch_data_out[73]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net133),
    .X(ch_data_out[74]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(ch_data_out[75]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(ch_data_out[76]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net136),
    .X(ch_data_out[77]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net137),
    .X(ch_data_out[78]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net138),
    .X(ch_data_out[79]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(ch_data_out[7]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(ch_data_out[109]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net140),
    .X(ch_data_out[80]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net141),
    .X(ch_data_out[81]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net142),
    .X(ch_data_out[82]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net143),
    .X(ch_data_out[83]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net144),
    .X(ch_data_out[84]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net145),
    .X(ch_data_out[85]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net146),
    .X(ch_data_out[86]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net147),
    .X(ch_data_out[87]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net148),
    .X(ch_data_out[88]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net149),
    .X(ch_data_out[89]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(ch_data_out[10]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net150),
    .X(ch_data_out[8]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net151),
    .X(ch_data_out[90]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net152),
    .X(ch_data_out[91]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net153),
    .X(ch_data_out[92]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net154),
    .X(ch_data_out[93]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net155),
    .X(ch_data_out[94]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net156),
    .X(ch_data_out[95]));
 sky130_fd_sc_hd__buf_2 output157 (.A(net157),
    .X(ch_data_out[96]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net158),
    .X(ch_data_out[97]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(ch_data_out[98]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(ch_data_out[110]));
 sky130_fd_sc_hd__buf_2 output160 (.A(net160),
    .X(ch_data_out[99]));
 sky130_fd_sc_hd__buf_2 output161 (.A(net161),
    .X(ch_data_out[9]));
 sky130_fd_sc_hd__buf_4 output162 (.A(net162),
    .X(m0_wbd_ack_o));
 sky130_fd_sc_hd__buf_6 output163 (.A(net163),
    .X(m0_wbd_dat_o[0]));
 sky130_fd_sc_hd__buf_6 output164 (.A(net164),
    .X(m0_wbd_dat_o[10]));
 sky130_fd_sc_hd__buf_4 output165 (.A(net165),
    .X(m0_wbd_dat_o[11]));
 sky130_fd_sc_hd__buf_6 output166 (.A(net166),
    .X(m0_wbd_dat_o[12]));
 sky130_fd_sc_hd__buf_4 output167 (.A(net167),
    .X(m0_wbd_dat_o[13]));
 sky130_fd_sc_hd__buf_2 output168 (.A(net168),
    .X(m0_wbd_dat_o[14]));
 sky130_fd_sc_hd__buf_4 output169 (.A(net169),
    .X(m0_wbd_dat_o[15]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(ch_data_out[111]));
 sky130_fd_sc_hd__buf_6 output170 (.A(net170),
    .X(m0_wbd_dat_o[16]));
 sky130_fd_sc_hd__buf_4 output171 (.A(net171),
    .X(m0_wbd_dat_o[17]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net172),
    .X(m0_wbd_dat_o[18]));
 sky130_fd_sc_hd__buf_4 output173 (.A(net173),
    .X(m0_wbd_dat_o[19]));
 sky130_fd_sc_hd__buf_4 output174 (.A(net174),
    .X(m0_wbd_dat_o[1]));
 sky130_fd_sc_hd__buf_6 output175 (.A(net175),
    .X(m0_wbd_dat_o[20]));
 sky130_fd_sc_hd__buf_4 output176 (.A(net176),
    .X(m0_wbd_dat_o[21]));
 sky130_fd_sc_hd__buf_2 output177 (.A(net177),
    .X(m0_wbd_dat_o[22]));
 sky130_fd_sc_hd__buf_6 output178 (.A(net178),
    .X(m0_wbd_dat_o[23]));
 sky130_fd_sc_hd__buf_4 output179 (.A(net179),
    .X(m0_wbd_dat_o[24]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net1489),
    .X(ch_data_out[112]));
 sky130_fd_sc_hd__buf_4 output180 (.A(net180),
    .X(m0_wbd_dat_o[25]));
 sky130_fd_sc_hd__buf_6 output181 (.A(net181),
    .X(m0_wbd_dat_o[26]));
 sky130_fd_sc_hd__buf_6 output182 (.A(net182),
    .X(m0_wbd_dat_o[27]));
 sky130_fd_sc_hd__buf_6 output183 (.A(net183),
    .X(m0_wbd_dat_o[28]));
 sky130_fd_sc_hd__buf_6 output184 (.A(net184),
    .X(m0_wbd_dat_o[29]));
 sky130_fd_sc_hd__buf_6 output185 (.A(net185),
    .X(m0_wbd_dat_o[2]));
 sky130_fd_sc_hd__buf_6 output186 (.A(net186),
    .X(m0_wbd_dat_o[30]));
 sky130_fd_sc_hd__buf_6 output187 (.A(net187),
    .X(m0_wbd_dat_o[31]));
 sky130_fd_sc_hd__buf_4 output188 (.A(net188),
    .X(m0_wbd_dat_o[3]));
 sky130_fd_sc_hd__buf_4 output189 (.A(net189),
    .X(m0_wbd_dat_o[4]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net1487),
    .X(ch_data_out[113]));
 sky130_fd_sc_hd__buf_4 output190 (.A(net190),
    .X(m0_wbd_dat_o[5]));
 sky130_fd_sc_hd__buf_4 output191 (.A(net191),
    .X(m0_wbd_dat_o[6]));
 sky130_fd_sc_hd__buf_4 output192 (.A(net192),
    .X(m0_wbd_dat_o[7]));
 sky130_fd_sc_hd__buf_4 output193 (.A(net193),
    .X(m0_wbd_dat_o[8]));
 sky130_fd_sc_hd__buf_6 output194 (.A(net194),
    .X(m0_wbd_dat_o[9]));
 sky130_fd_sc_hd__buf_2 output195 (.A(net195),
    .X(m0_wbd_lack_o));
 sky130_fd_sc_hd__buf_2 output196 (.A(net196),
    .X(m1_wbd_ack_o));
 sky130_fd_sc_hd__buf_2 output197 (.A(net197),
    .X(m1_wbd_dat_o[0]));
 sky130_fd_sc_hd__buf_2 output198 (.A(net198),
    .X(m1_wbd_dat_o[10]));
 sky130_fd_sc_hd__buf_2 output199 (.A(net199),
    .X(m1_wbd_dat_o[11]));
 sky130_fd_sc_hd__buf_2 output2 (.A(net2),
    .X(ch_clk_out[1]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net1485),
    .X(ch_data_out[114]));
 sky130_fd_sc_hd__buf_2 output200 (.A(net200),
    .X(m1_wbd_dat_o[12]));
 sky130_fd_sc_hd__buf_2 output201 (.A(net201),
    .X(m1_wbd_dat_o[13]));
 sky130_fd_sc_hd__buf_2 output202 (.A(net202),
    .X(m1_wbd_dat_o[14]));
 sky130_fd_sc_hd__buf_2 output203 (.A(net203),
    .X(m1_wbd_dat_o[15]));
 sky130_fd_sc_hd__buf_2 output204 (.A(net204),
    .X(m1_wbd_dat_o[16]));
 sky130_fd_sc_hd__buf_2 output205 (.A(net205),
    .X(m1_wbd_dat_o[17]));
 sky130_fd_sc_hd__buf_2 output206 (.A(net206),
    .X(m1_wbd_dat_o[18]));
 sky130_fd_sc_hd__clkbuf_4 output207 (.A(net207),
    .X(m1_wbd_dat_o[19]));
 sky130_fd_sc_hd__buf_2 output208 (.A(net208),
    .X(m1_wbd_dat_o[1]));
 sky130_fd_sc_hd__buf_2 output209 (.A(net209),
    .X(m1_wbd_dat_o[20]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net1483),
    .X(ch_data_out[115]));
 sky130_fd_sc_hd__buf_2 output210 (.A(net210),
    .X(m1_wbd_dat_o[21]));
 sky130_fd_sc_hd__buf_2 output211 (.A(net211),
    .X(m1_wbd_dat_o[22]));
 sky130_fd_sc_hd__buf_2 output212 (.A(net212),
    .X(m1_wbd_dat_o[23]));
 sky130_fd_sc_hd__buf_2 output213 (.A(net213),
    .X(m1_wbd_dat_o[24]));
 sky130_fd_sc_hd__buf_2 output214 (.A(net214),
    .X(m1_wbd_dat_o[25]));
 sky130_fd_sc_hd__buf_2 output215 (.A(net215),
    .X(m1_wbd_dat_o[26]));
 sky130_fd_sc_hd__buf_2 output216 (.A(net216),
    .X(m1_wbd_dat_o[27]));
 sky130_fd_sc_hd__buf_2 output217 (.A(net217),
    .X(m1_wbd_dat_o[28]));
 sky130_fd_sc_hd__buf_2 output218 (.A(net218),
    .X(m1_wbd_dat_o[29]));
 sky130_fd_sc_hd__buf_2 output219 (.A(net219),
    .X(m1_wbd_dat_o[2]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net1481),
    .X(ch_data_out[116]));
 sky130_fd_sc_hd__buf_2 output220 (.A(net220),
    .X(m1_wbd_dat_o[30]));
 sky130_fd_sc_hd__buf_2 output221 (.A(net221),
    .X(m1_wbd_dat_o[31]));
 sky130_fd_sc_hd__buf_2 output222 (.A(net222),
    .X(m1_wbd_dat_o[3]));
 sky130_fd_sc_hd__buf_2 output223 (.A(net223),
    .X(m1_wbd_dat_o[4]));
 sky130_fd_sc_hd__buf_2 output224 (.A(net224),
    .X(m1_wbd_dat_o[5]));
 sky130_fd_sc_hd__buf_2 output225 (.A(net225),
    .X(m1_wbd_dat_o[6]));
 sky130_fd_sc_hd__buf_2 output226 (.A(net226),
    .X(m1_wbd_dat_o[7]));
 sky130_fd_sc_hd__buf_2 output227 (.A(net227),
    .X(m1_wbd_dat_o[8]));
 sky130_fd_sc_hd__buf_2 output228 (.A(net228),
    .X(m1_wbd_dat_o[9]));
 sky130_fd_sc_hd__buf_2 output229 (.A(net229),
    .X(m1_wbd_lack_o));
 sky130_fd_sc_hd__buf_2 output23 (.A(net1479),
    .X(ch_data_out[117]));
 sky130_fd_sc_hd__buf_2 output230 (.A(net230),
    .X(m2_wbd_ack_o));
 sky130_fd_sc_hd__buf_2 output231 (.A(net231),
    .X(m2_wbd_dat_o[0]));
 sky130_fd_sc_hd__buf_2 output232 (.A(net232),
    .X(m2_wbd_dat_o[10]));
 sky130_fd_sc_hd__buf_2 output233 (.A(net233),
    .X(m2_wbd_dat_o[11]));
 sky130_fd_sc_hd__buf_2 output234 (.A(net234),
    .X(m2_wbd_dat_o[12]));
 sky130_fd_sc_hd__buf_2 output235 (.A(net235),
    .X(m2_wbd_dat_o[13]));
 sky130_fd_sc_hd__buf_2 output236 (.A(net236),
    .X(m2_wbd_dat_o[14]));
 sky130_fd_sc_hd__buf_2 output237 (.A(net237),
    .X(m2_wbd_dat_o[15]));
 sky130_fd_sc_hd__buf_2 output238 (.A(net238),
    .X(m2_wbd_dat_o[16]));
 sky130_fd_sc_hd__buf_2 output239 (.A(net239),
    .X(m2_wbd_dat_o[17]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net1477),
    .X(ch_data_out[118]));
 sky130_fd_sc_hd__buf_2 output240 (.A(net240),
    .X(m2_wbd_dat_o[18]));
 sky130_fd_sc_hd__buf_2 output241 (.A(net241),
    .X(m2_wbd_dat_o[19]));
 sky130_fd_sc_hd__buf_2 output242 (.A(net242),
    .X(m2_wbd_dat_o[1]));
 sky130_fd_sc_hd__buf_2 output243 (.A(net243),
    .X(m2_wbd_dat_o[20]));
 sky130_fd_sc_hd__buf_2 output244 (.A(net244),
    .X(m2_wbd_dat_o[21]));
 sky130_fd_sc_hd__buf_2 output245 (.A(net245),
    .X(m2_wbd_dat_o[22]));
 sky130_fd_sc_hd__buf_2 output246 (.A(net246),
    .X(m2_wbd_dat_o[23]));
 sky130_fd_sc_hd__buf_2 output247 (.A(net247),
    .X(m2_wbd_dat_o[24]));
 sky130_fd_sc_hd__buf_2 output248 (.A(net248),
    .X(m2_wbd_dat_o[25]));
 sky130_fd_sc_hd__buf_2 output249 (.A(net249),
    .X(m2_wbd_dat_o[26]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net1475),
    .X(ch_data_out[119]));
 sky130_fd_sc_hd__buf_2 output250 (.A(net250),
    .X(m2_wbd_dat_o[27]));
 sky130_fd_sc_hd__buf_2 output251 (.A(net251),
    .X(m2_wbd_dat_o[28]));
 sky130_fd_sc_hd__buf_2 output252 (.A(net252),
    .X(m2_wbd_dat_o[29]));
 sky130_fd_sc_hd__buf_2 output253 (.A(net253),
    .X(m2_wbd_dat_o[2]));
 sky130_fd_sc_hd__buf_2 output254 (.A(net254),
    .X(m2_wbd_dat_o[30]));
 sky130_fd_sc_hd__buf_2 output255 (.A(net255),
    .X(m2_wbd_dat_o[31]));
 sky130_fd_sc_hd__buf_2 output256 (.A(net256),
    .X(m2_wbd_dat_o[3]));
 sky130_fd_sc_hd__buf_4 output257 (.A(net257),
    .X(m2_wbd_dat_o[4]));
 sky130_fd_sc_hd__buf_2 output258 (.A(net258),
    .X(m2_wbd_dat_o[5]));
 sky130_fd_sc_hd__buf_2 output259 (.A(net259),
    .X(m2_wbd_dat_o[6]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net1491),
    .X(ch_data_out[11]));
 sky130_fd_sc_hd__buf_2 output260 (.A(net260),
    .X(m2_wbd_dat_o[7]));
 sky130_fd_sc_hd__buf_4 output261 (.A(net261),
    .X(m2_wbd_dat_o[8]));
 sky130_fd_sc_hd__buf_2 output262 (.A(net262),
    .X(m2_wbd_dat_o[9]));
 sky130_fd_sc_hd__buf_2 output263 (.A(net263),
    .X(m2_wbd_lack_o));
 sky130_fd_sc_hd__buf_2 output264 (.A(net264),
    .X(m3_wbd_ack_o));
 sky130_fd_sc_hd__buf_2 output265 (.A(net265),
    .X(m3_wbd_dat_o[0]));
 sky130_fd_sc_hd__buf_2 output266 (.A(net266),
    .X(m3_wbd_dat_o[10]));
 sky130_fd_sc_hd__buf_2 output267 (.A(net267),
    .X(m3_wbd_dat_o[11]));
 sky130_fd_sc_hd__buf_2 output268 (.A(net268),
    .X(m3_wbd_dat_o[12]));
 sky130_fd_sc_hd__buf_2 output269 (.A(net269),
    .X(m3_wbd_dat_o[13]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net1473),
    .X(ch_data_out[120]));
 sky130_fd_sc_hd__buf_2 output270 (.A(net270),
    .X(m3_wbd_dat_o[14]));
 sky130_fd_sc_hd__buf_2 output271 (.A(net271),
    .X(m3_wbd_dat_o[15]));
 sky130_fd_sc_hd__buf_2 output272 (.A(net272),
    .X(m3_wbd_dat_o[16]));
 sky130_fd_sc_hd__buf_2 output273 (.A(net273),
    .X(m3_wbd_dat_o[17]));
 sky130_fd_sc_hd__buf_2 output274 (.A(net274),
    .X(m3_wbd_dat_o[18]));
 sky130_fd_sc_hd__buf_2 output275 (.A(net275),
    .X(m3_wbd_dat_o[19]));
 sky130_fd_sc_hd__buf_2 output276 (.A(net276),
    .X(m3_wbd_dat_o[1]));
 sky130_fd_sc_hd__buf_2 output277 (.A(net277),
    .X(m3_wbd_dat_o[20]));
 sky130_fd_sc_hd__buf_2 output278 (.A(net278),
    .X(m3_wbd_dat_o[21]));
 sky130_fd_sc_hd__buf_2 output279 (.A(net279),
    .X(m3_wbd_dat_o[22]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net1471),
    .X(ch_data_out[121]));
 sky130_fd_sc_hd__buf_2 output280 (.A(net280),
    .X(m3_wbd_dat_o[23]));
 sky130_fd_sc_hd__buf_2 output281 (.A(net281),
    .X(m3_wbd_dat_o[24]));
 sky130_fd_sc_hd__buf_2 output282 (.A(net282),
    .X(m3_wbd_dat_o[25]));
 sky130_fd_sc_hd__buf_2 output283 (.A(net283),
    .X(m3_wbd_dat_o[26]));
 sky130_fd_sc_hd__buf_2 output284 (.A(net284),
    .X(m3_wbd_dat_o[27]));
 sky130_fd_sc_hd__buf_2 output285 (.A(net285),
    .X(m3_wbd_dat_o[28]));
 sky130_fd_sc_hd__buf_2 output286 (.A(net286),
    .X(m3_wbd_dat_o[29]));
 sky130_fd_sc_hd__buf_2 output287 (.A(net287),
    .X(m3_wbd_dat_o[2]));
 sky130_fd_sc_hd__buf_2 output288 (.A(net288),
    .X(m3_wbd_dat_o[30]));
 sky130_fd_sc_hd__buf_2 output289 (.A(net289),
    .X(m3_wbd_dat_o[31]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net1469),
    .X(ch_data_out[122]));
 sky130_fd_sc_hd__buf_2 output290 (.A(net290),
    .X(m3_wbd_dat_o[3]));
 sky130_fd_sc_hd__buf_2 output291 (.A(net291),
    .X(m3_wbd_dat_o[4]));
 sky130_fd_sc_hd__buf_2 output292 (.A(net292),
    .X(m3_wbd_dat_o[5]));
 sky130_fd_sc_hd__buf_2 output293 (.A(net293),
    .X(m3_wbd_dat_o[6]));
 sky130_fd_sc_hd__buf_2 output294 (.A(net294),
    .X(m3_wbd_dat_o[7]));
 sky130_fd_sc_hd__buf_2 output295 (.A(net295),
    .X(m3_wbd_dat_o[8]));
 sky130_fd_sc_hd__buf_2 output296 (.A(net296),
    .X(m3_wbd_dat_o[9]));
 sky130_fd_sc_hd__buf_2 output297 (.A(net297),
    .X(m3_wbd_lack_o));
 sky130_fd_sc_hd__clkbuf_1 output298 (.A(net298),
    .X(peri_wbclk));
 sky130_fd_sc_hd__clkbuf_1 output299 (.A(net299),
    .X(riscv_wbclk));
 sky130_fd_sc_hd__buf_2 output3 (.A(net3),
    .X(ch_clk_out[2]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net1467),
    .X(ch_data_out[123]));
 sky130_fd_sc_hd__clkbuf_1 output300 (.A(net300),
    .X(s0_mclk));
 sky130_fd_sc_hd__buf_2 output301 (.A(net301),
    .X(s0_wbd_adr_o[10]));
 sky130_fd_sc_hd__buf_2 output302 (.A(net302),
    .X(s0_wbd_adr_o[11]));
 sky130_fd_sc_hd__buf_2 output303 (.A(net303),
    .X(s0_wbd_adr_o[12]));
 sky130_fd_sc_hd__buf_2 output304 (.A(net304),
    .X(s0_wbd_adr_o[13]));
 sky130_fd_sc_hd__buf_2 output305 (.A(net305),
    .X(s0_wbd_adr_o[14]));
 sky130_fd_sc_hd__buf_2 output306 (.A(net306),
    .X(s0_wbd_adr_o[15]));
 sky130_fd_sc_hd__buf_2 output307 (.A(net307),
    .X(s0_wbd_adr_o[16]));
 sky130_fd_sc_hd__buf_2 output308 (.A(net308),
    .X(s0_wbd_adr_o[17]));
 sky130_fd_sc_hd__buf_2 output309 (.A(net309),
    .X(s0_wbd_adr_o[18]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net1465),
    .X(ch_data_out[124]));
 sky130_fd_sc_hd__buf_2 output310 (.A(net310),
    .X(s0_wbd_adr_o[19]));
 sky130_fd_sc_hd__buf_2 output311 (.A(net311),
    .X(s0_wbd_adr_o[20]));
 sky130_fd_sc_hd__buf_2 output312 (.A(net312),
    .X(s0_wbd_adr_o[21]));
 sky130_fd_sc_hd__buf_2 output313 (.A(net313),
    .X(s0_wbd_adr_o[22]));
 sky130_fd_sc_hd__buf_2 output314 (.A(net314),
    .X(s0_wbd_adr_o[23]));
 sky130_fd_sc_hd__buf_2 output315 (.A(net315),
    .X(s0_wbd_adr_o[24]));
 sky130_fd_sc_hd__buf_2 output316 (.A(net316),
    .X(s0_wbd_adr_o[25]));
 sky130_fd_sc_hd__buf_2 output317 (.A(net317),
    .X(s0_wbd_adr_o[26]));
 sky130_fd_sc_hd__buf_2 output318 (.A(net318),
    .X(s0_wbd_adr_o[27]));
 sky130_fd_sc_hd__buf_2 output319 (.A(net319),
    .X(s0_wbd_adr_o[28]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net1463),
    .X(ch_data_out[125]));
 sky130_fd_sc_hd__buf_2 output320 (.A(net320),
    .X(s0_wbd_adr_o[29]));
 sky130_fd_sc_hd__buf_2 output321 (.A(net321),
    .X(s0_wbd_adr_o[2]));
 sky130_fd_sc_hd__buf_2 output322 (.A(net322),
    .X(s0_wbd_adr_o[30]));
 sky130_fd_sc_hd__buf_2 output323 (.A(net323),
    .X(s0_wbd_adr_o[31]));
 sky130_fd_sc_hd__buf_2 output324 (.A(net324),
    .X(s0_wbd_adr_o[3]));
 sky130_fd_sc_hd__buf_2 output325 (.A(net325),
    .X(s0_wbd_adr_o[4]));
 sky130_fd_sc_hd__buf_2 output326 (.A(net326),
    .X(s0_wbd_adr_o[5]));
 sky130_fd_sc_hd__buf_2 output327 (.A(net327),
    .X(s0_wbd_adr_o[6]));
 sky130_fd_sc_hd__buf_2 output328 (.A(net328),
    .X(s0_wbd_adr_o[7]));
 sky130_fd_sc_hd__buf_2 output329 (.A(net329),
    .X(s0_wbd_adr_o[8]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net1461),
    .X(ch_data_out[126]));
 sky130_fd_sc_hd__buf_2 output330 (.A(net330),
    .X(s0_wbd_adr_o[9]));
 sky130_fd_sc_hd__buf_2 output331 (.A(net331),
    .X(s0_wbd_bl_o[0]));
 sky130_fd_sc_hd__buf_2 output332 (.A(net332),
    .X(s0_wbd_bl_o[1]));
 sky130_fd_sc_hd__buf_2 output333 (.A(net333),
    .X(s0_wbd_bl_o[2]));
 sky130_fd_sc_hd__buf_2 output334 (.A(net727),
    .X(s0_wbd_bl_o[3]));
 sky130_fd_sc_hd__buf_2 output335 (.A(net335),
    .X(s0_wbd_bl_o[4]));
 sky130_fd_sc_hd__buf_2 output336 (.A(net728),
    .X(s0_wbd_bl_o[5]));
 sky130_fd_sc_hd__buf_2 output337 (.A(net729),
    .X(s0_wbd_bl_o[6]));
 sky130_fd_sc_hd__buf_2 output338 (.A(net730),
    .X(s0_wbd_bl_o[7]));
 sky130_fd_sc_hd__buf_2 output339 (.A(net731),
    .X(s0_wbd_bl_o[8]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net1459),
    .X(ch_data_out[127]));
 sky130_fd_sc_hd__buf_2 output340 (.A(net340),
    .X(s0_wbd_bl_o[9]));
 sky130_fd_sc_hd__buf_2 output341 (.A(net341),
    .X(s0_wbd_bry_o));
 sky130_fd_sc_hd__buf_2 output342 (.A(net342),
    .X(s0_wbd_cyc_o));
 sky130_fd_sc_hd__buf_2 output343 (.A(net343),
    .X(s0_wbd_dat_o[0]));
 sky130_fd_sc_hd__buf_2 output344 (.A(net344),
    .X(s0_wbd_dat_o[10]));
 sky130_fd_sc_hd__buf_2 output345 (.A(net710),
    .X(s0_wbd_dat_o[11]));
 sky130_fd_sc_hd__buf_2 output346 (.A(net346),
    .X(s0_wbd_dat_o[12]));
 sky130_fd_sc_hd__buf_2 output347 (.A(net347),
    .X(s0_wbd_dat_o[13]));
 sky130_fd_sc_hd__buf_2 output348 (.A(net709),
    .X(s0_wbd_dat_o[14]));
 sky130_fd_sc_hd__buf_2 output349 (.A(net349),
    .X(s0_wbd_dat_o[15]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net1457),
    .X(ch_data_out[128]));
 sky130_fd_sc_hd__buf_2 output350 (.A(net350),
    .X(s0_wbd_dat_o[16]));
 sky130_fd_sc_hd__buf_2 output351 (.A(net351),
    .X(s0_wbd_dat_o[17]));
 sky130_fd_sc_hd__buf_2 output352 (.A(net352),
    .X(s0_wbd_dat_o[18]));
 sky130_fd_sc_hd__buf_2 output353 (.A(net353),
    .X(s0_wbd_dat_o[19]));
 sky130_fd_sc_hd__buf_2 output354 (.A(net354),
    .X(s0_wbd_dat_o[1]));
 sky130_fd_sc_hd__buf_2 output355 (.A(net355),
    .X(s0_wbd_dat_o[20]));
 sky130_fd_sc_hd__buf_2 output356 (.A(net356),
    .X(s0_wbd_dat_o[21]));
 sky130_fd_sc_hd__buf_2 output357 (.A(net357),
    .X(s0_wbd_dat_o[22]));
 sky130_fd_sc_hd__buf_2 output358 (.A(net358),
    .X(s0_wbd_dat_o[23]));
 sky130_fd_sc_hd__buf_2 output359 (.A(net359),
    .X(s0_wbd_dat_o[24]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net1455),
    .X(ch_data_out[129]));
 sky130_fd_sc_hd__buf_2 output360 (.A(net360),
    .X(s0_wbd_dat_o[25]));
 sky130_fd_sc_hd__buf_2 output361 (.A(net361),
    .X(s0_wbd_dat_o[26]));
 sky130_fd_sc_hd__buf_2 output362 (.A(net362),
    .X(s0_wbd_dat_o[27]));
 sky130_fd_sc_hd__buf_2 output363 (.A(net363),
    .X(s0_wbd_dat_o[28]));
 sky130_fd_sc_hd__buf_2 output364 (.A(net364),
    .X(s0_wbd_dat_o[29]));
 sky130_fd_sc_hd__buf_2 output365 (.A(net365),
    .X(s0_wbd_dat_o[2]));
 sky130_fd_sc_hd__buf_2 output366 (.A(net366),
    .X(s0_wbd_dat_o[30]));
 sky130_fd_sc_hd__buf_2 output367 (.A(net367),
    .X(s0_wbd_dat_o[31]));
 sky130_fd_sc_hd__buf_2 output368 (.A(net368),
    .X(s0_wbd_dat_o[3]));
 sky130_fd_sc_hd__buf_2 output369 (.A(net369),
    .X(s0_wbd_dat_o[4]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(ch_data_out[12]));
 sky130_fd_sc_hd__buf_2 output370 (.A(net370),
    .X(s0_wbd_dat_o[5]));
 sky130_fd_sc_hd__buf_2 output371 (.A(net371),
    .X(s0_wbd_dat_o[6]));
 sky130_fd_sc_hd__buf_2 output372 (.A(net372),
    .X(s0_wbd_dat_o[7]));
 sky130_fd_sc_hd__buf_2 output373 (.A(net373),
    .X(s0_wbd_dat_o[8]));
 sky130_fd_sc_hd__buf_2 output374 (.A(net374),
    .X(s0_wbd_dat_o[9]));
 sky130_fd_sc_hd__buf_2 output375 (.A(net375),
    .X(s0_wbd_sel_o[0]));
 sky130_fd_sc_hd__buf_2 output376 (.A(net376),
    .X(s0_wbd_sel_o[1]));
 sky130_fd_sc_hd__buf_2 output377 (.A(net377),
    .X(s0_wbd_sel_o[2]));
 sky130_fd_sc_hd__buf_2 output378 (.A(net378),
    .X(s0_wbd_sel_o[3]));
 sky130_fd_sc_hd__buf_2 output379 (.A(net379),
    .X(s0_wbd_stb_o));
 sky130_fd_sc_hd__buf_2 output38 (.A(net1453),
    .X(ch_data_out[130]));
 sky130_fd_sc_hd__buf_2 output380 (.A(net712),
    .X(s0_wbd_we_o));
 sky130_fd_sc_hd__clkbuf_1 output381 (.A(net381),
    .X(s1_mclk));
 sky130_fd_sc_hd__buf_2 output382 (.A(net382),
    .X(s1_wbd_adr_o[2]));
 sky130_fd_sc_hd__buf_2 output383 (.A(net383),
    .X(s1_wbd_adr_o[3]));
 sky130_fd_sc_hd__buf_2 output384 (.A(net384),
    .X(s1_wbd_adr_o[4]));
 sky130_fd_sc_hd__buf_2 output385 (.A(net385),
    .X(s1_wbd_adr_o[5]));
 sky130_fd_sc_hd__buf_2 output386 (.A(net386),
    .X(s1_wbd_adr_o[6]));
 sky130_fd_sc_hd__buf_2 output387 (.A(net387),
    .X(s1_wbd_adr_o[7]));
 sky130_fd_sc_hd__buf_2 output388 (.A(net388),
    .X(s1_wbd_adr_o[8]));
 sky130_fd_sc_hd__buf_2 output389 (.A(net389),
    .X(s1_wbd_cyc_o));
 sky130_fd_sc_hd__buf_2 output39 (.A(net1451),
    .X(ch_data_out[131]));
 sky130_fd_sc_hd__buf_2 output390 (.A(net390),
    .X(s1_wbd_dat_o[0]));
 sky130_fd_sc_hd__buf_2 output391 (.A(net391),
    .X(s1_wbd_dat_o[10]));
 sky130_fd_sc_hd__buf_2 output392 (.A(net392),
    .X(s1_wbd_dat_o[11]));
 sky130_fd_sc_hd__buf_2 output393 (.A(net393),
    .X(s1_wbd_dat_o[12]));
 sky130_fd_sc_hd__buf_2 output394 (.A(net394),
    .X(s1_wbd_dat_o[13]));
 sky130_fd_sc_hd__buf_2 output395 (.A(net395),
    .X(s1_wbd_dat_o[14]));
 sky130_fd_sc_hd__buf_2 output396 (.A(net396),
    .X(s1_wbd_dat_o[15]));
 sky130_fd_sc_hd__buf_2 output397 (.A(net397),
    .X(s1_wbd_dat_o[16]));
 sky130_fd_sc_hd__buf_2 output398 (.A(net398),
    .X(s1_wbd_dat_o[17]));
 sky130_fd_sc_hd__buf_2 output399 (.A(net399),
    .X(s1_wbd_dat_o[18]));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(ch_data_out[0]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net1450),
    .X(ch_data_out[132]));
 sky130_fd_sc_hd__buf_2 output400 (.A(net400),
    .X(s1_wbd_dat_o[19]));
 sky130_fd_sc_hd__buf_2 output401 (.A(net401),
    .X(s1_wbd_dat_o[1]));
 sky130_fd_sc_hd__buf_2 output402 (.A(net402),
    .X(s1_wbd_dat_o[20]));
 sky130_fd_sc_hd__buf_2 output403 (.A(net403),
    .X(s1_wbd_dat_o[21]));
 sky130_fd_sc_hd__buf_2 output404 (.A(net404),
    .X(s1_wbd_dat_o[22]));
 sky130_fd_sc_hd__buf_2 output405 (.A(net405),
    .X(s1_wbd_dat_o[23]));
 sky130_fd_sc_hd__buf_2 output406 (.A(net406),
    .X(s1_wbd_dat_o[24]));
 sky130_fd_sc_hd__buf_2 output407 (.A(net407),
    .X(s1_wbd_dat_o[25]));
 sky130_fd_sc_hd__buf_2 output408 (.A(net408),
    .X(s1_wbd_dat_o[26]));
 sky130_fd_sc_hd__buf_2 output409 (.A(net409),
    .X(s1_wbd_dat_o[27]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net1449),
    .X(ch_data_out[133]));
 sky130_fd_sc_hd__buf_2 output410 (.A(net410),
    .X(s1_wbd_dat_o[28]));
 sky130_fd_sc_hd__buf_2 output411 (.A(net411),
    .X(s1_wbd_dat_o[29]));
 sky130_fd_sc_hd__buf_2 output412 (.A(net412),
    .X(s1_wbd_dat_o[2]));
 sky130_fd_sc_hd__buf_2 output413 (.A(net413),
    .X(s1_wbd_dat_o[30]));
 sky130_fd_sc_hd__buf_2 output414 (.A(net414),
    .X(s1_wbd_dat_o[31]));
 sky130_fd_sc_hd__buf_2 output415 (.A(net415),
    .X(s1_wbd_dat_o[3]));
 sky130_fd_sc_hd__buf_2 output416 (.A(net416),
    .X(s1_wbd_dat_o[4]));
 sky130_fd_sc_hd__buf_2 output417 (.A(net417),
    .X(s1_wbd_dat_o[5]));
 sky130_fd_sc_hd__buf_2 output418 (.A(net418),
    .X(s1_wbd_dat_o[6]));
 sky130_fd_sc_hd__buf_2 output419 (.A(net419),
    .X(s1_wbd_dat_o[7]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net1448),
    .X(ch_data_out[134]));
 sky130_fd_sc_hd__buf_2 output420 (.A(net420),
    .X(s1_wbd_dat_o[8]));
 sky130_fd_sc_hd__buf_2 output421 (.A(net421),
    .X(s1_wbd_dat_o[9]));
 sky130_fd_sc_hd__buf_2 output422 (.A(net422),
    .X(s1_wbd_sel_o[0]));
 sky130_fd_sc_hd__buf_2 output423 (.A(net423),
    .X(s1_wbd_sel_o[1]));
 sky130_fd_sc_hd__buf_2 output424 (.A(net424),
    .X(s1_wbd_sel_o[2]));
 sky130_fd_sc_hd__buf_2 output425 (.A(net425),
    .X(s1_wbd_sel_o[3]));
 sky130_fd_sc_hd__buf_2 output426 (.A(net426),
    .X(s1_wbd_stb_o));
 sky130_fd_sc_hd__buf_2 output427 (.A(net427),
    .X(s1_wbd_we_o));
 sky130_fd_sc_hd__clkbuf_1 output428 (.A(net428),
    .X(s2_mclk));
 sky130_fd_sc_hd__buf_2 output429 (.A(net429),
    .X(s2_wbd_adr_o[10]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net1447),
    .X(ch_data_out[135]));
 sky130_fd_sc_hd__buf_2 output430 (.A(net430),
    .X(s2_wbd_adr_o[2]));
 sky130_fd_sc_hd__buf_2 output431 (.A(net431),
    .X(s2_wbd_adr_o[3]));
 sky130_fd_sc_hd__buf_2 output432 (.A(net432),
    .X(s2_wbd_adr_o[4]));
 sky130_fd_sc_hd__buf_2 output433 (.A(net433),
    .X(s2_wbd_adr_o[5]));
 sky130_fd_sc_hd__buf_2 output434 (.A(net434),
    .X(s2_wbd_adr_o[6]));
 sky130_fd_sc_hd__buf_2 output435 (.A(net435),
    .X(s2_wbd_adr_o[7]));
 sky130_fd_sc_hd__buf_2 output436 (.A(net436),
    .X(s2_wbd_adr_o[8]));
 sky130_fd_sc_hd__buf_2 output437 (.A(net437),
    .X(s2_wbd_adr_o[9]));
 sky130_fd_sc_hd__buf_2 output438 (.A(net438),
    .X(s2_wbd_cyc_o));
 sky130_fd_sc_hd__buf_2 output439 (.A(net439),
    .X(s2_wbd_dat_o[0]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net1446),
    .X(ch_data_out[136]));
 sky130_fd_sc_hd__buf_2 output440 (.A(net440),
    .X(s2_wbd_dat_o[10]));
 sky130_fd_sc_hd__buf_2 output441 (.A(net441),
    .X(s2_wbd_dat_o[11]));
 sky130_fd_sc_hd__buf_2 output442 (.A(net442),
    .X(s2_wbd_dat_o[12]));
 sky130_fd_sc_hd__buf_2 output443 (.A(net443),
    .X(s2_wbd_dat_o[13]));
 sky130_fd_sc_hd__buf_2 output444 (.A(net444),
    .X(s2_wbd_dat_o[14]));
 sky130_fd_sc_hd__buf_2 output445 (.A(net445),
    .X(s2_wbd_dat_o[15]));
 sky130_fd_sc_hd__buf_2 output446 (.A(net446),
    .X(s2_wbd_dat_o[16]));
 sky130_fd_sc_hd__buf_2 output447 (.A(net447),
    .X(s2_wbd_dat_o[17]));
 sky130_fd_sc_hd__buf_2 output448 (.A(net448),
    .X(s2_wbd_dat_o[18]));
 sky130_fd_sc_hd__buf_2 output449 (.A(net449),
    .X(s2_wbd_dat_o[19]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net1445),
    .X(ch_data_out[137]));
 sky130_fd_sc_hd__buf_2 output450 (.A(net450),
    .X(s2_wbd_dat_o[1]));
 sky130_fd_sc_hd__buf_2 output451 (.A(net451),
    .X(s2_wbd_dat_o[20]));
 sky130_fd_sc_hd__buf_2 output452 (.A(net452),
    .X(s2_wbd_dat_o[21]));
 sky130_fd_sc_hd__buf_2 output453 (.A(net453),
    .X(s2_wbd_dat_o[22]));
 sky130_fd_sc_hd__buf_2 output454 (.A(net454),
    .X(s2_wbd_dat_o[23]));
 sky130_fd_sc_hd__buf_2 output455 (.A(net455),
    .X(s2_wbd_dat_o[24]));
 sky130_fd_sc_hd__buf_2 output456 (.A(net456),
    .X(s2_wbd_dat_o[25]));
 sky130_fd_sc_hd__buf_2 output457 (.A(net457),
    .X(s2_wbd_dat_o[26]));
 sky130_fd_sc_hd__buf_2 output458 (.A(net458),
    .X(s2_wbd_dat_o[27]));
 sky130_fd_sc_hd__buf_2 output459 (.A(net459),
    .X(s2_wbd_dat_o[28]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net1444),
    .X(ch_data_out[138]));
 sky130_fd_sc_hd__buf_2 output460 (.A(net460),
    .X(s2_wbd_dat_o[29]));
 sky130_fd_sc_hd__buf_2 output461 (.A(net461),
    .X(s2_wbd_dat_o[2]));
 sky130_fd_sc_hd__buf_2 output462 (.A(net462),
    .X(s2_wbd_dat_o[30]));
 sky130_fd_sc_hd__buf_2 output463 (.A(net463),
    .X(s2_wbd_dat_o[31]));
 sky130_fd_sc_hd__buf_2 output464 (.A(net464),
    .X(s2_wbd_dat_o[3]));
 sky130_fd_sc_hd__buf_2 output465 (.A(net465),
    .X(s2_wbd_dat_o[4]));
 sky130_fd_sc_hd__buf_2 output466 (.A(net466),
    .X(s2_wbd_dat_o[5]));
 sky130_fd_sc_hd__buf_2 output467 (.A(net467),
    .X(s2_wbd_dat_o[6]));
 sky130_fd_sc_hd__buf_2 output468 (.A(net468),
    .X(s2_wbd_dat_o[7]));
 sky130_fd_sc_hd__buf_2 output469 (.A(net469),
    .X(s2_wbd_dat_o[8]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net1443),
    .X(ch_data_out[139]));
 sky130_fd_sc_hd__buf_2 output470 (.A(net470),
    .X(s2_wbd_dat_o[9]));
 sky130_fd_sc_hd__buf_2 output471 (.A(net471),
    .X(s2_wbd_sel_o[0]));
 sky130_fd_sc_hd__buf_2 output472 (.A(net472),
    .X(s2_wbd_sel_o[1]));
 sky130_fd_sc_hd__buf_2 output473 (.A(net473),
    .X(s2_wbd_sel_o[2]));
 sky130_fd_sc_hd__buf_2 output474 (.A(net474),
    .X(s2_wbd_sel_o[3]));
 sky130_fd_sc_hd__buf_2 output475 (.A(net475),
    .X(s2_wbd_stb_o));
 sky130_fd_sc_hd__buf_2 output476 (.A(net476),
    .X(s2_wbd_we_o));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(ch_data_out[13]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net1442),
    .X(ch_data_out[140]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(ch_data_out[100]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net1441),
    .X(ch_data_out[141]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net1440),
    .X(ch_data_out[142]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net1439),
    .X(ch_data_out[143]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net1438),
    .X(ch_data_out[144]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net1437),
    .X(ch_data_out[145]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net1434),
    .X(ch_data_out[146]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net1431),
    .X(ch_data_out[147]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net1428),
    .X(ch_data_out[148]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net1425),
    .X(ch_data_out[149]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(ch_data_out[14]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(ch_data_out[101]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(ch_data_out[150]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(ch_data_out[151]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net1422),
    .X(ch_data_out[152]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net1419),
    .X(ch_data_out[153]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net1416),
    .X(ch_data_out[154]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(ch_data_out[155]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(ch_data_out[156]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(ch_data_out[157]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(ch_data_out[15]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(ch_data_out[16]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(ch_data_out[102]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(ch_data_out[17]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(ch_data_out[18]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(ch_data_out[19]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(ch_data_out[1]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(ch_data_out[20]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(ch_data_out[21]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(ch_data_out[22]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(ch_data_out[23]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(ch_data_out[24]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(ch_data_out[25]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(ch_data_out[103]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(ch_data_out[26]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(ch_data_out[27]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(ch_data_out[28]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(ch_data_out[29]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(ch_data_out[2]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(ch_data_out[30]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(ch_data_out[31]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(ch_data_out[32]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(ch_data_out[33]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(ch_data_out[34]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(ch_data_out[104]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(ch_data_out[35]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(ch_data_out[36]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(ch_data_out[37]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(ch_data_out[38]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(ch_data_out[39]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(ch_data_out[3]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(ch_data_out[40]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(ch_data_out[41]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(ch_data_out[42]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(ch_data_out[43]));
 sky130_fd_sc_hd__buf_2 rebuffer1 (.A(_1855_),
    .X(net1774));
 sky130_fd_sc_hd__buf_2 rebuffer2 (.A(_1956_),
    .X(net1775));
 sky130_fd_sc_hd__buf_4 rebuffer3 (.A(_2259_),
    .X(net1776));
 sky130_fd_sc_hd__buf_6 split4 (.A(net814),
    .X(net1777));
 sky130_fd_sc_hd__dlclkp_2 \u_dcg_peri.u_clkgate.u_gate  (.CLK(net1772),
    .GATE(net1411),
    .GCLK(net298));
 sky130_fd_sc_hd__dlclkp_2 \u_dcg_riscv.u_clkgate.u_gate  (.CLK(net1768),
    .GATE(net1413),
    .GCLK(net299));
 sky130_fd_sc_hd__dlclkp_2 \u_dcg_s0.u_clkgate.u_gate  (.CLK(net1768),
    .GATE(net572),
    .GCLK(net300));
 sky130_fd_sc_hd__dlclkp_2 \u_dcg_s1.u_clkgate.u_gate  (.CLK(net1767),
    .GATE(\u_dcg_s1.clk_enb ),
    .GCLK(net381));
 sky130_fd_sc_hd__dlclkp_2 \u_dcg_s2.u_clkgate.u_gate  (.CLK(net1773),
    .GATE(net1415),
    .GCLK(net428));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[0].u_dsync0  (.CLK(\clknet_leaf_58_u_dsync.out_clk ),
    .D(\u_dcg_s0.clk_enb ),
    .RESET_B(net880),
    .Q(\u_dsync.in_data_s[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[0].u_dsync1  (.CLK(\clknet_leaf_37_u_dsync.out_clk ),
    .D(\u_dsync.in_data_s[0] ),
    .RESET_B(net878),
    .Q(\u_dsync.in_data_2s[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[0].u_dsync2  (.CLK(\clknet_leaf_37_u_dsync.out_clk ),
    .D(net1975),
    .RESET_B(net878),
    .Q(\u_dsync.out_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[1].u_dsync0  (.CLK(\clknet_leaf_7_u_dsync.out_clk ),
    .D(\u_dcg_s1.clk_enb ),
    .RESET_B(net857),
    .Q(\u_dsync.in_data_s[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[1].u_dsync1  (.CLK(\clknet_leaf_7_u_dsync.out_clk ),
    .D(net1969),
    .RESET_B(net857),
    .Q(\u_dsync.in_data_2s[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[1].u_dsync2  (.CLK(\clknet_leaf_6_u_dsync.out_clk ),
    .D(\u_dsync.in_data_2s[1] ),
    .RESET_B(net857),
    .Q(\u_dsync.out_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[2].u_dsync0  (.CLK(\clknet_leaf_12_u_dsync.out_clk ),
    .D(net1415),
    .RESET_B(net886),
    .Q(\u_dsync.in_data_s[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[2].u_dsync1  (.CLK(\clknet_leaf_12_u_dsync.out_clk ),
    .D(\u_dsync.in_data_s[2] ),
    .RESET_B(net883),
    .Q(\u_dsync.in_data_2s[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[2].u_dsync2  (.CLK(\clknet_leaf_12_u_dsync.out_clk ),
    .D(net1965),
    .RESET_B(net887),
    .Q(\u_dsync.out_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[3].u_dsync0  (.CLK(\clknet_leaf_14_u_dsync.out_clk ),
    .D(net1412),
    .RESET_B(net868),
    .Q(\u_dsync.in_data_s[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[3].u_dsync1  (.CLK(\clknet_leaf_14_u_dsync.out_clk ),
    .D(net1960),
    .RESET_B(net869),
    .Q(\u_dsync.in_data_2s[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[3].u_dsync2  (.CLK(\clknet_leaf_10_u_dsync.out_clk ),
    .D(net1940),
    .RESET_B(net869),
    .Q(\u_dsync.out_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[4].u_dsync0  (.CLK(\clknet_leaf_15_u_dsync.out_clk ),
    .D(\u_dcg_riscv.clk_enb ),
    .RESET_B(net876),
    .Q(\u_dsync.in_data_s[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[4].u_dsync1  (.CLK(\clknet_leaf_17_u_dsync.out_clk ),
    .D(\u_dsync.in_data_s[4] ),
    .RESET_B(net876),
    .Q(\u_dsync.in_data_2s[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[4].u_dsync2  (.CLK(\clknet_leaf_19_u_dsync.out_clk ),
    .D(net1944),
    .RESET_B(net884),
    .Q(\u_dsync.out_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[5].u_dsync0  (.CLK(\clknet_leaf_24_u_dsync.out_clk ),
    .D(net1717),
    .RESET_B(net911),
    .Q(\u_dsync.in_data_s[5] ));
 sky130_fd_sc_hd__conb_1 \u_dsync.bus_.bit_[5].u_dsync0_1717  (.LO(net1717));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[5].u_dsync1  (.CLK(\clknet_leaf_24_u_dsync.out_clk ),
    .D(net1959),
    .RESET_B(net912),
    .Q(\u_dsync.in_data_2s[5] ));
 sky130_fd_sc_hd__dfrtp_4 \u_dsync.bus_.bit_[5].u_dsync2  (.CLK(\clknet_leaf_24_u_dsync.out_clk ),
    .D(\u_dsync.in_data_2s[5] ),
    .RESET_B(net910),
    .Q(\u_dsync.out_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[6].u_dsync0  (.CLK(\clknet_leaf_21_u_dsync.out_clk ),
    .D(net1718),
    .RESET_B(net900),
    .Q(\u_dsync.in_data_s[6] ));
 sky130_fd_sc_hd__conb_1 \u_dsync.bus_.bit_[6].u_dsync0_1718  (.LO(net1718));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[6].u_dsync1  (.CLK(\clknet_leaf_26_u_dsync.out_clk ),
    .D(net1972),
    .RESET_B(net900),
    .Q(\u_dsync.in_data_2s[6] ));
 sky130_fd_sc_hd__dfrtp_2 \u_dsync.bus_.bit_[6].u_dsync2  (.CLK(\clknet_leaf_26_u_dsync.out_clk ),
    .D(net1966),
    .RESET_B(net900),
    .Q(\u_dsync.out_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[7].u_dsync0  (.CLK(\clknet_leaf_24_u_dsync.out_clk ),
    .D(net1719),
    .RESET_B(net910),
    .Q(\u_dsync.in_data_s[7] ));
 sky130_fd_sc_hd__conb_1 \u_dsync.bus_.bit_[7].u_dsync0_1719  (.LO(net1719));
 sky130_fd_sc_hd__dfrtp_1 \u_dsync.bus_.bit_[7].u_dsync1  (.CLK(\clknet_leaf_25_u_dsync.out_clk ),
    .D(net1956),
    .RESET_B(net911),
    .Q(\u_dsync.in_data_2s[7] ));
 sky130_fd_sc_hd__dfrtp_4 \u_dsync.bus_.bit_[7].u_dsync2  (.CLK(\clknet_leaf_29_u_dsync.out_clk ),
    .D(net1823),
    .RESET_B(net911),
    .Q(\u_dsync.out_data[7] ));
 sky130_fd_sc_hd__mux2_4 \u_rst_sync.u_buf.genblk1.u_mux  (.A0(net1878),
    .A1(rst_n),
    .S(net1720),
    .X(\u_dcg_peri.reset_n ));
 sky130_fd_sc_hd__conb_1 \u_rst_sync.u_buf.genblk1.u_mux_1720  (.LO(net1720));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_1.u_dly0  (.A(\u_skew_wi.clk_inbuf ),
    .X(\u_skew_wi.clkbuf_1.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_1.u_dly1  (.A(\u_skew_wi.clkbuf_1.X1 ),
    .X(\u_skew_wi.clkbuf_1.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_1.u_dly2  (.A(\u_skew_wi.clkbuf_1.X2 ),
    .X(\u_skew_wi.clkbuf_1.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_1.u_dly3  (.A(\u_skew_wi.clkbuf_1.X3 ),
    .X(\u_skew_wi.clk_d1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_10.u_dly0  (.A(\u_skew_wi.clk_d9 ),
    .X(\u_skew_wi.clkbuf_10.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_10.u_dly1  (.A(\u_skew_wi.clkbuf_10.X1 ),
    .X(\u_skew_wi.clkbuf_10.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_10.u_dly2  (.A(\u_skew_wi.clkbuf_10.X2 ),
    .X(\u_skew_wi.clkbuf_10.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_10.u_dly3  (.A(\u_skew_wi.clkbuf_10.X3 ),
    .X(\u_skew_wi.clk_d10 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_11.u_dly0  (.A(\u_skew_wi.clk_d10 ),
    .X(\u_skew_wi.clkbuf_11.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_11.u_dly1  (.A(\u_skew_wi.clkbuf_11.X1 ),
    .X(\u_skew_wi.clkbuf_11.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_11.u_dly2  (.A(\u_skew_wi.clkbuf_11.X2 ),
    .X(\u_skew_wi.clkbuf_11.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_11.u_dly3  (.A(\u_skew_wi.clkbuf_11.X3 ),
    .X(\u_skew_wi.clk_d11 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_12.u_dly0  (.A(\u_skew_wi.clk_d11 ),
    .X(\u_skew_wi.clkbuf_12.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_12.u_dly1  (.A(\u_skew_wi.clkbuf_12.X1 ),
    .X(\u_skew_wi.clkbuf_12.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_12.u_dly2  (.A(\u_skew_wi.clkbuf_12.X2 ),
    .X(\u_skew_wi.clkbuf_12.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_12.u_dly3  (.A(\u_skew_wi.clkbuf_12.X3 ),
    .X(\u_skew_wi.clk_d12 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_13.u_dly0  (.A(\u_skew_wi.clk_d12 ),
    .X(\u_skew_wi.clkbuf_13.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_13.u_dly1  (.A(\u_skew_wi.clkbuf_13.X1 ),
    .X(\u_skew_wi.clkbuf_13.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_13.u_dly2  (.A(\u_skew_wi.clkbuf_13.X2 ),
    .X(\u_skew_wi.clkbuf_13.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_13.u_dly3  (.A(\u_skew_wi.clkbuf_13.X3 ),
    .X(\u_skew_wi.clk_d13 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_14.u_dly0  (.A(\u_skew_wi.clk_d13 ),
    .X(\u_skew_wi.clkbuf_14.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_14.u_dly1  (.A(\u_skew_wi.clkbuf_14.X1 ),
    .X(\u_skew_wi.clkbuf_14.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_14.u_dly2  (.A(\u_skew_wi.clkbuf_14.X2 ),
    .X(\u_skew_wi.clkbuf_14.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_14.u_dly3  (.A(\u_skew_wi.clkbuf_14.X3 ),
    .X(\u_skew_wi.clk_d14 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_15.u_dly0  (.A(\u_skew_wi.clk_d14 ),
    .X(\u_skew_wi.clkbuf_15.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_15.u_dly1  (.A(\u_skew_wi.clkbuf_15.X1 ),
    .X(\u_skew_wi.clkbuf_15.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_15.u_dly2  (.A(\u_skew_wi.clkbuf_15.X2 ),
    .X(\u_skew_wi.clkbuf_15.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_15.u_dly3  (.A(\u_skew_wi.clkbuf_15.X3 ),
    .X(\u_skew_wi.clk_d15 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_2.u_dly0  (.A(\u_skew_wi.clk_d1 ),
    .X(\u_skew_wi.clkbuf_2.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_2.u_dly1  (.A(\u_skew_wi.clkbuf_2.X1 ),
    .X(\u_skew_wi.clkbuf_2.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_2.u_dly2  (.A(\u_skew_wi.clkbuf_2.X2 ),
    .X(\u_skew_wi.clkbuf_2.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_2.u_dly3  (.A(\u_skew_wi.clkbuf_2.X3 ),
    .X(\u_skew_wi.clk_d2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_3.u_dly0  (.A(\u_skew_wi.clk_d2 ),
    .X(\u_skew_wi.clkbuf_3.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_3.u_dly1  (.A(\u_skew_wi.clkbuf_3.X1 ),
    .X(\u_skew_wi.clkbuf_3.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_3.u_dly2  (.A(\u_skew_wi.clkbuf_3.X2 ),
    .X(\u_skew_wi.clkbuf_3.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_3.u_dly3  (.A(\u_skew_wi.clkbuf_3.X3 ),
    .X(\u_skew_wi.clk_d3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_4.u_dly0  (.A(\u_skew_wi.clk_d3 ),
    .X(\u_skew_wi.clkbuf_4.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_4.u_dly1  (.A(\u_skew_wi.clkbuf_4.X1 ),
    .X(\u_skew_wi.clkbuf_4.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_4.u_dly2  (.A(\u_skew_wi.clkbuf_4.X2 ),
    .X(\u_skew_wi.clkbuf_4.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_4.u_dly3  (.A(\u_skew_wi.clkbuf_4.X3 ),
    .X(\u_skew_wi.clk_d4 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_5.u_dly0  (.A(\u_skew_wi.clk_d4 ),
    .X(\u_skew_wi.clkbuf_5.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_5.u_dly1  (.A(\u_skew_wi.clkbuf_5.X1 ),
    .X(\u_skew_wi.clkbuf_5.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_5.u_dly2  (.A(\u_skew_wi.clkbuf_5.X2 ),
    .X(\u_skew_wi.clkbuf_5.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_5.u_dly3  (.A(\u_skew_wi.clkbuf_5.X3 ),
    .X(\u_skew_wi.clk_d5 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_6.u_dly0  (.A(\u_skew_wi.clk_d5 ),
    .X(\u_skew_wi.clkbuf_6.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_6.u_dly1  (.A(\u_skew_wi.clkbuf_6.X1 ),
    .X(\u_skew_wi.clkbuf_6.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_6.u_dly2  (.A(\u_skew_wi.clkbuf_6.X2 ),
    .X(\u_skew_wi.clkbuf_6.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_6.u_dly3  (.A(\u_skew_wi.clkbuf_6.X3 ),
    .X(\u_skew_wi.clk_d6 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_7.u_dly0  (.A(\u_skew_wi.clk_d6 ),
    .X(\u_skew_wi.clkbuf_7.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_7.u_dly1  (.A(\u_skew_wi.clkbuf_7.X1 ),
    .X(\u_skew_wi.clkbuf_7.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_7.u_dly2  (.A(\u_skew_wi.clkbuf_7.X2 ),
    .X(\u_skew_wi.clkbuf_7.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_7.u_dly3  (.A(\u_skew_wi.clkbuf_7.X3 ),
    .X(\u_skew_wi.clk_d7 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_8.u_dly0  (.A(\u_skew_wi.clk_d7 ),
    .X(\u_skew_wi.clkbuf_8.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_8.u_dly1  (.A(\u_skew_wi.clkbuf_8.X1 ),
    .X(\u_skew_wi.clkbuf_8.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_8.u_dly2  (.A(\u_skew_wi.clkbuf_8.X2 ),
    .X(\u_skew_wi.clkbuf_8.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_8.u_dly3  (.A(\u_skew_wi.clkbuf_8.X3 ),
    .X(\u_skew_wi.clk_d8 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_9.u_dly0  (.A(\u_skew_wi.clk_d8 ),
    .X(\u_skew_wi.clkbuf_9.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_9.u_dly1  (.A(\u_skew_wi.clkbuf_9.X1 ),
    .X(\u_skew_wi.clkbuf_9.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_9.u_dly2  (.A(\u_skew_wi.clkbuf_9.X2 ),
    .X(\u_skew_wi.clkbuf_9.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wi.clkbuf_9.u_dly3  (.A(\u_skew_wi.clkbuf_9.X3 ),
    .X(\u_skew_wi.clk_d9 ));
 sky130_fd_sc_hd__clkbuf_8 \u_skew_wi.u_clkbuf_in.u_buf  (.A(wbd_clk_int),
    .X(\u_skew_wi.clk_inbuf ));
 sky130_fd_sc_hd__clkbuf_8 \u_skew_wi.u_clkbuf_out.u_buf  (.A(\u_skew_wi.d30 ),
    .X(wbd_clk_wi));
 sky130_fd_sc_hd__mux2_2 \u_skew_wi.u_mux_level_00.genblk1.u_mux  (.A0(\u_skew_wi.in0 ),
    .A1(\u_skew_wi.in1 ),
    .S(cfg_cska_wi[0]),
    .X(\u_skew_wi.d00 ));
 sky130_fd_sc_hd__mux2_2 \u_skew_wi.u_mux_level_01.genblk1.u_mux  (.A0(\u_skew_wi.in2 ),
    .A1(\u_skew_wi.in3 ),
    .S(cfg_cska_wi[0]),
    .X(\u_skew_wi.d01 ));
 sky130_fd_sc_hd__mux2_2 \u_skew_wi.u_mux_level_02.genblk1.u_mux  (.A0(\u_skew_wi.in4 ),
    .A1(\u_skew_wi.in5 ),
    .S(cfg_cska_wi[0]),
    .X(\u_skew_wi.d02 ));
 sky130_fd_sc_hd__mux2_2 \u_skew_wi.u_mux_level_03.genblk1.u_mux  (.A0(\u_skew_wi.in6 ),
    .A1(\u_skew_wi.in7 ),
    .S(cfg_cska_wi[0]),
    .X(\u_skew_wi.d03 ));
 sky130_fd_sc_hd__mux2_2 \u_skew_wi.u_mux_level_04.genblk1.u_mux  (.A0(\u_skew_wi.in8 ),
    .A1(\u_skew_wi.in9 ),
    .S(cfg_cska_wi[0]),
    .X(\u_skew_wi.d04 ));
 sky130_fd_sc_hd__mux2_2 \u_skew_wi.u_mux_level_05.genblk1.u_mux  (.A0(\u_skew_wi.in10 ),
    .A1(\u_skew_wi.in11 ),
    .S(cfg_cska_wi[0]),
    .X(\u_skew_wi.d05 ));
 sky130_fd_sc_hd__mux2_2 \u_skew_wi.u_mux_level_06.genblk1.u_mux  (.A0(\u_skew_wi.in12 ),
    .A1(\u_skew_wi.in13 ),
    .S(cfg_cska_wi[0]),
    .X(\u_skew_wi.d06 ));
 sky130_fd_sc_hd__mux2_2 \u_skew_wi.u_mux_level_07.genblk1.u_mux  (.A0(\u_skew_wi.in14 ),
    .A1(\u_skew_wi.in15 ),
    .S(cfg_cska_wi[0]),
    .X(\u_skew_wi.d07 ));
 sky130_fd_sc_hd__mux2_2 \u_skew_wi.u_mux_level_10.genblk1.u_mux  (.A0(\u_skew_wi.d00 ),
    .A1(\u_skew_wi.d01 ),
    .S(cfg_cska_wi[1]),
    .X(\u_skew_wi.d10 ));
 sky130_fd_sc_hd__mux2_2 \u_skew_wi.u_mux_level_11.genblk1.u_mux  (.A0(\u_skew_wi.d02 ),
    .A1(\u_skew_wi.d03 ),
    .S(cfg_cska_wi[1]),
    .X(\u_skew_wi.d11 ));
 sky130_fd_sc_hd__mux2_2 \u_skew_wi.u_mux_level_12.genblk1.u_mux  (.A0(\u_skew_wi.d04 ),
    .A1(\u_skew_wi.d05 ),
    .S(cfg_cska_wi[1]),
    .X(\u_skew_wi.d12 ));
 sky130_fd_sc_hd__mux2_2 \u_skew_wi.u_mux_level_13.genblk1.u_mux  (.A0(\u_skew_wi.d06 ),
    .A1(\u_skew_wi.d07 ),
    .S(cfg_cska_wi[1]),
    .X(\u_skew_wi.d13 ));
 sky130_fd_sc_hd__mux2_2 \u_skew_wi.u_mux_level_20.genblk1.u_mux  (.A0(\u_skew_wi.d10 ),
    .A1(\u_skew_wi.d11 ),
    .S(cfg_cska_wi[2]),
    .X(\u_skew_wi.d20 ));
 sky130_fd_sc_hd__mux2_2 \u_skew_wi.u_mux_level_21.genblk1.u_mux  (.A0(\u_skew_wi.d12 ),
    .A1(\u_skew_wi.d13 ),
    .S(cfg_cska_wi[2]),
    .X(\u_skew_wi.d21 ));
 sky130_fd_sc_hd__mux2_4 \u_skew_wi.u_mux_level_30.genblk1.u_mux  (.A0(\u_skew_wi.d20 ),
    .A1(\u_skew_wi.d21 ),
    .S(cfg_cska_wi[3]),
    .X(\u_skew_wi.d30 ));
 sky130_fd_sc_hd__clkbuf_8 \u_skew_wi.u_tap_0.u_buf  (.A(\u_skew_wi.clk_inbuf ),
    .X(\u_skew_wi.in0 ));
 sky130_fd_sc_hd__clkbuf_8 \u_skew_wi.u_tap_1.u_buf  (.A(\u_skew_wi.clk_d1 ),
    .X(\u_skew_wi.in1 ));
 sky130_fd_sc_hd__clkbuf_8 \u_skew_wi.u_tap_10.u_buf  (.A(\u_skew_wi.clk_d10 ),
    .X(\u_skew_wi.in10 ));
 sky130_fd_sc_hd__clkbuf_8 \u_skew_wi.u_tap_11.u_buf  (.A(\u_skew_wi.clk_d11 ),
    .X(\u_skew_wi.in11 ));
 sky130_fd_sc_hd__clkbuf_8 \u_skew_wi.u_tap_12.u_buf  (.A(\u_skew_wi.clk_d12 ),
    .X(\u_skew_wi.in12 ));
 sky130_fd_sc_hd__clkbuf_8 \u_skew_wi.u_tap_13.u_buf  (.A(\u_skew_wi.clk_d13 ),
    .X(\u_skew_wi.in13 ));
 sky130_fd_sc_hd__clkbuf_8 \u_skew_wi.u_tap_14.u_buf  (.A(\u_skew_wi.clk_d14 ),
    .X(\u_skew_wi.in14 ));
 sky130_fd_sc_hd__clkbuf_8 \u_skew_wi.u_tap_15.u_buf  (.A(\u_skew_wi.clk_d15 ),
    .X(\u_skew_wi.in15 ));
 sky130_fd_sc_hd__clkbuf_8 \u_skew_wi.u_tap_2.u_buf  (.A(\u_skew_wi.clk_d2 ),
    .X(\u_skew_wi.in2 ));
 sky130_fd_sc_hd__clkbuf_8 \u_skew_wi.u_tap_3.u_buf  (.A(\u_skew_wi.clk_d3 ),
    .X(\u_skew_wi.in3 ));
 sky130_fd_sc_hd__clkbuf_8 \u_skew_wi.u_tap_4.u_buf  (.A(\u_skew_wi.clk_d4 ),
    .X(\u_skew_wi.in4 ));
 sky130_fd_sc_hd__clkbuf_8 \u_skew_wi.u_tap_5.u_buf  (.A(\u_skew_wi.clk_d5 ),
    .X(\u_skew_wi.in5 ));
 sky130_fd_sc_hd__clkbuf_8 \u_skew_wi.u_tap_6.u_buf  (.A(\u_skew_wi.clk_d6 ),
    .X(\u_skew_wi.in6 ));
 sky130_fd_sc_hd__clkbuf_8 \u_skew_wi.u_tap_7.u_buf  (.A(\u_skew_wi.clk_d7 ),
    .X(\u_skew_wi.in7 ));
 sky130_fd_sc_hd__clkbuf_8 \u_skew_wi.u_tap_8.u_buf  (.A(\u_skew_wi.clk_d8 ),
    .X(\u_skew_wi.in8 ));
 sky130_fd_sc_hd__clkbuf_8 \u_skew_wi.u_tap_9.u_buf  (.A(\u_skew_wi.clk_d9 ),
    .X(\u_skew_wi.in9 ));
 sky130_fd_sc_hd__dlclkp_2 \u_wbi_clkgate.u_gate  (.CLK(clk_i),
    .GATE(net1732),
    .GCLK(\u_dsync.out_clk ));
 sky130_fd_sc_hd__conb_1 \u_wbi_clkgate.u_gate_1732  (.HI(net1732));
 sky130_fd_sc_hd__conb_1 wb_interconnect_1721 (.LO(net1721));
 sky130_fd_sc_hd__conb_1 wb_interconnect_1722 (.LO(net1722));
 sky130_fd_sc_hd__conb_1 wb_interconnect_1723 (.LO(net1723));
 sky130_fd_sc_hd__conb_1 wb_interconnect_1724 (.LO(net1724));
 sky130_fd_sc_hd__conb_1 wb_interconnect_1725 (.LO(net1725));
 sky130_fd_sc_hd__conb_1 wb_interconnect_1726 (.LO(net1726));
 sky130_fd_sc_hd__conb_1 wb_interconnect_1727 (.LO(net1727));
 sky130_fd_sc_hd__conb_1 wb_interconnect_1728 (.LO(net1728));
 sky130_fd_sc_hd__conb_1 wb_interconnect_1729 (.LO(net1729));
 sky130_fd_sc_hd__conb_1 wb_interconnect_1730 (.LO(net1730));
 sky130_fd_sc_hd__buf_6 wire1 (.A(net1734),
    .X(net1733));
 sky130_fd_sc_hd__clkbuf_8 wire10 (.A(\clknet_3_0__leaf_u_dsync.out_clk ),
    .X(net1742));
 sky130_fd_sc_hd__buf_4 wire1007 (.A(_2187_),
    .X(net1007));
 sky130_fd_sc_hd__buf_4 wire1008 (.A(net1009),
    .X(net1008));
 sky130_fd_sc_hd__buf_4 wire1009 (.A(_2186_),
    .X(net1009));
 sky130_fd_sc_hd__buf_6 wire1010 (.A(_2184_),
    .X(net1010));
 sky130_fd_sc_hd__buf_4 wire1011 (.A(net1012),
    .X(net1011));
 sky130_fd_sc_hd__buf_6 wire1012 (.A(_2182_),
    .X(net1012));
 sky130_fd_sc_hd__buf_4 wire1013 (.A(_2181_),
    .X(net1013));
 sky130_fd_sc_hd__buf_4 wire1014 (.A(_2179_),
    .X(net1014));
 sky130_fd_sc_hd__buf_4 wire1015 (.A(net1016),
    .X(net1015));
 sky130_fd_sc_hd__buf_4 wire1016 (.A(_2177_),
    .X(net1016));
 sky130_fd_sc_hd__buf_4 wire1017 (.A(_2176_),
    .X(net1017));
 sky130_fd_sc_hd__buf_4 wire1018 (.A(_2174_),
    .X(net1018));
 sky130_fd_sc_hd__buf_4 wire1019 (.A(_2172_),
    .X(net1019));
 sky130_fd_sc_hd__buf_4 wire1020 (.A(net1021),
    .X(net1020));
 sky130_fd_sc_hd__buf_6 wire1021 (.A(_2171_),
    .X(net1021));
 sky130_fd_sc_hd__buf_4 wire1022 (.A(_2169_),
    .X(net1022));
 sky130_fd_sc_hd__buf_4 wire1023 (.A(net1024),
    .X(net1023));
 sky130_fd_sc_hd__buf_6 wire1024 (.A(net1025),
    .X(net1024));
 sky130_fd_sc_hd__buf_4 wire1025 (.A(_2167_),
    .X(net1025));
 sky130_fd_sc_hd__buf_4 wire1026 (.A(_2166_),
    .X(net1026));
 sky130_fd_sc_hd__buf_4 wire1027 (.A(_2164_),
    .X(net1027));
 sky130_fd_sc_hd__buf_4 wire1028 (.A(net1029),
    .X(net1028));
 sky130_fd_sc_hd__buf_4 wire1029 (.A(_2162_),
    .X(net1029));
 sky130_fd_sc_hd__buf_4 wire1030 (.A(_2161_),
    .X(net1030));
 sky130_fd_sc_hd__buf_4 wire1031 (.A(_2159_),
    .X(net1031));
 sky130_fd_sc_hd__buf_4 wire1032 (.A(net1033),
    .X(net1032));
 sky130_fd_sc_hd__buf_4 wire1033 (.A(_2157_),
    .X(net1033));
 sky130_fd_sc_hd__buf_4 wire1034 (.A(_2156_),
    .X(net1034));
 sky130_fd_sc_hd__buf_4 wire1035 (.A(_2154_),
    .X(net1035));
 sky130_fd_sc_hd__buf_12 wire1037 (.A(_2151_),
    .X(net1037));
 sky130_fd_sc_hd__clkbuf_8 wire1038 (.A(_2149_),
    .X(net1038));
 sky130_fd_sc_hd__buf_4 wire1039 (.A(_2147_),
    .X(net1039));
 sky130_fd_sc_hd__buf_4 wire1040 (.A(net1041),
    .X(net1040));
 sky130_fd_sc_hd__buf_6 wire1041 (.A(net1042),
    .X(net1041));
 sky130_fd_sc_hd__buf_4 wire1042 (.A(_2146_),
    .X(net1042));
 sky130_fd_sc_hd__buf_4 wire1043 (.A(_2142_),
    .X(net1043));
 sky130_fd_sc_hd__buf_4 wire1044 (.A(net1045),
    .X(net1044));
 sky130_fd_sc_hd__buf_6 wire1045 (.A(_2141_),
    .X(net1045));
 sky130_fd_sc_hd__buf_4 wire1046 (.A(_2139_),
    .X(net1046));
 sky130_fd_sc_hd__buf_4 wire1047 (.A(_2137_),
    .X(net1047));
 sky130_fd_sc_hd__buf_4 wire1048 (.A(net1049),
    .X(net1048));
 sky130_fd_sc_hd__buf_6 wire1049 (.A(_2136_),
    .X(net1049));
 sky130_fd_sc_hd__buf_4 wire1051 (.A(net1052),
    .X(net1051));
 sky130_fd_sc_hd__buf_6 wire1052 (.A(net1053),
    .X(net1052));
 sky130_fd_sc_hd__buf_4 wire1053 (.A(_2132_),
    .X(net1053));
 sky130_fd_sc_hd__buf_4 wire1054 (.A(_2131_),
    .X(net1054));
 sky130_fd_sc_hd__buf_4 wire1055 (.A(_2129_),
    .X(net1055));
 sky130_fd_sc_hd__buf_12 wire1056 (.A(_2127_),
    .X(net1056));
 sky130_fd_sc_hd__buf_6 wire1057 (.A(_2124_),
    .X(net1057));
 sky130_fd_sc_hd__buf_4 wire1058 (.A(net1059),
    .X(net1058));
 sky130_fd_sc_hd__buf_6 wire1059 (.A(_2122_),
    .X(net1059));
 sky130_fd_sc_hd__buf_4 wire1060 (.A(net1061),
    .X(net1060));
 sky130_fd_sc_hd__buf_6 wire1061 (.A(net1062),
    .X(net1061));
 sky130_fd_sc_hd__buf_4 wire1062 (.A(_2121_),
    .X(net1062));
 sky130_fd_sc_hd__buf_6 wire1063 (.A(_2119_),
    .X(net1063));
 sky130_fd_sc_hd__buf_12 wire1064 (.A(net1065),
    .X(net1064));
 sky130_fd_sc_hd__buf_6 wire1065 (.A(_2117_),
    .X(net1065));
 sky130_fd_sc_hd__buf_6 wire1066 (.A(_2116_),
    .X(net1066));
 sky130_fd_sc_hd__buf_6 wire1067 (.A(_2114_),
    .X(net1067));
 sky130_fd_sc_hd__buf_4 wire1068 (.A(net1069),
    .X(net1068));
 sky130_fd_sc_hd__buf_6 wire1069 (.A(_2112_),
    .X(net1069));
 sky130_fd_sc_hd__buf_4 wire1070 (.A(_2111_),
    .X(net1070));
 sky130_fd_sc_hd__clkbuf_8 wire1071 (.A(net1072),
    .X(net1071));
 sky130_fd_sc_hd__buf_4 wire1072 (.A(_2109_),
    .X(net1072));
 sky130_fd_sc_hd__buf_4 wire1073 (.A(net1074),
    .X(net1073));
 sky130_fd_sc_hd__buf_4 wire1074 (.A(_2107_),
    .X(net1074));
 sky130_fd_sc_hd__buf_4 wire1075 (.A(net1076),
    .X(net1075));
 sky130_fd_sc_hd__buf_6 wire1076 (.A(_2106_),
    .X(net1076));
 sky130_fd_sc_hd__buf_4 wire1077 (.A(_2104_),
    .X(net1077));
 sky130_fd_sc_hd__clkbuf_8 wire1078 (.A(net1079),
    .X(net1078));
 sky130_fd_sc_hd__buf_6 wire1079 (.A(_2102_),
    .X(net1079));
 sky130_fd_sc_hd__buf_4 wire1080 (.A(_2101_),
    .X(net1080));
 sky130_fd_sc_hd__clkbuf_8 wire1081 (.A(_2099_),
    .X(net1081));
 sky130_fd_sc_hd__buf_4 wire1082 (.A(net1083),
    .X(net1082));
 sky130_fd_sc_hd__buf_6 wire1083 (.A(_2097_),
    .X(net1083));
 sky130_fd_sc_hd__buf_4 wire1084 (.A(_2096_),
    .X(net1084));
 sky130_fd_sc_hd__buf_4 wire1085 (.A(_2094_),
    .X(net1085));
 sky130_fd_sc_hd__buf_6 wire1086 (.A(net1087),
    .X(net1086));
 sky130_fd_sc_hd__buf_6 wire1087 (.A(net1088),
    .X(net1087));
 sky130_fd_sc_hd__buf_4 wire1088 (.A(_2092_),
    .X(net1088));
 sky130_fd_sc_hd__buf_4 wire1089 (.A(_2091_),
    .X(net1089));
 sky130_fd_sc_hd__buf_6 wire1090 (.A(_2089_),
    .X(net1090));
 sky130_fd_sc_hd__buf_6 wire1091 (.A(_2087_),
    .X(net1091));
 sky130_fd_sc_hd__buf_12 wire1092 (.A(_2086_),
    .X(net1092));
 sky130_fd_sc_hd__buf_4 wire1093 (.A(_2084_),
    .X(net1093));
 sky130_fd_sc_hd__buf_4 wire1094 (.A(net1095),
    .X(net1094));
 sky130_fd_sc_hd__buf_6 wire1095 (.A(net1096),
    .X(net1095));
 sky130_fd_sc_hd__buf_6 wire1096 (.A(_2082_),
    .X(net1096));
 sky130_fd_sc_hd__buf_4 wire1098 (.A(_2079_),
    .X(net1098));
 sky130_fd_sc_hd__clkbuf_8 wire1099 (.A(net1100),
    .X(net1099));
 sky130_fd_sc_hd__buf_6 wire1100 (.A(_2077_),
    .X(net1100));
 sky130_fd_sc_hd__clkbuf_8 wire1102 (.A(_2074_),
    .X(net1102));
 sky130_fd_sc_hd__buf_4 wire1103 (.A(net1104),
    .X(net1103));
 sky130_fd_sc_hd__buf_6 wire1104 (.A(net1105),
    .X(net1104));
 sky130_fd_sc_hd__buf_4 wire1105 (.A(_2072_),
    .X(net1105));
 sky130_fd_sc_hd__buf_4 wire1106 (.A(net1107),
    .X(net1106));
 sky130_fd_sc_hd__buf_4 wire1107 (.A(_2069_),
    .X(net1107));
 sky130_fd_sc_hd__buf_6 wire1108 (.A(_2067_),
    .X(net1108));
 sky130_fd_sc_hd__buf_6 wire1109 (.A(net1110),
    .X(net1109));
 sky130_fd_sc_hd__buf_4 wire1110 (.A(_2066_),
    .X(net1110));
 sky130_fd_sc_hd__buf_4 wire1111 (.A(_2064_),
    .X(net1111));
 sky130_fd_sc_hd__buf_12 wire1112 (.A(net1113),
    .X(net1112));
 sky130_fd_sc_hd__buf_4 wire1113 (.A(_2062_),
    .X(net1113));
 sky130_fd_sc_hd__buf_6 wire1114 (.A(_2061_),
    .X(net1114));
 sky130_fd_sc_hd__buf_12 wire1115 (.A(_2059_),
    .X(net1115));
 sky130_fd_sc_hd__buf_4 wire1116 (.A(net1117),
    .X(net1116));
 sky130_fd_sc_hd__buf_6 wire1117 (.A(net1118),
    .X(net1117));
 sky130_fd_sc_hd__buf_4 wire1118 (.A(_2057_),
    .X(net1118));
 sky130_fd_sc_hd__buf_4 wire1120 (.A(net1121),
    .X(net1120));
 sky130_fd_sc_hd__buf_4 wire1121 (.A(_2054_),
    .X(net1121));
 sky130_fd_sc_hd__buf_8 wire1122 (.A(_2052_),
    .X(net1122));
 sky130_fd_sc_hd__buf_12 wire1123 (.A(net1124),
    .X(net1123));
 sky130_fd_sc_hd__buf_6 wire1124 (.A(_2051_),
    .X(net1124));
 sky130_fd_sc_hd__buf_6 wire1125 (.A(_2049_),
    .X(net1125));
 sky130_fd_sc_hd__buf_12 wire1126 (.A(net1127),
    .X(net1126));
 sky130_fd_sc_hd__buf_6 wire1127 (.A(_2047_),
    .X(net1127));
 sky130_fd_sc_hd__buf_8 wire1128 (.A(_2044_),
    .X(net1128));
 sky130_fd_sc_hd__buf_4 wire1129 (.A(net1130),
    .X(net1129));
 sky130_fd_sc_hd__buf_6 wire1130 (.A(_2042_),
    .X(net1130));
 sky130_fd_sc_hd__buf_4 wire1131 (.A(net1132),
    .X(net1131));
 sky130_fd_sc_hd__buf_6 wire1132 (.A(net1133),
    .X(net1132));
 sky130_fd_sc_hd__buf_4 wire1133 (.A(_2041_),
    .X(net1133));
 sky130_fd_sc_hd__buf_6 wire1134 (.A(_2039_),
    .X(net1134));
 sky130_fd_sc_hd__buf_12 wire1135 (.A(net1136),
    .X(net1135));
 sky130_fd_sc_hd__buf_6 wire1136 (.A(_2037_),
    .X(net1136));
 sky130_fd_sc_hd__buf_6 wire1137 (.A(_2034_),
    .X(net1137));
 sky130_fd_sc_hd__buf_4 wire1138 (.A(net1139),
    .X(net1138));
 sky130_fd_sc_hd__buf_4 wire1139 (.A(_2032_),
    .X(net1139));
 sky130_fd_sc_hd__buf_4 wire1140 (.A(net1141),
    .X(net1140));
 sky130_fd_sc_hd__buf_6 wire1141 (.A(_2031_),
    .X(net1141));
 sky130_fd_sc_hd__buf_4 wire1142 (.A(_2029_),
    .X(net1142));
 sky130_fd_sc_hd__buf_4 wire1181 (.A(_1911_),
    .X(net1181));
 sky130_fd_sc_hd__buf_4 wire1279 (.A(\u_dcg_s0.cfg_mode[1] ),
    .X(net1279));
 sky130_fd_sc_hd__buf_8 wire1280 (.A(\u_reg.reg_rdata[31] ),
    .X(net1280));
 sky130_fd_sc_hd__buf_4 wire1281 (.A(\u_reg.reg_rdata[30] ),
    .X(net1281));
 sky130_fd_sc_hd__buf_4 wire1282 (.A(net1283),
    .X(net1282));
 sky130_fd_sc_hd__buf_4 wire1283 (.A(\u_reg.reg_rdata[29] ),
    .X(net1283));
 sky130_fd_sc_hd__buf_4 wire1284 (.A(\u_reg.reg_rdata[28] ),
    .X(net1284));
 sky130_fd_sc_hd__buf_4 wire1285 (.A(\u_reg.reg_rdata[27] ),
    .X(net1285));
 sky130_fd_sc_hd__buf_4 wire1286 (.A(net1287),
    .X(net1286));
 sky130_fd_sc_hd__buf_6 wire1287 (.A(\u_reg.reg_rdata[26] ),
    .X(net1287));
 sky130_fd_sc_hd__buf_4 wire1288 (.A(\u_reg.reg_rdata[25] ),
    .X(net1288));
 sky130_fd_sc_hd__buf_6 wire1289 (.A(\u_reg.reg_rdata[24] ),
    .X(net1289));
 sky130_fd_sc_hd__buf_4 wire1290 (.A(\u_reg.reg_rdata[22] ),
    .X(net1290));
 sky130_fd_sc_hd__buf_4 wire1291 (.A(net1292),
    .X(net1291));
 sky130_fd_sc_hd__buf_4 wire1292 (.A(\u_reg.reg_rdata[21] ),
    .X(net1292));
 sky130_fd_sc_hd__buf_4 wire1293 (.A(net1294),
    .X(net1293));
 sky130_fd_sc_hd__buf_6 wire1294 (.A(\u_reg.reg_rdata[20] ),
    .X(net1294));
 sky130_fd_sc_hd__buf_8 wire1295 (.A(\u_reg.reg_rdata[17] ),
    .X(net1295));
 sky130_fd_sc_hd__clkbuf_8 wire1296 (.A(net1297),
    .X(net1296));
 sky130_fd_sc_hd__buf_6 wire1297 (.A(\u_reg.reg_rdata[16] ),
    .X(net1297));
 sky130_fd_sc_hd__buf_4 wire1298 (.A(net1299),
    .X(net1298));
 sky130_fd_sc_hd__buf_4 wire1299 (.A(\u_reg.reg_rdata[15] ),
    .X(net1299));
 sky130_fd_sc_hd__buf_4 wire13 (.A(\clknet_3_1__leaf_u_dsync.out_clk ),
    .X(net1745));
 sky130_fd_sc_hd__clkbuf_8 wire1300 (.A(net1301),
    .X(net1300));
 sky130_fd_sc_hd__buf_4 wire1301 (.A(\u_reg.reg_rdata[14] ),
    .X(net1301));
 sky130_fd_sc_hd__buf_4 wire1302 (.A(net1303),
    .X(net1302));
 sky130_fd_sc_hd__buf_4 wire1303 (.A(\u_reg.reg_rdata[13] ),
    .X(net1303));
 sky130_fd_sc_hd__buf_6 wire1304 (.A(\u_reg.reg_rdata[12] ),
    .X(net1304));
 sky130_fd_sc_hd__buf_6 wire1305 (.A(\u_reg.reg_rdata[11] ),
    .X(net1305));
 sky130_fd_sc_hd__buf_4 wire1306 (.A(\u_reg.reg_rdata[10] ),
    .X(net1306));
 sky130_fd_sc_hd__clkbuf_8 wire1307 (.A(\u_reg.reg_rdata[9] ),
    .X(net1307));
 sky130_fd_sc_hd__buf_4 wire1308 (.A(\u_reg.reg_rdata[8] ),
    .X(net1308));
 sky130_fd_sc_hd__clkbuf_8 wire1309 (.A(\u_reg.reg_rdata[7] ),
    .X(net1309));
 sky130_fd_sc_hd__buf_4 wire1310 (.A(\u_reg.reg_rdata[5] ),
    .X(net1310));
 sky130_fd_sc_hd__buf_6 wire1311 (.A(\u_reg.reg_rdata[4] ),
    .X(net1311));
 sky130_fd_sc_hd__buf_4 wire1312 (.A(\u_reg.reg_rdata[0] ),
    .X(net1312));
 sky130_fd_sc_hd__buf_4 wire1366 (.A(\u_s1.u_sync_wbb.wbm_lack_o ),
    .X(net1366));
 sky130_fd_sc_hd__buf_6 wire1367 (.A(\u_s1.u_sync_wbb.wbm_ack_o ),
    .X(net1367));
 sky130_fd_sc_hd__buf_6 wire1401 (.A(net1400),
    .X(net1401));
 sky130_fd_sc_hd__buf_12 wire1402 (.A(net1403),
    .X(net1402));
 sky130_fd_sc_hd__buf_6 wire1411 (.A(net1412),
    .X(net1411));
 sky130_fd_sc_hd__buf_4 wire1412 (.A(\u_dcg_peri.clk_enb ),
    .X(net1412));
 sky130_fd_sc_hd__buf_6 wire1413 (.A(net1414),
    .X(net1413));
 sky130_fd_sc_hd__buf_4 wire1414 (.A(\u_dcg_riscv.clk_enb ),
    .X(net1414));
 sky130_fd_sc_hd__buf_4 wire1415 (.A(\u_dcg_s2.clk_enb ),
    .X(net1415));
 sky130_fd_sc_hd__buf_6 wire1416 (.A(net1417),
    .X(net1416));
 sky130_fd_sc_hd__buf_6 wire1417 (.A(net1418),
    .X(net1417));
 sky130_fd_sc_hd__buf_6 wire1418 (.A(net64),
    .X(net1418));
 sky130_fd_sc_hd__buf_6 wire1419 (.A(net1420),
    .X(net1419));
 sky130_fd_sc_hd__buf_6 wire1420 (.A(net1421),
    .X(net1420));
 sky130_fd_sc_hd__buf_6 wire1421 (.A(net63),
    .X(net1421));
 sky130_fd_sc_hd__buf_6 wire1422 (.A(net1423),
    .X(net1422));
 sky130_fd_sc_hd__buf_6 wire1423 (.A(net1424),
    .X(net1423));
 sky130_fd_sc_hd__buf_6 wire1424 (.A(net62),
    .X(net1424));
 sky130_fd_sc_hd__buf_6 wire1425 (.A(net1426),
    .X(net1425));
 sky130_fd_sc_hd__buf_6 wire1426 (.A(net1427),
    .X(net1426));
 sky130_fd_sc_hd__buf_6 wire1427 (.A(net58),
    .X(net1427));
 sky130_fd_sc_hd__buf_6 wire1428 (.A(net1429),
    .X(net1428));
 sky130_fd_sc_hd__buf_6 wire1429 (.A(net1430),
    .X(net1429));
 sky130_fd_sc_hd__buf_6 wire1430 (.A(net57),
    .X(net1430));
 sky130_fd_sc_hd__buf_6 wire1431 (.A(net1432),
    .X(net1431));
 sky130_fd_sc_hd__buf_6 wire1432 (.A(net1433),
    .X(net1432));
 sky130_fd_sc_hd__buf_6 wire1433 (.A(net56),
    .X(net1433));
 sky130_fd_sc_hd__buf_6 wire1434 (.A(net1435),
    .X(net1434));
 sky130_fd_sc_hd__buf_6 wire1435 (.A(net1436),
    .X(net1435));
 sky130_fd_sc_hd__buf_6 wire1436 (.A(net55),
    .X(net1436));
 sky130_fd_sc_hd__buf_4 wire1437 (.A(net54),
    .X(net1437));
 sky130_fd_sc_hd__buf_6 wire1438 (.A(net53),
    .X(net1438));
 sky130_fd_sc_hd__buf_4 wire1439 (.A(net52),
    .X(net1439));
 sky130_fd_sc_hd__buf_4 wire1440 (.A(net51),
    .X(net1440));
 sky130_fd_sc_hd__buf_4 wire1441 (.A(net50),
    .X(net1441));
 sky130_fd_sc_hd__buf_4 wire1442 (.A(net49),
    .X(net1442));
 sky130_fd_sc_hd__buf_4 wire1443 (.A(net47),
    .X(net1443));
 sky130_fd_sc_hd__buf_4 wire1444 (.A(net46),
    .X(net1444));
 sky130_fd_sc_hd__buf_6 wire1445 (.A(net45),
    .X(net1445));
 sky130_fd_sc_hd__buf_6 wire1446 (.A(net44),
    .X(net1446));
 sky130_fd_sc_hd__buf_6 wire1447 (.A(net43),
    .X(net1447));
 sky130_fd_sc_hd__buf_6 wire1448 (.A(net42),
    .X(net1448));
 sky130_fd_sc_hd__buf_6 wire1449 (.A(net41),
    .X(net1449));
 sky130_fd_sc_hd__buf_6 wire1450 (.A(net40),
    .X(net1450));
 sky130_fd_sc_hd__buf_6 wire1451 (.A(net1452),
    .X(net1451));
 sky130_fd_sc_hd__buf_4 wire1452 (.A(net39),
    .X(net1452));
 sky130_fd_sc_hd__buf_6 wire1453 (.A(net1454),
    .X(net1453));
 sky130_fd_sc_hd__buf_4 wire1454 (.A(net38),
    .X(net1454));
 sky130_fd_sc_hd__buf_6 wire1455 (.A(net1456),
    .X(net1455));
 sky130_fd_sc_hd__buf_4 wire1456 (.A(net36),
    .X(net1456));
 sky130_fd_sc_hd__buf_6 wire1457 (.A(net1458),
    .X(net1457));
 sky130_fd_sc_hd__buf_4 wire1458 (.A(net35),
    .X(net1458));
 sky130_fd_sc_hd__buf_6 wire1459 (.A(net1460),
    .X(net1459));
 sky130_fd_sc_hd__buf_4 wire1460 (.A(net34),
    .X(net1460));
 sky130_fd_sc_hd__buf_6 wire1461 (.A(net1462),
    .X(net1461));
 sky130_fd_sc_hd__buf_4 wire1462 (.A(net33),
    .X(net1462));
 sky130_fd_sc_hd__buf_6 wire1463 (.A(net1464),
    .X(net1463));
 sky130_fd_sc_hd__buf_4 wire1464 (.A(net32),
    .X(net1464));
 sky130_fd_sc_hd__buf_6 wire1465 (.A(net1466),
    .X(net1465));
 sky130_fd_sc_hd__buf_4 wire1466 (.A(net31),
    .X(net1466));
 sky130_fd_sc_hd__buf_6 wire1467 (.A(net1468),
    .X(net1467));
 sky130_fd_sc_hd__buf_4 wire1468 (.A(net30),
    .X(net1468));
 sky130_fd_sc_hd__buf_6 wire1469 (.A(net1470),
    .X(net1469));
 sky130_fd_sc_hd__buf_4 wire1470 (.A(net29),
    .X(net1470));
 sky130_fd_sc_hd__buf_6 wire1471 (.A(net1472),
    .X(net1471));
 sky130_fd_sc_hd__buf_4 wire1472 (.A(net28),
    .X(net1472));
 sky130_fd_sc_hd__buf_6 wire1473 (.A(net1474),
    .X(net1473));
 sky130_fd_sc_hd__buf_4 wire1474 (.A(net27),
    .X(net1474));
 sky130_fd_sc_hd__buf_6 wire1475 (.A(net1476),
    .X(net1475));
 sky130_fd_sc_hd__buf_4 wire1476 (.A(net25),
    .X(net1476));
 sky130_fd_sc_hd__buf_6 wire1477 (.A(net1478),
    .X(net1477));
 sky130_fd_sc_hd__buf_4 wire1478 (.A(net24),
    .X(net1478));
 sky130_fd_sc_hd__buf_6 wire1479 (.A(net1480),
    .X(net1479));
 sky130_fd_sc_hd__buf_6 wire1480 (.A(net23),
    .X(net1480));
 sky130_fd_sc_hd__buf_6 wire1481 (.A(net1482),
    .X(net1481));
 sky130_fd_sc_hd__buf_6 wire1482 (.A(net22),
    .X(net1482));
 sky130_fd_sc_hd__buf_6 wire1483 (.A(net1484),
    .X(net1483));
 sky130_fd_sc_hd__buf_4 wire1484 (.A(net21),
    .X(net1484));
 sky130_fd_sc_hd__buf_6 wire1485 (.A(net1486),
    .X(net1485));
 sky130_fd_sc_hd__buf_6 wire1486 (.A(net20),
    .X(net1486));
 sky130_fd_sc_hd__buf_6 wire1487 (.A(net1488),
    .X(net1487));
 sky130_fd_sc_hd__buf_4 wire1488 (.A(net19),
    .X(net1488));
 sky130_fd_sc_hd__buf_6 wire1489 (.A(net1490),
    .X(net1489));
 sky130_fd_sc_hd__buf_4 wire1490 (.A(net18),
    .X(net1490));
 sky130_fd_sc_hd__buf_4 wire1491 (.A(net26),
    .X(net1491));
 sky130_fd_sc_hd__buf_4 wire1492 (.A(\u_dcg_riscv.cfg_mode_ss[1] ),
    .X(net1492));
 sky130_fd_sc_hd__buf_4 wire1493 (.A(net2081),
    .X(net1493));
 sky130_fd_sc_hd__buf_4 wire1494 (.A(net2070),
    .X(net1494));
 sky130_fd_sc_hd__buf_6 wire1511 (.A(net1512),
    .X(net1511));
 sky130_fd_sc_hd__buf_4 wire1512 (.A(s0_idle),
    .X(net1512));
 sky130_fd_sc_hd__buf_6 wire1513 (.A(m2_wbd_dat_i[9]),
    .X(net1513));
 sky130_fd_sc_hd__buf_4 wire1514 (.A(m2_wbd_dat_i[8]),
    .X(net1514));
 sky130_fd_sc_hd__buf_4 wire1515 (.A(m2_wbd_dat_i[7]),
    .X(net1515));
 sky130_fd_sc_hd__buf_6 wire1516 (.A(m2_wbd_dat_i[6]),
    .X(net1516));
 sky130_fd_sc_hd__buf_6 wire1517 (.A(m2_wbd_dat_i[5]),
    .X(net1517));
 sky130_fd_sc_hd__buf_4 wire1519 (.A(m2_wbd_dat_i[31]),
    .X(net1519));
 sky130_fd_sc_hd__buf_4 wire1520 (.A(net1964),
    .X(net1520));
 sky130_fd_sc_hd__buf_4 wire1522 (.A(net2041),
    .X(net1522));
 sky130_fd_sc_hd__buf_4 wire1523 (.A(net1955),
    .X(net1523));
 sky130_fd_sc_hd__buf_4 wire1524 (.A(m2_wbd_dat_i[23]),
    .X(net1524));
 sky130_fd_sc_hd__buf_4 wire1525 (.A(m2_wbd_dat_i[21]),
    .X(net1525));
 sky130_fd_sc_hd__buf_4 wire1526 (.A(net1950),
    .X(net1526));
 sky130_fd_sc_hd__buf_4 wire1527 (.A(net2054),
    .X(net1527));
 sky130_fd_sc_hd__buf_6 wire1528 (.A(net2019),
    .X(net1528));
 sky130_fd_sc_hd__buf_4 wire1529 (.A(net2076),
    .X(net1529));
 sky130_fd_sc_hd__buf_4 wire1531 (.A(net2072),
    .X(net1531));
 sky130_fd_sc_hd__buf_4 wire1532 (.A(m2_wbd_dat_i[12]),
    .X(net1532));
 sky130_fd_sc_hd__buf_6 wire1533 (.A(net1947),
    .X(net1533));
 sky130_fd_sc_hd__buf_6 wire1534 (.A(m2_wbd_dat_i[10]),
    .X(net1534));
 sky130_fd_sc_hd__buf_8 wire1535 (.A(m1_wbd_dat_i[9]),
    .X(net1535));
 sky130_fd_sc_hd__buf_4 wire1536 (.A(m1_wbd_dat_i[8]),
    .X(net1536));
 sky130_fd_sc_hd__buf_4 wire1537 (.A(m1_wbd_dat_i[7]),
    .X(net1537));
 sky130_fd_sc_hd__buf_8 wire1538 (.A(m1_wbd_dat_i[6]),
    .X(net1538));
 sky130_fd_sc_hd__buf_8 wire1539 (.A(m1_wbd_dat_i[5]),
    .X(net1539));
 sky130_fd_sc_hd__buf_4 wire1540 (.A(m1_wbd_dat_i[4]),
    .X(net1540));
 sky130_fd_sc_hd__buf_6 wire1541 (.A(m1_wbd_dat_i[31]),
    .X(net1541));
 sky130_fd_sc_hd__buf_6 wire1542 (.A(net2071),
    .X(net1542));
 sky130_fd_sc_hd__buf_6 wire1543 (.A(net2052),
    .X(net1543));
 sky130_fd_sc_hd__buf_4 wire1544 (.A(net2023),
    .X(net1544));
 sky130_fd_sc_hd__buf_6 wire1545 (.A(net1945),
    .X(net1545));
 sky130_fd_sc_hd__buf_4 wire1546 (.A(m1_wbd_dat_i[26]),
    .X(net1546));
 sky130_fd_sc_hd__buf_6 wire1547 (.A(m1_wbd_dat_i[23]),
    .X(net1547));
 sky130_fd_sc_hd__buf_6 wire1548 (.A(m1_wbd_dat_i[22]),
    .X(net1548));
 sky130_fd_sc_hd__buf_6 wire1549 (.A(m1_wbd_dat_i[21]),
    .X(net1549));
 sky130_fd_sc_hd__buf_4 wire1550 (.A(net2064),
    .X(net1550));
 sky130_fd_sc_hd__buf_4 wire1551 (.A(m1_wbd_dat_i[1]),
    .X(net1551));
 sky130_fd_sc_hd__buf_4 wire1552 (.A(net2008),
    .X(net1552));
 sky130_fd_sc_hd__buf_6 wire1553 (.A(m1_wbd_dat_i[18]),
    .X(net1553));
 sky130_fd_sc_hd__buf_6 wire1554 (.A(net1949),
    .X(net1554));
 sky130_fd_sc_hd__buf_4 wire1555 (.A(m1_wbd_dat_i[16]),
    .X(net1555));
 sky130_fd_sc_hd__buf_6 wire1556 (.A(m1_wbd_dat_i[15]),
    .X(net1556));
 sky130_fd_sc_hd__buf_6 wire1557 (.A(m1_wbd_dat_i[14]),
    .X(net1557));
 sky130_fd_sc_hd__buf_6 wire1558 (.A(m1_wbd_dat_i[13]),
    .X(net1558));
 sky130_fd_sc_hd__buf_6 wire1559 (.A(m1_wbd_dat_i[12]),
    .X(net1559));
 sky130_fd_sc_hd__buf_6 wire1560 (.A(m1_wbd_dat_i[11]),
    .X(net1560));
 sky130_fd_sc_hd__buf_6 wire1561 (.A(net2068),
    .X(net1561));
 sky130_fd_sc_hd__buf_4 wire1562 (.A(m1_wbd_dat_i[0]),
    .X(net1562));
 sky130_fd_sc_hd__buf_4 wire1563 (.A(m1_wbd_bry_i),
    .X(net1563));
 sky130_fd_sc_hd__buf_4 wire1564 (.A(m1_wbd_bl_i[0]),
    .X(net1564));
 sky130_fd_sc_hd__buf_4 wire1565 (.A(m0_wbd_sel_i[0]),
    .X(net1565));
 sky130_fd_sc_hd__buf_8 wire1566 (.A(m0_wbd_dat_i[9]),
    .X(net1566));
 sky130_fd_sc_hd__buf_4 wire1567 (.A(m0_wbd_dat_i[8]),
    .X(net1567));
 sky130_fd_sc_hd__clkbuf_8 wire1568 (.A(net1967),
    .X(net1568));
 sky130_fd_sc_hd__buf_6 wire1569 (.A(m0_wbd_dat_i[6]),
    .X(net1569));
 sky130_fd_sc_hd__buf_8 wire1570 (.A(m0_wbd_dat_i[5]),
    .X(net1570));
 sky130_fd_sc_hd__buf_4 wire1571 (.A(net2062),
    .X(net1571));
 sky130_fd_sc_hd__buf_4 wire1572 (.A(m0_wbd_dat_i[31]),
    .X(net1572));
 sky130_fd_sc_hd__buf_6 wire1573 (.A(net1985),
    .X(net1573));
 sky130_fd_sc_hd__buf_6 wire1574 (.A(m0_wbd_dat_i[2]),
    .X(net1574));
 sky130_fd_sc_hd__buf_6 wire1575 (.A(net2028),
    .X(net1575));
 sky130_fd_sc_hd__buf_6 wire1576 (.A(net2010),
    .X(net1576));
 sky130_fd_sc_hd__buf_4 wire1577 (.A(net2018),
    .X(net1577));
 sky130_fd_sc_hd__buf_6 wire1578 (.A(m0_wbd_dat_i[23]),
    .X(net1578));
 sky130_fd_sc_hd__buf_6 wire1579 (.A(m0_wbd_dat_i[22]),
    .X(net1579));
 sky130_fd_sc_hd__buf_6 wire1580 (.A(m0_wbd_dat_i[21]),
    .X(net1580));
 sky130_fd_sc_hd__buf_4 wire1581 (.A(net2075),
    .X(net1581));
 sky130_fd_sc_hd__buf_4 wire1582 (.A(m0_wbd_dat_i[1]),
    .X(net1582));
 sky130_fd_sc_hd__buf_6 wire1583 (.A(net1976),
    .X(net1583));
 sky130_fd_sc_hd__buf_4 wire1584 (.A(m0_wbd_dat_i[18]),
    .X(net1584));
 sky130_fd_sc_hd__buf_6 wire1585 (.A(m0_wbd_dat_i[17]),
    .X(net1585));
 sky130_fd_sc_hd__buf_4 wire1586 (.A(m0_wbd_dat_i[16]),
    .X(net1586));
 sky130_fd_sc_hd__buf_6 wire1587 (.A(m0_wbd_dat_i[15]),
    .X(net1587));
 sky130_fd_sc_hd__buf_6 wire1588 (.A(m0_wbd_dat_i[14]),
    .X(net1588));
 sky130_fd_sc_hd__buf_6 wire1589 (.A(m0_wbd_dat_i[13]),
    .X(net1589));
 sky130_fd_sc_hd__buf_6 wire1590 (.A(m0_wbd_dat_i[12]),
    .X(net1590));
 sky130_fd_sc_hd__buf_6 wire1591 (.A(m0_wbd_dat_i[11]),
    .X(net1591));
 sky130_fd_sc_hd__buf_6 wire1592 (.A(m0_wbd_dat_i[10]),
    .X(net1592));
 sky130_fd_sc_hd__buf_6 wire1593 (.A(m0_wbd_dat_i[0]),
    .X(net1593));
 sky130_fd_sc_hd__buf_4 wire1594 (.A(m0_wbd_adr_i[7]),
    .X(net1594));
 sky130_fd_sc_hd__buf_4 wire1595 (.A(m0_wbd_adr_i[5]),
    .X(net1595));
 sky130_fd_sc_hd__buf_6 wire1596 (.A(m0_wbd_adr_i[4]),
    .X(net1596));
 sky130_fd_sc_hd__buf_6 wire1597 (.A(net2093),
    .X(net1597));
 sky130_fd_sc_hd__buf_4 wire1598 (.A(m0_wbd_adr_i[2]),
    .X(net1598));
 sky130_fd_sc_hd__buf_6 wire1599 (.A(ch_data_in[99]),
    .X(net1599));
 sky130_fd_sc_hd__buf_6 wire1600 (.A(ch_data_in[98]),
    .X(net1600));
 sky130_fd_sc_hd__buf_6 wire1601 (.A(net1602),
    .X(net1601));
 sky130_fd_sc_hd__buf_4 wire1602 (.A(ch_data_in[97]),
    .X(net1602));
 sky130_fd_sc_hd__buf_6 wire1603 (.A(net1604),
    .X(net1603));
 sky130_fd_sc_hd__buf_4 wire1604 (.A(ch_data_in[96]),
    .X(net1604));
 sky130_fd_sc_hd__buf_6 wire1605 (.A(net1606),
    .X(net1605));
 sky130_fd_sc_hd__buf_4 wire1606 (.A(ch_data_in[95]),
    .X(net1606));
 sky130_fd_sc_hd__buf_6 wire1607 (.A(net1608),
    .X(net1607));
 sky130_fd_sc_hd__buf_4 wire1608 (.A(ch_data_in[94]),
    .X(net1608));
 sky130_fd_sc_hd__buf_6 wire1609 (.A(net1610),
    .X(net1609));
 sky130_fd_sc_hd__buf_4 wire1610 (.A(ch_data_in[93]),
    .X(net1610));
 sky130_fd_sc_hd__buf_6 wire1611 (.A(net1612),
    .X(net1611));
 sky130_fd_sc_hd__buf_4 wire1612 (.A(ch_data_in[92]),
    .X(net1612));
 sky130_fd_sc_hd__buf_6 wire1613 (.A(net1614),
    .X(net1613));
 sky130_fd_sc_hd__buf_6 wire1614 (.A(ch_data_in[91]),
    .X(net1614));
 sky130_fd_sc_hd__buf_6 wire1615 (.A(net1616),
    .X(net1615));
 sky130_fd_sc_hd__buf_4 wire1616 (.A(ch_data_in[90]),
    .X(net1616));
 sky130_fd_sc_hd__buf_6 wire1617 (.A(net1618),
    .X(net1617));
 sky130_fd_sc_hd__buf_6 wire1618 (.A(ch_data_in[89]),
    .X(net1618));
 sky130_fd_sc_hd__buf_6 wire1619 (.A(net1620),
    .X(net1619));
 sky130_fd_sc_hd__buf_4 wire1620 (.A(ch_data_in[88]),
    .X(net1620));
 sky130_fd_sc_hd__buf_6 wire1621 (.A(net1622),
    .X(net1621));
 sky130_fd_sc_hd__buf_4 wire1622 (.A(ch_data_in[87]),
    .X(net1622));
 sky130_fd_sc_hd__buf_6 wire1623 (.A(net1624),
    .X(net1623));
 sky130_fd_sc_hd__buf_4 wire1624 (.A(ch_data_in[86]),
    .X(net1624));
 sky130_fd_sc_hd__buf_6 wire1625 (.A(net1626),
    .X(net1625));
 sky130_fd_sc_hd__buf_4 wire1626 (.A(ch_data_in[85]),
    .X(net1626));
 sky130_fd_sc_hd__buf_6 wire1627 (.A(net1628),
    .X(net1627));
 sky130_fd_sc_hd__buf_6 wire1628 (.A(ch_data_in[84]),
    .X(net1628));
 sky130_fd_sc_hd__buf_6 wire1629 (.A(net1630),
    .X(net1629));
 sky130_fd_sc_hd__buf_6 wire1630 (.A(ch_data_in[83]),
    .X(net1630));
 sky130_fd_sc_hd__buf_6 wire1631 (.A(net1632),
    .X(net1631));
 sky130_fd_sc_hd__buf_6 wire1632 (.A(ch_data_in[82]),
    .X(net1632));
 sky130_fd_sc_hd__buf_6 wire1633 (.A(net1634),
    .X(net1633));
 sky130_fd_sc_hd__buf_6 wire1634 (.A(ch_data_in[81]),
    .X(net1634));
 sky130_fd_sc_hd__buf_6 wire1635 (.A(net1636),
    .X(net1635));
 sky130_fd_sc_hd__buf_6 wire1636 (.A(ch_data_in[80]),
    .X(net1636));
 sky130_fd_sc_hd__buf_6 wire1637 (.A(net1638),
    .X(net1637));
 sky130_fd_sc_hd__buf_6 wire1638 (.A(ch_data_in[79]),
    .X(net1638));
 sky130_fd_sc_hd__buf_6 wire1639 (.A(net1640),
    .X(net1639));
 sky130_fd_sc_hd__buf_6 wire1640 (.A(ch_data_in[78]),
    .X(net1640));
 sky130_fd_sc_hd__buf_6 wire1641 (.A(net1642),
    .X(net1641));
 sky130_fd_sc_hd__buf_6 wire1642 (.A(ch_data_in[77]),
    .X(net1642));
 sky130_fd_sc_hd__buf_4 wire1643 (.A(ch_data_in[43]),
    .X(net1643));
 sky130_fd_sc_hd__buf_4 wire1644 (.A(ch_data_in[42]),
    .X(net1644));
 sky130_fd_sc_hd__buf_4 wire1645 (.A(ch_data_in[41]),
    .X(net1645));
 sky130_fd_sc_hd__buf_4 wire1646 (.A(ch_data_in[40]),
    .X(net1646));
 sky130_fd_sc_hd__buf_4 wire1647 (.A(ch_data_in[39]),
    .X(net1647));
 sky130_fd_sc_hd__buf_4 wire1648 (.A(ch_data_in[38]),
    .X(net1648));
 sky130_fd_sc_hd__buf_4 wire1649 (.A(ch_data_in[37]),
    .X(net1649));
 sky130_fd_sc_hd__buf_4 wire1650 (.A(ch_data_in[36]),
    .X(net1650));
 sky130_fd_sc_hd__buf_4 wire1651 (.A(ch_data_in[35]),
    .X(net1651));
 sky130_fd_sc_hd__buf_4 wire1652 (.A(ch_data_in[34]),
    .X(net1652));
 sky130_fd_sc_hd__buf_4 wire1653 (.A(ch_data_in[33]),
    .X(net1653));
 sky130_fd_sc_hd__buf_4 wire1654 (.A(ch_data_in[32]),
    .X(net1654));
 sky130_fd_sc_hd__buf_4 wire1655 (.A(ch_data_in[31]),
    .X(net1655));
 sky130_fd_sc_hd__buf_4 wire1656 (.A(ch_data_in[30]),
    .X(net1656));
 sky130_fd_sc_hd__buf_4 wire1657 (.A(ch_data_in[29]),
    .X(net1657));
 sky130_fd_sc_hd__buf_4 wire1658 (.A(ch_data_in[28]),
    .X(net1658));
 sky130_fd_sc_hd__buf_6 wire1659 (.A(ch_data_in[27]),
    .X(net1659));
 sky130_fd_sc_hd__buf_6 wire1660 (.A(ch_data_in[26]),
    .X(net1660));
 sky130_fd_sc_hd__buf_6 wire1661 (.A(ch_data_in[25]),
    .X(net1661));
 sky130_fd_sc_hd__buf_6 wire1662 (.A(ch_data_in[24]),
    .X(net1662));
 sky130_fd_sc_hd__buf_6 wire1663 (.A(net1664),
    .X(net1663));
 sky130_fd_sc_hd__buf_6 wire1664 (.A(ch_data_in[15]),
    .X(net1664));
 sky130_fd_sc_hd__buf_6 wire1665 (.A(net1666),
    .X(net1665));
 sky130_fd_sc_hd__buf_6 wire1666 (.A(net1667),
    .X(net1666));
 sky130_fd_sc_hd__buf_6 wire1667 (.A(ch_data_in[157]),
    .X(net1667));
 sky130_fd_sc_hd__buf_6 wire1668 (.A(net1669),
    .X(net1668));
 sky130_fd_sc_hd__buf_6 wire1669 (.A(net1670),
    .X(net1669));
 sky130_fd_sc_hd__buf_6 wire1670 (.A(ch_data_in[156]),
    .X(net1670));
 sky130_fd_sc_hd__buf_6 wire1671 (.A(net1672),
    .X(net1671));
 sky130_fd_sc_hd__buf_6 wire1672 (.A(net1673),
    .X(net1672));
 sky130_fd_sc_hd__buf_6 wire1673 (.A(ch_data_in[155]),
    .X(net1673));
 sky130_fd_sc_hd__buf_6 wire1674 (.A(net1675),
    .X(net1674));
 sky130_fd_sc_hd__buf_6 wire1675 (.A(net1676),
    .X(net1675));
 sky130_fd_sc_hd__buf_4 wire1676 (.A(ch_data_in[151]),
    .X(net1676));
 sky130_fd_sc_hd__buf_6 wire1677 (.A(net1678),
    .X(net1677));
 sky130_fd_sc_hd__buf_6 wire1678 (.A(net1679),
    .X(net1678));
 sky130_fd_sc_hd__buf_4 wire1679 (.A(ch_data_in[150]),
    .X(net1679));
 sky130_fd_sc_hd__buf_6 wire1680 (.A(net1681),
    .X(net1680));
 sky130_fd_sc_hd__buf_6 wire1681 (.A(ch_data_in[14]),
    .X(net1681));
 sky130_fd_sc_hd__clkbuf_4 wire1682 (.A(ch_data_in[143]),
    .X(net1682));
 sky130_fd_sc_hd__buf_4 wire1683 (.A(ch_data_in[142]),
    .X(net1683));
 sky130_fd_sc_hd__buf_4 wire1684 (.A(ch_data_in[141]),
    .X(net1684));
 sky130_fd_sc_hd__buf_4 wire1685 (.A(ch_data_in[140]),
    .X(net1685));
 sky130_fd_sc_hd__buf_6 wire1686 (.A(net1687),
    .X(net1686));
 sky130_fd_sc_hd__buf_6 wire1687 (.A(ch_data_in[13]),
    .X(net1687));
 sky130_fd_sc_hd__clkbuf_4 wire1688 (.A(ch_data_in[139]),
    .X(net1688));
 sky130_fd_sc_hd__buf_6 wire1689 (.A(net1690),
    .X(net1689));
 sky130_fd_sc_hd__buf_6 wire1690 (.A(ch_data_in[12]),
    .X(net1690));
 sky130_fd_sc_hd__buf_6 wire1691 (.A(net1692),
    .X(net1691));
 sky130_fd_sc_hd__buf_4 wire1692 (.A(ch_data_in[111]),
    .X(net1692));
 sky130_fd_sc_hd__buf_6 wire1693 (.A(net1694),
    .X(net1693));
 sky130_fd_sc_hd__buf_6 wire1694 (.A(ch_data_in[110]),
    .X(net1694));
 sky130_fd_sc_hd__buf_6 wire1695 (.A(net1696),
    .X(net1695));
 sky130_fd_sc_hd__buf_6 wire1696 (.A(ch_data_in[109]),
    .X(net1696));
 sky130_fd_sc_hd__buf_6 wire1697 (.A(net1698),
    .X(net1697));
 sky130_fd_sc_hd__buf_6 wire1698 (.A(ch_data_in[108]),
    .X(net1698));
 sky130_fd_sc_hd__buf_6 wire1699 (.A(net1700),
    .X(net1699));
 sky130_fd_sc_hd__buf_4 wire1700 (.A(ch_data_in[107]),
    .X(net1700));
 sky130_fd_sc_hd__buf_6 wire1701 (.A(net1702),
    .X(net1701));
 sky130_fd_sc_hd__buf_6 wire1702 (.A(ch_data_in[106]),
    .X(net1702));
 sky130_fd_sc_hd__buf_6 wire1703 (.A(net1704),
    .X(net1703));
 sky130_fd_sc_hd__buf_6 wire1704 (.A(ch_data_in[105]),
    .X(net1704));
 sky130_fd_sc_hd__buf_6 wire1705 (.A(net1706),
    .X(net1705));
 sky130_fd_sc_hd__buf_6 wire1706 (.A(ch_data_in[104]),
    .X(net1706));
 sky130_fd_sc_hd__buf_6 wire1707 (.A(net1708),
    .X(net1707));
 sky130_fd_sc_hd__buf_6 wire1708 (.A(ch_data_in[103]),
    .X(net1708));
 sky130_fd_sc_hd__buf_6 wire1709 (.A(net1710),
    .X(net1709));
 sky130_fd_sc_hd__buf_4 wire1710 (.A(ch_data_in[102]),
    .X(net1710));
 sky130_fd_sc_hd__buf_6 wire1711 (.A(net1712),
    .X(net1711));
 sky130_fd_sc_hd__buf_4 wire1712 (.A(ch_data_in[101]),
    .X(net1712));
 sky130_fd_sc_hd__buf_6 wire1713 (.A(net1714),
    .X(net1713));
 sky130_fd_sc_hd__buf_4 wire1714 (.A(ch_data_in[100]),
    .X(net1714));
 sky130_fd_sc_hd__buf_6 wire1715 (.A(ch_clk_in[2]),
    .X(net1715));
 sky130_fd_sc_hd__buf_4 wire1716 (.A(ch_clk_in[1]),
    .X(net1716));
 sky130_fd_sc_hd__buf_4 wire2 (.A(net1735),
    .X(net1734));
 sky130_fd_sc_hd__buf_4 wire21 (.A(net1754),
    .X(net1753));
 sky130_fd_sc_hd__buf_4 wire23 (.A(net1758),
    .X(net1755));
 sky130_fd_sc_hd__buf_4 wire24 (.A(net1757),
    .X(net1756));
 sky130_fd_sc_hd__clkbuf_8 wire25 (.A(\clknet_3_5__leaf_u_dsync.out_clk ),
    .X(net1757));
 sky130_fd_sc_hd__buf_4 wire27 (.A(\clknet_3_7__leaf_u_dsync.out_clk ),
    .X(net1759));
 sky130_fd_sc_hd__clkbuf_4 wire28 (.A(\clknet_3_7__leaf_u_dsync.out_clk ),
    .X(net1760));
 sky130_fd_sc_hd__buf_6 wire29 (.A(net1762),
    .X(net1761));
 sky130_fd_sc_hd__clkbuf_2 wire3 (.A(\u_dsync.out_clk ),
    .X(net1735));
 sky130_fd_sc_hd__buf_4 wire30 (.A(net1763),
    .X(net1762));
 sky130_fd_sc_hd__clkbuf_2 wire31 (.A(mclk_raw),
    .X(net1763));
 sky130_fd_sc_hd__buf_2 wire32 (.A(clknet_0_mclk_raw),
    .X(net1764));
 sky130_fd_sc_hd__buf_2 wire33 (.A(clknet_0_mclk_raw),
    .X(net1765));
 sky130_fd_sc_hd__clkbuf_4 wire34 (.A(net1767),
    .X(net1766));
 sky130_fd_sc_hd__clkbuf_4 wire35 (.A(clknet_2_0__leaf_mclk_raw),
    .X(net1767));
 sky130_fd_sc_hd__buf_6 wire36 (.A(net1769),
    .X(net1768));
 sky130_fd_sc_hd__clkbuf_4 wire38 (.A(clknet_2_2__leaf_mclk_raw),
    .X(net1770));
 sky130_fd_sc_hd__buf_2 wire39 (.A(clknet_2_2__leaf_mclk_raw),
    .X(net1771));
 sky130_fd_sc_hd__buf_2 wire4 (.A(\clknet_0_u_dsync.out_clk ),
    .X(net1736));
 sky130_fd_sc_hd__clkbuf_2 wire40 (.A(net1773),
    .X(net1772));
 sky130_fd_sc_hd__clkbuf_4 wire41 (.A(clknet_2_3__leaf_mclk_raw),
    .X(net1773));
 sky130_fd_sc_hd__clkbuf_4 wire477 (.A(_3577_),
    .X(net477));
 sky130_fd_sc_hd__buf_4 wire478 (.A(_3565_),
    .X(net478));
 sky130_fd_sc_hd__buf_4 wire479 (.A(_3557_),
    .X(net479));
 sky130_fd_sc_hd__buf_4 wire480 (.A(_3553_),
    .X(net480));
 sky130_fd_sc_hd__buf_4 wire485 (.A(_3478_),
    .X(net485));
 sky130_fd_sc_hd__buf_2 wire5 (.A(\clknet_0_u_dsync.out_clk ),
    .X(net1737));
 sky130_fd_sc_hd__buf_6 wire510 (.A(_2783_),
    .X(net510));
 sky130_fd_sc_hd__buf_6 wire511 (.A(_2782_),
    .X(net511));
 sky130_fd_sc_hd__buf_6 wire512 (.A(_2781_),
    .X(net512));
 sky130_fd_sc_hd__buf_6 wire515 (.A(_3586_),
    .X(net515));
 sky130_fd_sc_hd__buf_6 wire516 (.A(_3585_),
    .X(net516));
 sky130_fd_sc_hd__buf_4 wire517 (.A(_3584_),
    .X(net517));
 sky130_fd_sc_hd__buf_4 wire519 (.A(net518),
    .X(net519));
 sky130_fd_sc_hd__buf_4 wire549 (.A(_2780_),
    .X(net549));
 sky130_fd_sc_hd__buf_6 wire550 (.A(_2778_),
    .X(net550));
 sky130_fd_sc_hd__buf_6 wire551 (.A(_2777_),
    .X(net551));
 sky130_fd_sc_hd__buf_6 wire552 (.A(_2773_),
    .X(net552));
 sky130_fd_sc_hd__buf_6 wire553 (.A(_2752_),
    .X(net553));
 sky130_fd_sc_hd__buf_6 wire555 (.A(_2745_),
    .X(net555));
 sky130_fd_sc_hd__clkbuf_8 wire556 (.A(_2743_),
    .X(net556));
 sky130_fd_sc_hd__buf_6 wire557 (.A(_2742_),
    .X(net557));
 sky130_fd_sc_hd__buf_6 wire558 (.A(_2741_),
    .X(net558));
 sky130_fd_sc_hd__clkbuf_8 wire559 (.A(_2740_),
    .X(net559));
 sky130_fd_sc_hd__buf_6 wire560 (.A(_2736_),
    .X(net560));
 sky130_fd_sc_hd__buf_6 wire561 (.A(_2669_),
    .X(net561));
 sky130_fd_sc_hd__buf_6 wire572 (.A(net573),
    .X(net572));
 sky130_fd_sc_hd__buf_4 wire573 (.A(\u_dcg_s0.clk_enb ),
    .X(net573));
 sky130_fd_sc_hd__buf_6 wire575 (.A(net574),
    .X(net575));
 sky130_fd_sc_hd__buf_6 wire579 (.A(net578),
    .X(net579));
 sky130_fd_sc_hd__buf_8 wire585 (.A(net1885),
    .X(net585));
 sky130_fd_sc_hd__buf_6 wire590 (.A(net589),
    .X(net590));
 sky130_fd_sc_hd__buf_6 wire591 (.A(_2775_),
    .X(net591));
 sky130_fd_sc_hd__buf_8 wire592 (.A(_2751_),
    .X(net592));
 sky130_fd_sc_hd__buf_4 wire597 (.A(_2748_),
    .X(net597));
 sky130_fd_sc_hd__buf_4 wire6 (.A(\clknet_1_0_0_u_dsync.out_clk ),
    .X(net1738));
 sky130_fd_sc_hd__buf_6 wire602 (.A(_2744_),
    .X(net602));
 sky130_fd_sc_hd__buf_4 wire607 (.A(net606),
    .X(net607));
 sky130_fd_sc_hd__buf_6 wire609 (.A(_2717_),
    .X(net609));
 sky130_fd_sc_hd__buf_6 wire613 (.A(net612),
    .X(net613));
 sky130_fd_sc_hd__buf_4 wire615 (.A(net616),
    .X(net615));
 sky130_fd_sc_hd__clkbuf_8 wire616 (.A(net614),
    .X(net616));
 sky130_fd_sc_hd__buf_4 wire617 (.A(_2668_),
    .X(net617));
 sky130_fd_sc_hd__buf_4 wire625 (.A(_2663_),
    .X(net625));
 sky130_fd_sc_hd__buf_6 wire628 (.A(_2024_),
    .X(net628));
 sky130_fd_sc_hd__buf_6 wire629 (.A(_1963_),
    .X(net629));
 sky130_fd_sc_hd__buf_8 wire630 (.A(_1882_),
    .X(net630));
 sky130_fd_sc_hd__buf_6 wire631 (.A(_3248_),
    .X(net631));
 sky130_fd_sc_hd__buf_6 wire632 (.A(_3245_),
    .X(net632));
 sky130_fd_sc_hd__buf_6 wire633 (.A(net634),
    .X(net633));
 sky130_fd_sc_hd__buf_4 wire634 (.A(net2026),
    .X(net634));
 sky130_fd_sc_hd__buf_6 wire635 (.A(_3239_),
    .X(net635));
 sky130_fd_sc_hd__buf_6 wire636 (.A(net1833),
    .X(net636));
 sky130_fd_sc_hd__buf_6 wire637 (.A(net1888),
    .X(net637));
 sky130_fd_sc_hd__buf_6 wire638 (.A(net1919),
    .X(net638));
 sky130_fd_sc_hd__buf_6 wire639 (.A(net1933),
    .X(net639));
 sky130_fd_sc_hd__buf_4 wire640 (.A(_3221_),
    .X(net640));
 sky130_fd_sc_hd__buf_6 wire641 (.A(_3219_),
    .X(net641));
 sky130_fd_sc_hd__buf_6 wire642 (.A(net2014),
    .X(net642));
 sky130_fd_sc_hd__buf_6 wire643 (.A(_3212_),
    .X(net643));
 sky130_fd_sc_hd__buf_6 wire644 (.A(_3209_),
    .X(net644));
 sky130_fd_sc_hd__buf_6 wire645 (.A(net646),
    .X(net645));
 sky130_fd_sc_hd__buf_4 wire646 (.A(net1935),
    .X(net646));
 sky130_fd_sc_hd__buf_6 wire647 (.A(net1840),
    .X(net647));
 sky130_fd_sc_hd__buf_4 wire648 (.A(_3202_),
    .X(net648));
 sky130_fd_sc_hd__buf_6 wire649 (.A(_3200_),
    .X(net649));
 sky130_fd_sc_hd__buf_4 wire650 (.A(_3197_),
    .X(net650));
 sky130_fd_sc_hd__buf_6 wire651 (.A(_3193_),
    .X(net651));
 sky130_fd_sc_hd__buf_6 wire652 (.A(net653),
    .X(net652));
 sky130_fd_sc_hd__buf_4 wire653 (.A(_3191_),
    .X(net653));
 sky130_fd_sc_hd__buf_6 wire654 (.A(net2020),
    .X(net654));
 sky130_fd_sc_hd__buf_6 wire655 (.A(_3185_),
    .X(net655));
 sky130_fd_sc_hd__buf_6 wire656 (.A(_3182_),
    .X(net656));
 sky130_fd_sc_hd__buf_6 wire657 (.A(net2073),
    .X(net657));
 sky130_fd_sc_hd__buf_4 wire658 (.A(_3176_),
    .X(net658));
 sky130_fd_sc_hd__buf_4 wire659 (.A(_3174_),
    .X(net659));
 sky130_fd_sc_hd__buf_4 wire660 (.A(_3172_),
    .X(net660));
 sky130_fd_sc_hd__buf_6 wire661 (.A(net2069),
    .X(net661));
 sky130_fd_sc_hd__buf_4 wire662 (.A(_3167_),
    .X(net662));
 sky130_fd_sc_hd__buf_6 wire663 (.A(net1968),
    .X(net663));
 sky130_fd_sc_hd__buf_4 wire664 (.A(_3160_),
    .X(net664));
 sky130_fd_sc_hd__buf_4 wire665 (.A(_3157_),
    .X(net665));
 sky130_fd_sc_hd__buf_6 wire666 (.A(_3155_),
    .X(net666));
 sky130_fd_sc_hd__buf_6 wire667 (.A(net668),
    .X(net667));
 sky130_fd_sc_hd__buf_4 wire668 (.A(_3153_),
    .X(net668));
 sky130_fd_sc_hd__buf_6 wire669 (.A(net2053),
    .X(net669));
 sky130_fd_sc_hd__buf_6 wire670 (.A(_3147_),
    .X(net670));
 sky130_fd_sc_hd__buf_6 wire671 (.A(_3145_),
    .X(net671));
 sky130_fd_sc_hd__buf_6 wire672 (.A(_3143_),
    .X(net672));
 sky130_fd_sc_hd__buf_6 wire673 (.A(net674),
    .X(net673));
 sky130_fd_sc_hd__buf_4 wire674 (.A(_3140_),
    .X(net674));
 sky130_fd_sc_hd__buf_8 wire675 (.A(net676),
    .X(net675));
 sky130_fd_sc_hd__buf_6 wire676 (.A(net1916),
    .X(net676));
 sky130_fd_sc_hd__buf_8 wire677 (.A(net678),
    .X(net677));
 sky130_fd_sc_hd__buf_6 wire678 (.A(net2083),
    .X(net678));
 sky130_fd_sc_hd__buf_6 wire679 (.A(_2879_),
    .X(net679));
 sky130_fd_sc_hd__buf_4 wire680 (.A(_2871_),
    .X(net680));
 sky130_fd_sc_hd__buf_4 wire681 (.A(_2820_),
    .X(net681));
 sky130_fd_sc_hd__buf_4 wire682 (.A(_2814_),
    .X(net682));
 sky130_fd_sc_hd__buf_6 wire683 (.A(_2812_),
    .X(net683));
 sky130_fd_sc_hd__buf_4 wire684 (.A(_2809_),
    .X(net684));
 sky130_fd_sc_hd__buf_4 wire685 (.A(_2806_),
    .X(net685));
 sky130_fd_sc_hd__buf_4 wire686 (.A(_2803_),
    .X(net686));
 sky130_fd_sc_hd__buf_4 wire687 (.A(_2772_),
    .X(net687));
 sky130_fd_sc_hd__buf_8 wire688 (.A(net1986),
    .X(net688));
 sky130_fd_sc_hd__buf_6 wire689 (.A(net2024),
    .X(net689));
 sky130_fd_sc_hd__buf_8 wire690 (.A(net1896),
    .X(net690));
 sky130_fd_sc_hd__buf_8 wire691 (.A(net2011),
    .X(net691));
 sky130_fd_sc_hd__buf_6 wire692 (.A(_2759_),
    .X(net692));
 sky130_fd_sc_hd__buf_12 wire693 (.A(net694),
    .X(net693));
 sky130_fd_sc_hd__buf_6 wire694 (.A(_2757_),
    .X(net694));
 sky130_fd_sc_hd__buf_8 wire695 (.A(net696),
    .X(net695));
 sky130_fd_sc_hd__buf_6 wire696 (.A(_2755_),
    .X(net696));
 sky130_fd_sc_hd__buf_4 wire697 (.A(net698),
    .X(net697));
 sky130_fd_sc_hd__buf_4 wire698 (.A(_2735_),
    .X(net698));
 sky130_fd_sc_hd__buf_8 wire699 (.A(_2733_),
    .X(net699));
 sky130_fd_sc_hd__buf_6 wire700 (.A(_2731_),
    .X(net700));
 sky130_fd_sc_hd__buf_4 wire701 (.A(_2729_),
    .X(net701));
 sky130_fd_sc_hd__buf_6 wire702 (.A(net1948),
    .X(net702));
 sky130_fd_sc_hd__buf_4 wire703 (.A(_2723_),
    .X(net703));
 sky130_fd_sc_hd__buf_6 wire705 (.A(_2686_),
    .X(net705));
 sky130_fd_sc_hd__buf_6 wire706 (.A(_2684_),
    .X(net706));
 sky130_fd_sc_hd__buf_6 wire707 (.A(_2675_),
    .X(net707));
 sky130_fd_sc_hd__buf_6 wire708 (.A(_2672_),
    .X(net708));
 sky130_fd_sc_hd__buf_4 wire709 (.A(net348),
    .X(net709));
 sky130_fd_sc_hd__buf_4 wire710 (.A(net345),
    .X(net710));
 sky130_fd_sc_hd__buf_4 wire711 (.A(_2023_),
    .X(net711));
 sky130_fd_sc_hd__buf_4 wire712 (.A(net380),
    .X(net712));
 sky130_fd_sc_hd__buf_6 wire719 (.A(_1970_),
    .X(net719));
 sky130_fd_sc_hd__buf_6 wire720 (.A(_1967_),
    .X(net720));
 sky130_fd_sc_hd__buf_8 wire725 (.A(_1953_),
    .X(net725));
 sky130_fd_sc_hd__buf_12 wire726 (.A(_1944_),
    .X(net726));
 sky130_fd_sc_hd__buf_4 wire727 (.A(net334),
    .X(net727));
 sky130_fd_sc_hd__clkbuf_4 wire728 (.A(net336),
    .X(net728));
 sky130_fd_sc_hd__clkbuf_4 wire729 (.A(net337),
    .X(net729));
 sky130_fd_sc_hd__buf_4 wire730 (.A(net338),
    .X(net730));
 sky130_fd_sc_hd__buf_4 wire731 (.A(net339),
    .X(net731));
 sky130_fd_sc_hd__buf_6 wire732 (.A(_1837_),
    .X(net732));
 sky130_fd_sc_hd__buf_6 wire737 (.A(net738),
    .X(net737));
 sky130_fd_sc_hd__buf_4 wire738 (.A(_1719_),
    .X(net738));
 sky130_fd_sc_hd__buf_8 wire783 (.A(_1939_),
    .X(net783));
 sky130_fd_sc_hd__buf_6 wire784 (.A(_1938_),
    .X(net784));
 sky130_fd_sc_hd__buf_8 wire785 (.A(_1934_),
    .X(net785));
 sky130_fd_sc_hd__buf_4 wire786 (.A(_1932_),
    .X(net786));
 sky130_fd_sc_hd__buf_6 wire787 (.A(_1931_),
    .X(net787));
 sky130_fd_sc_hd__buf_8 wire788 (.A(_1929_),
    .X(net788));
 sky130_fd_sc_hd__buf_6 wire789 (.A(_1927_),
    .X(net789));
 sky130_fd_sc_hd__buf_6 wire790 (.A(_1926_),
    .X(net790));
 sky130_fd_sc_hd__buf_8 wire791 (.A(_1924_),
    .X(net791));
 sky130_fd_sc_hd__buf_4 wire792 (.A(net793),
    .X(net792));
 sky130_fd_sc_hd__buf_4 wire793 (.A(_1922_),
    .X(net793));
 sky130_fd_sc_hd__buf_8 wire794 (.A(_1921_),
    .X(net794));
 sky130_fd_sc_hd__buf_4 wire795 (.A(net796),
    .X(net795));
 sky130_fd_sc_hd__buf_4 wire796 (.A(_1918_),
    .X(net796));
 sky130_fd_sc_hd__buf_4 wire797 (.A(_1863_),
    .X(net797));
 sky130_fd_sc_hd__buf_4 wire798 (.A(_1858_),
    .X(net798));
 sky130_fd_sc_hd__buf_4 wire8 (.A(net1741),
    .X(net1740));
 sky130_fd_sc_hd__buf_4 wire807 (.A(_1847_),
    .X(net807));
 sky130_fd_sc_hd__buf_6 wire867 (.A(net866),
    .X(net867));
 sky130_fd_sc_hd__buf_4 wire920 (.A(\u_dcg_peri.reset_n ),
    .X(net920));
 assign m0_wbd_err_o = net1721;
 assign m1_wbd_err_o = net1722;
 assign m2_wbd_err_o = net1723;
 assign m3_wbd_err_o = net1724;
 assign s0_wbd_adr_o[0] = net1725;
 assign s0_wbd_adr_o[1] = net1726;
 assign s1_wbd_adr_o[0] = net1727;
 assign s1_wbd_adr_o[1] = net1728;
 assign s2_wbd_adr_o[0] = net1729;
 assign s2_wbd_adr_o[1] = net1730;
endmodule

