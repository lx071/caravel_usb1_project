magic
tech sky130A
magscale 1 2
timestamp 1698804265
<< viali >>
rect 213653 5185 213687 5219
rect 116225 4981 116259 5015
rect 116869 4981 116903 5015
rect 117513 4981 117547 5015
rect 118249 4981 118283 5015
rect 210985 4981 211019 5015
rect 211629 4981 211663 5015
rect 214297 4981 214331 5015
rect 214849 4981 214883 5015
rect 215401 4981 215435 5015
rect 216229 4981 216263 5015
rect 216781 4981 216815 5015
rect 306205 4981 306239 5015
rect 306757 4981 306791 5015
rect 307585 4981 307619 5015
rect 308045 4981 308079 5015
rect 308689 4981 308723 5015
rect 308505 4777 308539 4811
rect 308321 4573 308355 4607
rect 215769 4505 215803 4539
rect 115489 4437 115523 4471
rect 116041 4437 116075 4471
rect 116593 4437 116627 4471
rect 117881 4437 117915 4471
rect 118433 4437 118467 4471
rect 118985 4437 119019 4471
rect 119537 4437 119571 4471
rect 120733 4437 120767 4471
rect 121377 4437 121411 4471
rect 122481 4437 122515 4471
rect 210433 4437 210467 4471
rect 211077 4437 211111 4471
rect 211629 4437 211663 4471
rect 212365 4437 212399 4471
rect 213009 4437 213043 4471
rect 213561 4437 213595 4471
rect 214021 4437 214055 4471
rect 214665 4437 214699 4471
rect 216781 4437 216815 4471
rect 217241 4437 217275 4471
rect 217885 4437 217919 4471
rect 305653 4437 305687 4471
rect 306205 4437 306239 4471
rect 306757 4437 306791 4471
rect 307401 4437 307435 4471
rect 309149 4437 309183 4471
rect 309609 4437 309643 4471
rect 310437 4437 310471 4471
rect 211813 4165 211847 4199
rect 115765 4097 115799 4131
rect 116869 4097 116903 4131
rect 118709 4097 118743 4131
rect 120733 4097 120767 4131
rect 121929 4097 121963 4131
rect 124505 4097 124539 4131
rect 125149 4097 125183 4131
rect 209053 4097 209087 4131
rect 210157 4097 210191 4131
rect 211261 4097 211295 4131
rect 212825 4097 212859 4131
rect 213377 4097 213411 4131
rect 213929 4097 213963 4131
rect 215493 4097 215527 4131
rect 217011 4097 217045 4131
rect 306481 4097 306515 4131
rect 307493 4097 307527 4131
rect 309149 4097 309183 4131
rect 310529 4097 310563 4131
rect 115213 4029 115247 4063
rect 117421 4029 117455 4063
rect 118157 4029 118191 4063
rect 121653 4029 121687 4063
rect 122573 4029 122607 4063
rect 123493 4029 123527 4063
rect 209605 4029 209639 4063
rect 214941 4029 214975 4063
rect 216689 4029 216723 4063
rect 304181 4029 304215 4063
rect 304825 4029 304859 4063
rect 306205 4029 306239 4063
rect 308873 4029 308907 4063
rect 310713 3961 310747 3995
rect 119353 3893 119387 3927
rect 120273 3893 120307 3927
rect 208409 3893 208443 3927
rect 217793 3893 217827 3927
rect 218529 3893 218563 3927
rect 219541 3893 219575 3927
rect 305469 3893 305503 3927
rect 307033 3893 307067 3927
rect 307677 3893 307711 3927
rect 309701 3893 309735 3927
rect 311357 3893 311391 3927
rect 113833 3689 113867 3723
rect 125885 3689 125919 3723
rect 126437 3689 126471 3723
rect 220461 3689 220495 3723
rect 313197 3689 313231 3723
rect 211629 3553 211663 3587
rect 216505 3553 216539 3587
rect 309057 3553 309091 3587
rect 309977 3553 310011 3587
rect 114385 3485 114419 3519
rect 115489 3485 115523 3519
rect 116685 3485 116719 3519
rect 118157 3485 118191 3519
rect 118801 3485 118835 3519
rect 119353 3485 119387 3519
rect 120089 3485 120123 3519
rect 120549 3485 120583 3519
rect 121285 3485 121319 3519
rect 124321 3485 124355 3519
rect 125333 3485 125367 3519
rect 208317 3485 208351 3519
rect 208869 3485 208903 3519
rect 209421 3485 209455 3519
rect 210985 3485 211019 3519
rect 212181 3485 212215 3519
rect 213377 3485 213411 3519
rect 214573 3485 214607 3519
rect 215309 3485 215343 3519
rect 217057 3485 217091 3519
rect 217701 3485 217735 3519
rect 218253 3485 218287 3519
rect 218897 3485 218931 3519
rect 219449 3485 219483 3519
rect 303445 3485 303479 3519
rect 303997 3485 304031 3519
rect 304549 3485 304583 3519
rect 305285 3485 305319 3519
rect 305561 3485 305595 3519
rect 306205 3485 306239 3519
rect 306481 3485 306515 3519
rect 307401 3485 307435 3519
rect 308137 3485 308171 3519
rect 308413 3485 308447 3519
rect 309333 3485 309367 3519
rect 310253 3485 310287 3519
rect 310897 3485 310931 3519
rect 311173 3485 311207 3519
rect 114937 3417 114971 3451
rect 116133 3417 116167 3451
rect 117605 3417 117639 3451
rect 121837 3417 121871 3451
rect 123769 3417 123803 3451
rect 125057 3417 125091 3451
rect 210433 3417 210467 3451
rect 212825 3417 212859 3451
rect 214021 3417 214055 3451
rect 215861 3417 215895 3451
rect 300869 3417 300903 3451
rect 307125 3417 307159 3451
rect 311725 3417 311759 3451
rect 122573 3349 122607 3383
rect 123217 3349 123251 3383
rect 300133 3349 300167 3383
rect 302801 3349 302835 3383
rect 312277 3349 312311 3383
rect 357173 3349 357207 3383
rect 393605 3349 393639 3383
rect 394249 3349 394283 3383
rect 394709 3349 394743 3383
rect 396733 3349 396767 3383
rect 221105 3145 221139 3179
rect 309149 3145 309183 3179
rect 314761 3145 314795 3179
rect 317889 3145 317923 3179
rect 331321 3145 331355 3179
rect 340061 3145 340095 3179
rect 344293 3145 344327 3179
rect 345029 3145 345063 3179
rect 353309 3145 353343 3179
rect 353953 3145 353987 3179
rect 357541 3145 357575 3179
rect 115121 3077 115155 3111
rect 116317 3077 116351 3111
rect 118709 3077 118743 3111
rect 120273 3077 120307 3111
rect 123861 3077 123895 3111
rect 127265 3077 127299 3111
rect 213009 3077 213043 3111
rect 214205 3077 214239 3111
rect 216597 3077 216631 3111
rect 219909 3077 219943 3111
rect 307401 3077 307435 3111
rect 309425 3077 309459 3111
rect 310713 3077 310747 3111
rect 344385 3077 344419 3111
rect 362233 3077 362267 3111
rect 416329 3077 416363 3111
rect 114109 3009 114143 3043
rect 115673 3009 115707 3043
rect 116869 3009 116903 3043
rect 118065 3009 118099 3043
rect 119261 3009 119295 3043
rect 120825 3009 120859 3043
rect 122021 3009 122055 3043
rect 123217 3009 123251 3043
rect 124413 3009 124447 3043
rect 125425 3009 125459 3043
rect 125701 3009 125735 3043
rect 126253 3009 126287 3043
rect 145849 3009 145883 3043
rect 164341 3009 164375 3043
rect 168665 3009 168699 3043
rect 202429 3009 202463 3043
rect 202797 3009 202831 3043
rect 205465 3009 205499 3043
rect 207581 3009 207615 3043
rect 209605 3009 209639 3043
rect 210801 3009 210835 3043
rect 211997 3009 212031 3043
rect 213561 3009 213595 3043
rect 214757 3009 214791 3043
rect 215953 3009 215987 3043
rect 217149 3009 217183 3043
rect 218713 3009 218747 3043
rect 219265 3009 219299 3043
rect 220461 3009 220495 3043
rect 254041 3009 254075 3043
rect 259101 3009 259135 3043
rect 259653 3009 259687 3043
rect 296545 3009 296579 3043
rect 297373 3009 297407 3043
rect 298017 3009 298051 3043
rect 298661 3009 298695 3043
rect 300225 3009 300259 3043
rect 300593 3009 300627 3043
rect 301145 3009 301179 3043
rect 303169 3009 303203 3043
rect 304365 3009 304399 3043
rect 305837 3009 305871 3043
rect 306665 3009 306699 3043
rect 307677 3009 307711 3043
rect 308597 3009 308631 3043
rect 310989 3009 311023 3043
rect 311909 3009 311943 3043
rect 312737 3009 312771 3043
rect 314025 3009 314059 3043
rect 314577 3009 314611 3043
rect 317337 3009 317371 3043
rect 331413 3009 331447 3043
rect 340153 3009 340187 3043
rect 340797 3009 340831 3043
rect 353769 3009 353803 3043
rect 357357 3009 357391 3043
rect 390201 3009 390235 3043
rect 390569 3009 390603 3043
rect 392961 3009 392995 3043
rect 393329 3009 393363 3043
rect 394433 3009 394467 3043
rect 396733 3009 396767 3043
rect 397101 3009 397135 3043
rect 398113 3009 398147 3043
rect 452853 3009 452887 3043
rect 453405 3009 453439 3043
rect 113557 2941 113591 2975
rect 117513 2941 117547 2975
rect 121561 2941 121595 2975
rect 122941 2941 122975 2975
rect 169217 2941 169251 2975
rect 204913 2941 204947 2975
rect 208133 2941 208167 2975
rect 209053 2941 209087 2975
rect 210249 2941 210283 2975
rect 211445 2941 211479 2975
rect 215401 2941 215435 2975
rect 302893 2941 302927 2975
rect 303813 2941 303847 2975
rect 305561 2941 305595 2975
rect 308321 2941 308355 2975
rect 311633 2941 311667 2975
rect 312461 2941 312495 2975
rect 315773 2941 315807 2975
rect 391673 2941 391707 2975
rect 394985 2941 395019 2975
rect 452577 2941 452611 2975
rect 126713 2873 126747 2907
rect 297557 2873 297591 2907
rect 301329 2873 301363 2907
rect 306481 2873 306515 2907
rect 317153 2873 317187 2907
rect 332057 2873 332091 2907
rect 470425 2873 470459 2907
rect 37657 2805 37691 2839
rect 74549 2805 74583 2839
rect 75009 2805 75043 2839
rect 108221 2805 108255 2839
rect 112177 2805 112211 2839
rect 113005 2805 113039 2839
rect 143181 2805 143215 2839
rect 152289 2805 152323 2839
rect 164801 2805 164835 2839
rect 168021 2805 168055 2839
rect 201693 2805 201727 2839
rect 206109 2805 206143 2839
rect 206845 2805 206879 2839
rect 218161 2805 218195 2839
rect 221657 2805 221691 2839
rect 247233 2805 247267 2839
rect 251557 2805 251591 2839
rect 260297 2805 260331 2839
rect 295993 2805 296027 2839
rect 299581 2805 299615 2839
rect 301789 2805 301823 2839
rect 313381 2805 313415 2839
rect 319085 2805 319119 2839
rect 319637 2805 319671 2839
rect 323777 2805 323811 2839
rect 324789 2805 324823 2839
rect 325341 2805 325375 2839
rect 332609 2805 332643 2839
rect 337485 2805 337519 2839
rect 338129 2805 338163 2839
rect 341533 2805 341567 2839
rect 342085 2805 342119 2839
rect 345581 2805 345615 2839
rect 346685 2805 346719 2839
rect 348617 2805 348651 2839
rect 349905 2805 349939 2839
rect 350549 2805 350583 2839
rect 352573 2805 352607 2839
rect 354505 2805 354539 2839
rect 356161 2805 356195 2839
rect 358185 2805 358219 2839
rect 380909 2805 380943 2839
rect 391213 2805 391247 2839
rect 396181 2805 396215 2839
rect 398941 2805 398975 2839
rect 400045 2805 400079 2839
rect 400965 2805 400999 2839
rect 408509 2805 408543 2839
rect 435005 2805 435039 2839
rect 435833 2805 435867 2839
rect 1869 2601 1903 2635
rect 19901 2601 19935 2635
rect 55965 2601 55999 2635
rect 58173 2601 58207 2635
rect 70409 2601 70443 2635
rect 73997 2601 74031 2635
rect 182189 2601 182223 2635
rect 301513 2601 301547 2635
rect 302893 2601 302927 2635
rect 304733 2601 304767 2635
rect 308413 2601 308447 2635
rect 314393 2601 314427 2635
rect 318349 2601 318383 2635
rect 319637 2601 319671 2635
rect 348341 2601 348375 2635
rect 350457 2601 350491 2635
rect 355149 2601 355183 2635
rect 355885 2601 355919 2635
rect 359565 2601 359599 2635
rect 362509 2601 362543 2635
rect 380541 2601 380575 2635
rect 382749 2601 382783 2635
rect 387165 2601 387199 2635
rect 395629 2601 395663 2635
rect 398573 2601 398607 2635
rect 56701 2533 56735 2567
rect 148241 2533 148275 2567
rect 242909 2533 242943 2567
rect 325341 2533 325375 2567
rect 341441 2533 341475 2567
rect 422585 2533 422619 2567
rect 434637 2533 434671 2567
rect 71605 2465 71639 2499
rect 110797 2465 110831 2499
rect 113557 2465 113591 2499
rect 114937 2465 114971 2499
rect 116777 2465 116811 2499
rect 149345 2465 149379 2499
rect 211813 2465 211847 2499
rect 219173 2465 219207 2499
rect 291117 2465 291151 2499
rect 293785 2465 293819 2499
rect 297741 2465 297775 2499
rect 367293 2465 367327 2499
rect 368489 2465 368523 2499
rect 385325 2465 385359 2499
rect 404001 2465 404035 2499
rect 407221 2465 407255 2499
rect 411821 2465 411855 2499
rect 461041 2465 461075 2499
rect 2053 2397 2087 2431
rect 20085 2397 20119 2431
rect 20637 2397 20671 2431
rect 36450 2397 36484 2431
rect 38117 2397 38151 2431
rect 42625 2397 42659 2431
rect 48881 2397 48915 2431
rect 53849 2397 53883 2431
rect 54401 2397 54435 2431
rect 54677 2397 54711 2431
rect 56149 2397 56183 2431
rect 58725 2397 58759 2431
rect 63233 2397 63267 2431
rect 63509 2397 63543 2431
rect 66821 2397 66855 2431
rect 71053 2397 71087 2431
rect 74181 2397 74215 2431
rect 74733 2397 74767 2431
rect 92029 2397 92063 2431
rect 92673 2397 92707 2431
rect 98101 2397 98135 2431
rect 98653 2397 98687 2431
rect 103897 2397 103931 2431
rect 104541 2397 104575 2431
rect 107393 2397 107427 2431
rect 107669 2397 107703 2431
rect 108405 2397 108439 2431
rect 110245 2397 110279 2431
rect 112361 2397 112395 2431
rect 114109 2397 114143 2431
rect 116133 2397 116167 2431
rect 118065 2397 118099 2431
rect 119261 2397 119295 2431
rect 120641 2397 120675 2431
rect 121837 2397 121871 2431
rect 123217 2397 123251 2431
rect 124413 2397 124447 2431
rect 125517 2397 125551 2431
rect 126069 2397 126103 2431
rect 126621 2397 126655 2431
rect 128277 2397 128311 2431
rect 130853 2397 130887 2431
rect 131405 2397 131439 2431
rect 136741 2397 136775 2431
rect 137293 2397 137327 2431
rect 143365 2397 143399 2431
rect 143917 2397 143951 2431
rect 146309 2397 146343 2431
rect 148885 2397 148919 2431
rect 152197 2397 152231 2431
rect 153485 2397 153519 2431
rect 156705 2397 156739 2431
rect 157349 2397 157383 2431
rect 161305 2397 161339 2431
rect 164341 2397 164375 2431
rect 165077 2397 165111 2431
rect 170229 2397 170263 2431
rect 182373 2397 182407 2431
rect 192217 2397 192251 2431
rect 193045 2397 193079 2431
rect 198565 2397 198599 2431
rect 200221 2397 200255 2431
rect 200865 2397 200899 2431
rect 203349 2397 203383 2431
rect 203901 2397 203935 2431
rect 205557 2397 205591 2431
rect 207673 2397 207707 2431
rect 208225 2397 208259 2431
rect 209421 2397 209455 2431
rect 211077 2397 211111 2431
rect 211537 2397 211571 2431
rect 213377 2397 213411 2431
rect 214573 2397 214607 2431
rect 215953 2397 215987 2431
rect 217149 2397 217183 2431
rect 218437 2397 218471 2431
rect 219725 2397 219759 2431
rect 220461 2397 220495 2431
rect 221013 2397 221047 2431
rect 223589 2397 223623 2431
rect 224969 2397 225003 2431
rect 225613 2397 225647 2431
rect 230765 2397 230799 2431
rect 231409 2397 231443 2431
rect 236469 2397 236503 2431
rect 237757 2397 237791 2431
rect 238493 2397 238527 2431
rect 239045 2397 239079 2431
rect 243645 2397 243679 2431
rect 247141 2397 247175 2431
rect 248797 2397 248831 2431
rect 249349 2397 249383 2431
rect 251741 2397 251775 2431
rect 254501 2397 254535 2431
rect 256525 2397 256559 2431
rect 259469 2397 259503 2431
rect 260021 2397 260055 2431
rect 262321 2397 262355 2431
rect 262965 2397 262999 2431
rect 263517 2397 263551 2431
rect 265173 2397 265207 2431
rect 272533 2397 272567 2431
rect 273085 2397 273119 2431
rect 277685 2397 277719 2431
rect 286517 2397 286551 2431
rect 287437 2397 287471 2431
rect 290565 2397 290599 2431
rect 293233 2397 293267 2431
rect 295441 2397 295475 2431
rect 296453 2397 296487 2431
rect 297005 2397 297039 2431
rect 298017 2397 298051 2431
rect 299581 2397 299615 2431
rect 300317 2397 300351 2431
rect 301789 2397 301823 2431
rect 303445 2397 303479 2431
rect 304549 2397 304583 2431
rect 306021 2397 306055 2431
rect 306757 2397 306791 2431
rect 309517 2397 309551 2431
rect 310713 2397 310747 2431
rect 310989 2397 311023 2431
rect 312369 2397 312403 2431
rect 313749 2397 313783 2431
rect 315681 2397 315715 2431
rect 317613 2397 317647 2431
rect 318993 2397 319027 2431
rect 319453 2397 319487 2431
rect 323593 2397 323627 2431
rect 324697 2397 324731 2431
rect 325157 2397 325191 2431
rect 326629 2397 326663 2431
rect 327181 2397 327215 2431
rect 329389 2397 329423 2431
rect 330033 2397 330067 2431
rect 331781 2397 331815 2431
rect 332333 2397 332367 2431
rect 333069 2397 333103 2431
rect 335461 2397 335495 2431
rect 336381 2397 336415 2431
rect 337853 2397 337887 2431
rect 340521 2397 340555 2431
rect 341625 2397 341659 2431
rect 342177 2397 342211 2431
rect 342913 2397 342947 2431
rect 344661 2397 344695 2431
rect 346593 2397 346627 2431
rect 347329 2397 347363 2431
rect 350273 2397 350307 2431
rect 353677 2397 353711 2431
rect 356069 2397 356103 2431
rect 357265 2397 357299 2431
rect 358461 2397 358495 2431
rect 362601 2397 362635 2431
rect 367845 2397 367879 2431
rect 371709 2397 371743 2431
rect 380725 2397 380759 2431
rect 381277 2397 381311 2431
rect 381829 2397 381863 2431
rect 385877 2397 385911 2431
rect 387901 2397 387935 2431
rect 388453 2397 388487 2431
rect 389557 2397 389591 2431
rect 391121 2397 391155 2431
rect 394433 2397 394467 2431
rect 396917 2397 396951 2431
rect 397377 2397 397411 2431
rect 398757 2397 398791 2431
rect 399861 2397 399895 2431
rect 401149 2397 401183 2431
rect 404645 2397 404679 2431
rect 407773 2397 407807 2431
rect 408417 2397 408451 2431
rect 409337 2397 409371 2431
rect 412373 2397 412407 2431
rect 416789 2397 416823 2431
rect 421389 2397 421423 2431
rect 421941 2397 421975 2431
rect 425713 2397 425747 2431
rect 434821 2397 434855 2431
rect 435741 2397 435775 2431
rect 439973 2397 440007 2431
rect 448069 2397 448103 2431
rect 452853 2397 452887 2431
rect 461317 2397 461351 2431
rect 465733 2397 465767 2431
rect 466009 2397 466043 2431
rect 470885 2397 470919 2431
rect 474657 2397 474691 2431
rect 479257 2397 479291 2431
rect 36737 2329 36771 2363
rect 42901 2329 42935 2363
rect 49157 2329 49191 2363
rect 59001 2329 59035 2363
rect 67097 2329 67131 2363
rect 75285 2329 75319 2363
rect 96905 2329 96939 2363
rect 105093 2329 105127 2363
rect 108957 2329 108991 2363
rect 112913 2329 112947 2363
rect 117513 2329 117547 2363
rect 118709 2329 118743 2363
rect 120181 2329 120215 2363
rect 121469 2329 121503 2363
rect 122849 2329 122883 2363
rect 123861 2329 123895 2363
rect 125241 2329 125275 2363
rect 151001 2329 151035 2363
rect 154037 2329 154071 2363
rect 157901 2329 157935 2363
rect 161857 2329 161891 2363
rect 165537 2329 165571 2363
rect 169033 2329 169067 2363
rect 199117 2329 199151 2363
rect 206109 2329 206143 2363
rect 206937 2329 206971 2363
rect 208869 2329 208903 2363
rect 210249 2329 210283 2363
rect 212825 2329 212859 2363
rect 214021 2329 214055 2363
rect 215401 2329 215435 2363
rect 216597 2329 216631 2363
rect 221565 2329 221599 2363
rect 223037 2329 223071 2363
rect 226165 2329 226199 2363
rect 231961 2329 231995 2363
rect 244197 2329 244231 2363
rect 246313 2329 246347 2363
rect 252293 2329 252327 2363
rect 257077 2329 257111 2363
rect 264345 2329 264379 2363
rect 277133 2329 277167 2363
rect 285965 2329 285999 2363
rect 295809 2329 295843 2363
rect 299029 2329 299063 2363
rect 300777 2329 300811 2363
rect 303997 2329 304031 2363
rect 305469 2329 305503 2363
rect 307309 2329 307343 2363
rect 308505 2329 308539 2363
rect 309241 2329 309275 2363
rect 311817 2329 311851 2363
rect 313289 2329 313323 2363
rect 314669 2329 314703 2363
rect 317061 2329 317095 2363
rect 331229 2329 331263 2363
rect 335277 2329 335311 2363
rect 337301 2329 337335 2363
rect 339969 2329 340003 2363
rect 345765 2329 345799 2363
rect 348433 2329 348467 2363
rect 349721 2329 349755 2363
rect 352389 2329 352423 2363
rect 353309 2329 353343 2363
rect 354505 2329 354539 2363
rect 357909 2329 357943 2363
rect 371157 2329 371191 2363
rect 372445 2329 372479 2363
rect 389281 2329 389315 2363
rect 391673 2329 391707 2363
rect 393881 2329 393915 2363
rect 395905 2329 395939 2363
rect 399309 2329 399343 2363
rect 401517 2329 401551 2363
rect 405197 2329 405231 2363
rect 408693 2329 408727 2363
rect 425161 2329 425195 2363
rect 435465 2329 435499 2363
rect 439421 2329 439455 2363
rect 447793 2329 447827 2363
rect 474381 2329 474415 2363
rect 478981 2329 479015 2363
rect 492413 2329 492447 2363
rect 2605 2261 2639 2295
rect 35909 2261 35943 2295
rect 37933 2261 37967 2295
rect 41981 2261 42015 2295
rect 48329 2261 48363 2295
rect 62589 2261 62623 2295
rect 66269 2261 66303 2295
rect 92213 2261 92247 2295
rect 110061 2261 110095 2295
rect 128093 2261 128127 2295
rect 128829 2261 128863 2295
rect 130209 2261 130243 2295
rect 136097 2261 136131 2295
rect 146125 2261 146159 2295
rect 152749 2261 152783 2295
rect 160477 2261 160511 2295
rect 164157 2261 164191 2295
rect 170781 2261 170815 2295
rect 182925 2261 182959 2295
rect 193597 2261 193631 2295
rect 197921 2261 197955 2295
rect 200405 2261 200439 2295
rect 202705 2261 202739 2295
rect 204913 2261 204947 2295
rect 218253 2261 218287 2295
rect 224233 2261 224267 2295
rect 236285 2261 236319 2295
rect 237021 2261 237055 2295
rect 248061 2261 248095 2295
rect 254317 2261 254351 2295
rect 255789 2261 255823 2295
rect 258365 2261 258399 2295
rect 265725 2261 265759 2295
rect 272349 2261 272383 2295
rect 278329 2261 278363 2295
rect 290381 2261 290415 2295
rect 292589 2261 292623 2295
rect 311541 2261 311575 2295
rect 318809 2261 318843 2295
rect 323409 2261 323443 2295
rect 324513 2261 324547 2295
rect 326445 2261 326479 2295
rect 329297 2261 329331 2295
rect 332517 2261 332551 2295
rect 337209 2261 337243 2295
rect 338037 2261 338071 2295
rect 342361 2261 342395 2295
rect 344477 2261 344511 2295
rect 345673 2261 345707 2295
rect 346777 2261 346811 2295
rect 349629 2261 349663 2295
rect 352297 2261 352331 2295
rect 354413 2261 354447 2295
rect 357081 2261 357115 2295
rect 386521 2261 386555 2295
rect 390477 2261 390511 2295
rect 413017 2261 413051 2295
rect 416605 2261 416639 2295
rect 426541 2261 426575 2295
rect 440617 2261 440651 2295
rect 448621 2261 448655 2295
rect 452669 2261 452703 2295
rect 453405 2261 453439 2295
rect 461869 2261 461903 2295
rect 466561 2261 466595 2295
rect 470701 2261 470735 2295
rect 475485 2261 475519 2295
rect 479809 2261 479843 2295
rect 492137 2261 492171 2295
rect 493517 2261 493551 2295
<< metal1 >>
rect 74 9228 130 10000
rect 1854 9228 1860 9240
rect 74 9200 1860 9228
rect 1854 9188 1860 9200
rect 1912 9188 1918 9240
rect 17074 9228 17130 10000
rect 17052 9200 17130 9228
rect 34074 9228 34130 10000
rect 34422 9228 34428 9240
rect 34074 9200 34428 9228
rect 17052 9160 17080 9200
rect 34422 9188 34428 9200
rect 34480 9188 34486 9240
rect 51074 9228 51130 10000
rect 52362 9228 52368 9240
rect 51074 9200 52368 9228
rect 52362 9188 52368 9200
rect 52420 9188 52426 9240
rect 68074 9228 68130 10000
rect 68922 9228 68928 9240
rect 68074 9200 68928 9228
rect 68922 9188 68928 9200
rect 68980 9188 68986 9240
rect 85074 9228 85130 10000
rect 85040 9200 85130 9228
rect 102074 9228 102130 10000
rect 102226 9228 102232 9240
rect 102074 9200 102232 9228
rect 85040 9160 85068 9200
rect 102226 9188 102232 9200
rect 102284 9188 102290 9240
rect 119074 9228 119130 10000
rect 119982 9228 119988 9240
rect 119074 9200 119988 9228
rect 119982 9188 119988 9200
rect 120040 9188 120046 9240
rect 136074 9228 136130 10000
rect 136542 9228 136548 9240
rect 136074 9200 136548 9228
rect 136542 9188 136548 9200
rect 136600 9188 136606 9240
rect 153074 9228 153130 10000
rect 170074 9228 170130 10000
rect 153074 9200 153148 9228
rect 153120 9160 153148 9200
rect 17052 9132 17126 9160
rect 85040 9132 85114 9160
rect 17098 8888 17126 9132
rect 17862 8888 17868 8900
rect 17098 8860 17868 8888
rect 17862 8848 17868 8860
rect 17920 8848 17926 8900
rect 85086 8888 85114 9132
rect 153074 9132 153148 9160
rect 170048 9200 170130 9228
rect 187074 9228 187130 10000
rect 187602 9228 187608 9240
rect 187074 9200 187608 9228
rect 170048 9160 170076 9200
rect 187602 9188 187608 9200
rect 187660 9188 187666 9240
rect 204074 9228 204130 10000
rect 204162 9228 204168 9240
rect 204074 9200 204168 9228
rect 204162 9188 204168 9200
rect 204220 9188 204226 9240
rect 221074 9228 221130 10000
rect 222102 9228 222108 9240
rect 221074 9200 222108 9228
rect 222102 9188 222108 9200
rect 222160 9188 222166 9240
rect 238074 9228 238130 10000
rect 255074 9228 255130 10000
rect 238074 9200 238156 9228
rect 238128 9160 238156 9200
rect 170048 9132 170122 9160
rect 153074 8968 153102 9132
rect 153074 8928 153108 8968
rect 153102 8916 153108 8928
rect 153160 8916 153166 8968
rect 170094 8956 170122 9132
rect 238082 9132 238156 9160
rect 255056 9200 255130 9228
rect 272074 9228 272130 10000
rect 273162 9228 273168 9240
rect 272074 9200 273168 9228
rect 255056 9160 255084 9200
rect 273162 9188 273168 9200
rect 273220 9188 273226 9240
rect 289074 9228 289130 10000
rect 289446 9228 289452 9240
rect 289074 9200 289452 9228
rect 289446 9188 289452 9200
rect 289504 9188 289510 9240
rect 306074 9228 306130 10000
rect 306024 9200 306130 9228
rect 323074 9228 323130 10000
rect 340074 9228 340130 10000
rect 340782 9228 340788 9240
rect 323074 9200 323164 9228
rect 340074 9200 340788 9228
rect 306024 9160 306052 9200
rect 323136 9160 323164 9200
rect 340782 9188 340788 9200
rect 340840 9188 340846 9240
rect 357074 9228 357130 10000
rect 357250 9228 357256 9240
rect 357074 9200 357256 9228
rect 357250 9188 357256 9200
rect 357308 9188 357314 9240
rect 374074 9228 374130 10000
rect 375282 9228 375288 9240
rect 374074 9200 375288 9228
rect 375282 9188 375288 9200
rect 375340 9188 375346 9240
rect 391074 9228 391130 10000
rect 408074 9228 408130 10000
rect 391032 9200 391130 9228
rect 408052 9200 408130 9228
rect 425074 9228 425130 10000
rect 426342 9228 426348 9240
rect 425074 9200 426348 9228
rect 255056 9132 255130 9160
rect 306024 9132 306116 9160
rect 171042 8956 171048 8968
rect 170094 8928 171048 8956
rect 171042 8916 171048 8928
rect 171100 8916 171106 8968
rect 238082 8956 238110 9132
rect 238662 8956 238668 8968
rect 238082 8928 238668 8956
rect 238662 8916 238668 8928
rect 238720 8916 238726 8968
rect 85482 8888 85488 8900
rect 85086 8860 85488 8888
rect 85482 8848 85488 8860
rect 85540 8848 85546 8900
rect 255102 8888 255130 9132
rect 306088 8956 306116 9132
rect 323090 9132 323164 9160
rect 391032 9160 391060 9200
rect 408052 9160 408080 9200
rect 426342 9188 426348 9200
rect 426400 9188 426406 9240
rect 442074 9228 442130 10000
rect 442902 9228 442908 9240
rect 442074 9200 442908 9228
rect 442902 9188 442908 9200
rect 442960 9188 442966 9240
rect 391032 9132 391106 9160
rect 408052 9132 408126 9160
rect 306282 8956 306288 8968
rect 306088 8928 306288 8956
rect 306282 8916 306288 8928
rect 306340 8916 306346 8968
rect 323090 8956 323118 9132
rect 324222 8956 324228 8968
rect 323090 8928 324228 8956
rect 324222 8916 324228 8928
rect 324280 8916 324286 8968
rect 391078 8956 391106 9132
rect 391842 8956 391848 8968
rect 391078 8928 391848 8956
rect 391842 8916 391848 8928
rect 391900 8916 391906 8968
rect 408098 8956 408126 9132
rect 408402 8956 408408 8968
rect 408098 8928 408408 8956
rect 408402 8916 408408 8928
rect 408460 8916 408466 8968
rect 255222 8888 255228 8900
rect 255102 8860 255228 8888
rect 255222 8848 255228 8860
rect 255280 8848 255286 8900
rect 302878 8440 302884 8492
rect 302936 8480 302942 8492
rect 395614 8480 395620 8492
rect 302936 8452 395620 8480
rect 302936 8440 302942 8452
rect 395614 8440 395620 8452
rect 395672 8440 395678 8492
rect 293770 8372 293776 8424
rect 293828 8412 293834 8424
rect 387150 8412 387156 8424
rect 293828 8384 387156 8412
rect 293828 8372 293834 8384
rect 387150 8372 387156 8384
rect 387208 8372 387214 8424
rect 308398 8304 308404 8356
rect 308456 8344 308462 8356
rect 403986 8344 403992 8356
rect 308456 8316 403992 8344
rect 308456 8304 308462 8316
rect 403986 8304 403992 8316
rect 404044 8304 404050 8356
rect 362494 7692 362500 7744
rect 362552 7732 362558 7744
rect 408310 7732 408316 7744
rect 362552 7704 408316 7732
rect 362552 7692 362558 7704
rect 408310 7692 408316 7704
rect 408368 7692 408374 7744
rect 1104 7642 528816 7664
rect 1104 7590 67574 7642
rect 67626 7590 67638 7642
rect 67690 7590 67702 7642
rect 67754 7590 67766 7642
rect 67818 7590 67830 7642
rect 67882 7590 199502 7642
rect 199554 7590 199566 7642
rect 199618 7590 199630 7642
rect 199682 7590 199694 7642
rect 199746 7590 199758 7642
rect 199810 7590 331430 7642
rect 331482 7590 331494 7642
rect 331546 7590 331558 7642
rect 331610 7590 331622 7642
rect 331674 7590 331686 7642
rect 331738 7590 463358 7642
rect 463410 7590 463422 7642
rect 463474 7590 463486 7642
rect 463538 7590 463550 7642
rect 463602 7590 463614 7642
rect 463666 7590 528816 7642
rect 1104 7568 528816 7590
rect 319622 7488 319628 7540
rect 319680 7528 319686 7540
rect 404538 7528 404544 7540
rect 319680 7500 404544 7528
rect 319680 7488 319686 7500
rect 404538 7488 404544 7500
rect 404596 7488 404602 7540
rect 218514 7420 218520 7472
rect 218572 7460 218578 7472
rect 306650 7460 306656 7472
rect 218572 7432 306656 7460
rect 218572 7420 218578 7432
rect 306650 7420 306656 7432
rect 306708 7420 306714 7472
rect 314746 7420 314752 7472
rect 314804 7460 314810 7472
rect 403710 7460 403716 7472
rect 314804 7432 403716 7460
rect 314804 7420 314810 7432
rect 403710 7420 403716 7432
rect 403768 7420 403774 7472
rect 219526 7352 219532 7404
rect 219584 7392 219590 7404
rect 300210 7392 300216 7404
rect 219584 7364 300216 7392
rect 219584 7352 219590 7364
rect 300210 7352 300216 7364
rect 300268 7352 300274 7404
rect 315942 7352 315948 7404
rect 316000 7392 316006 7404
rect 407206 7392 407212 7404
rect 316000 7364 407212 7392
rect 316000 7352 316006 7364
rect 407206 7352 407212 7364
rect 407264 7352 407270 7404
rect 220446 7284 220452 7336
rect 220504 7324 220510 7336
rect 301406 7324 301412 7336
rect 220504 7296 301412 7324
rect 220504 7284 220510 7296
rect 301406 7284 301412 7296
rect 301464 7284 301470 7336
rect 310698 7284 310704 7336
rect 310756 7324 310762 7336
rect 403066 7324 403072 7336
rect 310756 7296 403072 7324
rect 310756 7284 310762 7296
rect 403066 7284 403072 7296
rect 403124 7284 403130 7336
rect 202782 7216 202788 7268
rect 202840 7256 202846 7268
rect 296530 7256 296536 7268
rect 202840 7228 296536 7256
rect 202840 7216 202846 7228
rect 296530 7216 296536 7228
rect 296588 7216 296594 7268
rect 303430 7216 303436 7268
rect 303488 7256 303494 7268
rect 396718 7256 396724 7268
rect 303488 7228 396724 7256
rect 303488 7216 303494 7228
rect 396718 7216 396724 7228
rect 396776 7216 396782 7268
rect 31294 7148 31300 7200
rect 31352 7188 31358 7200
rect 125410 7188 125416 7200
rect 31352 7160 125416 7188
rect 31352 7148 31358 7160
rect 125410 7148 125416 7160
rect 125468 7148 125474 7200
rect 125870 7148 125876 7200
rect 125928 7188 125934 7200
rect 218698 7188 218704 7200
rect 125928 7160 218704 7188
rect 125928 7148 125934 7160
rect 218698 7148 218704 7160
rect 218756 7148 218762 7200
rect 291102 7148 291108 7200
rect 291160 7188 291166 7200
rect 385310 7188 385316 7200
rect 291160 7160 385316 7188
rect 291160 7148 291166 7160
rect 385310 7148 385316 7160
rect 385368 7148 385374 7200
rect 1104 7098 528816 7120
rect 1104 7046 66914 7098
rect 66966 7046 66978 7098
rect 67030 7046 67042 7098
rect 67094 7046 67106 7098
rect 67158 7046 67170 7098
rect 67222 7046 198842 7098
rect 198894 7046 198906 7098
rect 198958 7046 198970 7098
rect 199022 7046 199034 7098
rect 199086 7046 199098 7098
rect 199150 7046 330770 7098
rect 330822 7046 330834 7098
rect 330886 7046 330898 7098
rect 330950 7046 330962 7098
rect 331014 7046 331026 7098
rect 331078 7046 462698 7098
rect 462750 7046 462762 7098
rect 462814 7046 462826 7098
rect 462878 7046 462890 7098
rect 462942 7046 462954 7098
rect 463006 7046 528816 7098
rect 1104 7024 528816 7046
rect 125134 6944 125140 6996
rect 125192 6984 125198 6996
rect 217134 6984 217140 6996
rect 125192 6956 217140 6984
rect 125192 6944 125198 6956
rect 217134 6944 217140 6956
rect 217192 6944 217198 6996
rect 218054 6944 218060 6996
rect 218112 6984 218118 6996
rect 314286 6984 314292 6996
rect 218112 6956 314292 6984
rect 218112 6944 218118 6956
rect 314286 6944 314292 6956
rect 314344 6944 314350 6996
rect 318334 6944 318340 6996
rect 318392 6984 318398 6996
rect 411806 6984 411812 6996
rect 318392 6956 411812 6984
rect 318392 6944 318398 6956
rect 411806 6944 411812 6956
rect 411864 6944 411870 6996
rect 124490 6876 124496 6928
rect 124548 6916 124554 6928
rect 218882 6916 218888 6928
rect 124548 6888 218888 6916
rect 124548 6876 124554 6888
rect 218882 6876 218888 6888
rect 218940 6876 218946 6928
rect 304718 6876 304724 6928
rect 304776 6916 304782 6928
rect 402054 6916 402060 6928
rect 304776 6888 402060 6916
rect 304776 6876 304782 6888
rect 402054 6876 402060 6888
rect 402112 6876 402118 6928
rect 17862 6808 17868 6860
rect 17920 6848 17926 6860
rect 19886 6848 19892 6860
rect 17920 6820 19892 6848
rect 17920 6808 17926 6820
rect 19886 6808 19892 6820
rect 19944 6808 19950 6860
rect 34422 6808 34428 6860
rect 34480 6848 34486 6860
rect 37642 6848 37648 6860
rect 34480 6820 37648 6848
rect 34480 6808 34486 6820
rect 37642 6808 37648 6820
rect 37700 6808 37706 6860
rect 52362 6808 52368 6860
rect 52420 6848 52426 6860
rect 53834 6848 53840 6860
rect 52420 6820 53840 6848
rect 52420 6808 52426 6820
rect 53834 6808 53840 6820
rect 53892 6808 53898 6860
rect 68922 6808 68928 6860
rect 68980 6848 68986 6860
rect 73982 6848 73988 6860
rect 68980 6820 73988 6848
rect 68980 6808 68986 6820
rect 73982 6808 73988 6820
rect 74040 6808 74046 6860
rect 85482 6808 85488 6860
rect 85540 6848 85546 6860
rect 92014 6848 92020 6860
rect 85540 6820 92020 6848
rect 85540 6808 85546 6820
rect 92014 6808 92020 6820
rect 92072 6808 92078 6860
rect 119982 6808 119988 6860
rect 120040 6848 120046 6860
rect 126790 6848 126796 6860
rect 120040 6820 126796 6848
rect 120040 6808 120046 6820
rect 126790 6808 126796 6820
rect 126848 6808 126854 6860
rect 1104 6554 528816 6576
rect 1104 6502 67574 6554
rect 67626 6502 67638 6554
rect 67690 6502 67702 6554
rect 67754 6502 67766 6554
rect 67818 6502 67830 6554
rect 67882 6502 199502 6554
rect 199554 6502 199566 6554
rect 199618 6502 199630 6554
rect 199682 6502 199694 6554
rect 199746 6502 199758 6554
rect 199810 6502 331430 6554
rect 331482 6502 331494 6554
rect 331546 6502 331558 6554
rect 331610 6502 331622 6554
rect 331674 6502 331686 6554
rect 331738 6502 463358 6554
rect 463410 6502 463422 6554
rect 463474 6502 463486 6554
rect 463538 6502 463550 6554
rect 463602 6502 463614 6554
rect 463666 6502 528816 6554
rect 1104 6480 528816 6502
rect 300854 6264 300860 6316
rect 300912 6304 300918 6316
rect 351914 6304 351920 6316
rect 300912 6276 351920 6304
rect 300912 6264 300918 6276
rect 351914 6264 351920 6276
rect 351972 6264 351978 6316
rect 114186 6196 114192 6248
rect 114244 6236 114250 6248
rect 208578 6236 208584 6248
rect 114244 6208 208584 6236
rect 114244 6196 114250 6208
rect 208578 6196 208584 6208
rect 208636 6196 208642 6248
rect 209406 6196 209412 6248
rect 209464 6236 209470 6248
rect 306098 6236 306104 6248
rect 209464 6208 306104 6236
rect 209464 6196 209470 6208
rect 306098 6196 306104 6208
rect 306156 6196 306162 6248
rect 324222 6196 324228 6248
rect 324280 6236 324286 6248
rect 341978 6236 341984 6248
rect 324280 6208 341984 6236
rect 324280 6196 324286 6208
rect 341978 6196 341984 6208
rect 342036 6196 342042 6248
rect 357250 6196 357256 6248
rect 357308 6236 357314 6248
rect 380526 6236 380532 6248
rect 357308 6208 380532 6236
rect 357308 6196 357314 6208
rect 380526 6196 380532 6208
rect 380584 6196 380590 6248
rect 391842 6196 391848 6248
rect 391900 6236 391906 6248
rect 416314 6236 416320 6248
rect 391900 6208 416320 6236
rect 391900 6196 391906 6208
rect 416314 6196 416320 6208
rect 416372 6196 416378 6248
rect 426342 6196 426348 6248
rect 426400 6236 426406 6248
rect 442810 6236 442816 6248
rect 426400 6208 442816 6236
rect 426400 6196 426406 6208
rect 442810 6196 442816 6208
rect 442868 6196 442874 6248
rect 102226 6128 102232 6180
rect 102284 6168 102290 6180
rect 110046 6168 110052 6180
rect 102284 6140 110052 6168
rect 102284 6128 102290 6140
rect 110046 6128 110052 6140
rect 110104 6128 110110 6180
rect 136542 6128 136548 6180
rect 136600 6168 136606 6180
rect 145834 6168 145840 6180
rect 136600 6140 145840 6168
rect 136600 6128 136606 6140
rect 145834 6128 145840 6140
rect 145892 6128 145898 6180
rect 153102 6128 153108 6180
rect 153160 6168 153166 6180
rect 164142 6168 164148 6180
rect 153160 6140 164148 6168
rect 153160 6128 153166 6140
rect 164142 6128 164148 6140
rect 164200 6128 164206 6180
rect 171042 6128 171048 6180
rect 171100 6168 171106 6180
rect 179414 6168 179420 6180
rect 171100 6140 179420 6168
rect 171100 6128 171106 6140
rect 179414 6128 179420 6140
rect 179472 6128 179478 6180
rect 187602 6128 187608 6180
rect 187660 6168 187666 6180
rect 200206 6168 200212 6180
rect 187660 6140 200212 6168
rect 187660 6128 187666 6140
rect 200206 6128 200212 6140
rect 200264 6128 200270 6180
rect 204162 6128 204168 6180
rect 204220 6168 204226 6180
rect 217410 6168 217416 6180
rect 204220 6140 217416 6168
rect 204220 6128 204226 6140
rect 217410 6128 217416 6140
rect 217468 6128 217474 6180
rect 222102 6128 222108 6180
rect 222160 6168 222166 6180
rect 236270 6168 236276 6180
rect 222160 6140 236276 6168
rect 222160 6128 222166 6140
rect 236270 6128 236276 6140
rect 236328 6128 236334 6180
rect 238662 6128 238668 6180
rect 238720 6168 238726 6180
rect 254026 6168 254032 6180
rect 238720 6140 254032 6168
rect 238720 6128 238726 6140
rect 254026 6128 254032 6140
rect 254084 6128 254090 6180
rect 255222 6128 255228 6180
rect 255280 6168 255286 6180
rect 271782 6168 271788 6180
rect 255280 6140 271788 6168
rect 255280 6128 255286 6140
rect 271782 6128 271788 6140
rect 271840 6128 271846 6180
rect 273162 6128 273168 6180
rect 273220 6168 273226 6180
rect 288342 6168 288348 6180
rect 273220 6140 288348 6168
rect 273220 6128 273226 6140
rect 288342 6128 288348 6140
rect 288400 6128 288406 6180
rect 289446 6128 289452 6180
rect 289504 6168 289510 6180
rect 304994 6168 305000 6180
rect 289504 6140 305000 6168
rect 289504 6128 289510 6140
rect 304994 6128 305000 6140
rect 305052 6128 305058 6180
rect 306282 6128 306288 6180
rect 306340 6168 306346 6180
rect 326430 6168 326436 6180
rect 306340 6140 326436 6168
rect 306340 6128 306346 6140
rect 326430 6128 326436 6140
rect 326488 6128 326494 6180
rect 340782 6128 340788 6180
rect 340840 6168 340846 6180
rect 362218 6168 362224 6180
rect 340840 6140 362224 6168
rect 340840 6128 340846 6140
rect 362218 6128 362224 6140
rect 362276 6128 362282 6180
rect 375282 6128 375288 6180
rect 375340 6168 375346 6180
rect 398558 6168 398564 6180
rect 375340 6140 398564 6168
rect 375340 6128 375346 6140
rect 398558 6128 398564 6140
rect 398616 6128 398622 6180
rect 408402 6128 408408 6180
rect 408460 6168 408466 6180
rect 434622 6168 434628 6180
rect 408460 6140 434628 6168
rect 408460 6128 408466 6140
rect 434622 6128 434628 6140
rect 434680 6128 434686 6180
rect 442902 6128 442908 6180
rect 442960 6168 442966 6180
rect 470410 6168 470416 6180
rect 442960 6140 470416 6168
rect 442960 6128 442966 6140
rect 470410 6128 470416 6140
rect 470468 6128 470474 6180
rect 27706 6060 27712 6112
rect 27764 6100 27770 6112
rect 120258 6100 120264 6112
rect 27764 6072 120264 6100
rect 27764 6060 27770 6072
rect 120258 6060 120264 6072
rect 120316 6060 120322 6112
rect 126238 6060 126244 6112
rect 126296 6100 126302 6112
rect 219158 6100 219164 6112
rect 126296 6072 219164 6100
rect 126296 6060 126302 6072
rect 219158 6060 219164 6072
rect 219216 6060 219222 6112
rect 304810 6060 304816 6112
rect 304868 6100 304874 6112
rect 355778 6100 355784 6112
rect 304868 6072 355784 6100
rect 304868 6060 304874 6072
rect 355778 6060 355784 6072
rect 355836 6060 355842 6112
rect 1104 6010 528816 6032
rect 1104 5958 66914 6010
rect 66966 5958 66978 6010
rect 67030 5958 67042 6010
rect 67094 5958 67106 6010
rect 67158 5958 67170 6010
rect 67222 5958 198842 6010
rect 198894 5958 198906 6010
rect 198958 5958 198970 6010
rect 199022 5958 199034 6010
rect 199086 5958 199098 6010
rect 199150 5958 330770 6010
rect 330822 5958 330834 6010
rect 330886 5958 330898 6010
rect 330950 5958 330962 6010
rect 331014 5958 331026 6010
rect 331078 5958 462698 6010
rect 462750 5958 462762 6010
rect 462814 5958 462826 6010
rect 462878 5958 462890 6010
rect 462942 5958 462954 6010
rect 463006 5958 528816 6010
rect 1104 5936 528816 5958
rect 29730 5856 29736 5908
rect 29788 5896 29794 5908
rect 123846 5896 123852 5908
rect 29788 5868 123852 5896
rect 29788 5856 29794 5868
rect 123846 5856 123852 5868
rect 123904 5856 123910 5908
rect 169202 5856 169208 5908
rect 169260 5896 169266 5908
rect 262306 5896 262312 5908
rect 169260 5868 262312 5896
rect 169260 5856 169266 5868
rect 262306 5856 262312 5868
rect 262364 5856 262370 5908
rect 263502 5856 263508 5908
rect 263560 5896 263566 5908
rect 340874 5896 340880 5908
rect 263560 5868 340880 5896
rect 263560 5856 263566 5868
rect 340874 5856 340880 5868
rect 340932 5856 340938 5908
rect 355134 5856 355140 5908
rect 355192 5896 355198 5908
rect 409966 5896 409972 5908
rect 355192 5868 409972 5896
rect 355192 5856 355198 5868
rect 409966 5856 409972 5868
rect 410024 5856 410030 5908
rect 117314 5788 117320 5840
rect 117372 5828 117378 5840
rect 207658 5828 207664 5840
rect 117372 5800 207664 5828
rect 117372 5788 117378 5800
rect 207658 5788 207664 5800
rect 207716 5788 207722 5840
rect 209038 5788 209044 5840
rect 209096 5828 209102 5840
rect 303798 5828 303804 5840
rect 209096 5800 303804 5828
rect 209096 5788 209102 5800
rect 303798 5788 303804 5800
rect 303856 5788 303862 5840
rect 342346 5788 342352 5840
rect 342404 5828 342410 5840
rect 407758 5828 407764 5840
rect 342404 5800 407764 5828
rect 342404 5788 342410 5800
rect 407758 5788 407764 5800
rect 407816 5788 407822 5840
rect 26418 5720 26424 5772
rect 26476 5760 26482 5772
rect 120074 5760 120080 5772
rect 26476 5732 120080 5760
rect 26476 5720 26482 5732
rect 120074 5720 120080 5732
rect 120132 5720 120138 5772
rect 212810 5720 212816 5772
rect 212868 5760 212874 5772
rect 308122 5760 308128 5772
rect 212868 5732 308128 5760
rect 212868 5720 212874 5732
rect 308122 5720 308128 5732
rect 308180 5720 308186 5772
rect 338022 5720 338028 5772
rect 338080 5760 338086 5772
rect 407114 5760 407120 5772
rect 338080 5732 407120 5760
rect 338080 5720 338086 5732
rect 407114 5720 407120 5732
rect 407172 5720 407178 5772
rect 117406 5652 117412 5704
rect 117464 5692 117470 5704
rect 208854 5692 208860 5704
rect 117464 5664 208860 5692
rect 117464 5652 117470 5664
rect 208854 5652 208860 5664
rect 208912 5652 208918 5704
rect 209590 5652 209596 5704
rect 209648 5692 209654 5704
rect 305270 5692 305276 5704
rect 209648 5664 305276 5692
rect 209648 5652 209654 5664
rect 305270 5652 305276 5664
rect 305328 5652 305334 5704
rect 332502 5652 332508 5704
rect 332560 5692 332566 5704
rect 406102 5692 406108 5704
rect 332560 5664 406108 5692
rect 332560 5652 332566 5664
rect 406102 5652 406108 5664
rect 406160 5652 406166 5704
rect 24578 5584 24584 5636
rect 24636 5624 24642 5636
rect 118786 5624 118792 5636
rect 24636 5596 118792 5624
rect 24636 5584 24642 5596
rect 118786 5584 118792 5596
rect 118844 5584 118850 5636
rect 119338 5584 119344 5636
rect 119396 5624 119402 5636
rect 213362 5624 213368 5636
rect 119396 5596 213368 5624
rect 119396 5584 119402 5596
rect 213362 5584 213368 5596
rect 213420 5584 213426 5636
rect 298646 5584 298652 5636
rect 298704 5624 298710 5636
rect 390186 5624 390192 5636
rect 298704 5596 390192 5624
rect 298704 5584 298710 5596
rect 390186 5584 390192 5596
rect 390244 5584 390250 5636
rect 25406 5516 25412 5568
rect 25464 5556 25470 5568
rect 118694 5556 118700 5568
rect 25464 5528 118700 5556
rect 25464 5516 25470 5528
rect 118694 5516 118700 5528
rect 118752 5516 118758 5568
rect 208394 5516 208400 5568
rect 208452 5556 208458 5568
rect 305362 5556 305368 5568
rect 208452 5528 305368 5556
rect 208452 5516 208458 5528
rect 305362 5516 305368 5528
rect 305420 5516 305426 5568
rect 327166 5516 327172 5568
rect 327224 5556 327230 5568
rect 421374 5556 421380 5568
rect 327224 5528 421380 5556
rect 327224 5516 327230 5528
rect 421374 5516 421380 5528
rect 421432 5516 421438 5568
rect 1104 5466 528816 5488
rect 1104 5414 67574 5466
rect 67626 5414 67638 5466
rect 67690 5414 67702 5466
rect 67754 5414 67766 5466
rect 67818 5414 67830 5466
rect 67882 5414 199502 5466
rect 199554 5414 199566 5466
rect 199618 5414 199630 5466
rect 199682 5414 199694 5466
rect 199746 5414 199758 5466
rect 199810 5414 331430 5466
rect 331482 5414 331494 5466
rect 331546 5414 331558 5466
rect 331610 5414 331622 5466
rect 331674 5414 331686 5466
rect 331738 5414 463358 5466
rect 463410 5414 463422 5466
rect 463474 5414 463486 5466
rect 463538 5414 463550 5466
rect 463602 5414 463614 5466
rect 463666 5414 528816 5466
rect 1104 5392 528816 5414
rect 110782 5176 110788 5228
rect 110840 5216 110846 5228
rect 204898 5216 204904 5228
rect 110840 5188 204904 5216
rect 110840 5176 110846 5188
rect 204898 5176 204904 5188
rect 204956 5176 204962 5228
rect 213638 5176 213644 5228
rect 213696 5216 213702 5228
rect 218146 5216 218152 5228
rect 213696 5188 218152 5216
rect 213696 5176 213702 5188
rect 218146 5176 218152 5188
rect 218204 5176 218210 5228
rect 63586 5108 63592 5160
rect 63644 5148 63650 5160
rect 150986 5148 150992 5160
rect 63644 5120 150992 5148
rect 63644 5108 63650 5120
rect 150986 5108 150992 5120
rect 151044 5108 151050 5160
rect 214466 5108 214472 5160
rect 214524 5148 214530 5160
rect 220354 5148 220360 5160
rect 214524 5120 220360 5148
rect 214524 5108 214530 5120
rect 220354 5108 220360 5120
rect 220412 5108 220418 5160
rect 239030 5108 239036 5160
rect 239088 5148 239094 5160
rect 332318 5148 332324 5160
rect 239088 5120 332324 5148
rect 239088 5108 239094 5120
rect 332318 5108 332324 5120
rect 332376 5108 332382 5160
rect 137278 5040 137284 5092
rect 137336 5080 137342 5092
rect 230750 5080 230756 5092
rect 137336 5052 230756 5080
rect 137336 5040 137342 5052
rect 230750 5040 230756 5052
rect 230808 5040 230814 5092
rect 308490 5040 308496 5092
rect 308548 5080 308554 5092
rect 355870 5080 355876 5092
rect 308548 5052 355876 5080
rect 308548 5040 308554 5052
rect 355870 5040 355876 5052
rect 355928 5040 355934 5092
rect 116210 4972 116216 5024
rect 116268 4972 116274 5024
rect 116670 4972 116676 5024
rect 116728 5012 116734 5024
rect 116857 5015 116915 5021
rect 116857 5012 116869 5015
rect 116728 4984 116869 5012
rect 116728 4972 116734 4984
rect 116857 4981 116869 4984
rect 116903 4981 116915 5015
rect 116857 4975 116915 4981
rect 117498 4972 117504 5024
rect 117556 4972 117562 5024
rect 118050 4972 118056 5024
rect 118108 5012 118114 5024
rect 118237 5015 118295 5021
rect 118237 5012 118249 5015
rect 118108 4984 118249 5012
rect 118108 4972 118114 4984
rect 118237 4981 118249 4984
rect 118283 4981 118295 5015
rect 118237 4975 118295 4981
rect 210786 4972 210792 5024
rect 210844 5012 210850 5024
rect 210973 5015 211031 5021
rect 210973 5012 210985 5015
rect 210844 4984 210985 5012
rect 210844 4972 210850 4984
rect 210973 4981 210985 4984
rect 211019 4981 211031 5015
rect 210973 4975 211031 4981
rect 211614 4972 211620 5024
rect 211672 4972 211678 5024
rect 214282 4972 214288 5024
rect 214340 4972 214346 5024
rect 214834 4972 214840 5024
rect 214892 4972 214898 5024
rect 215386 4972 215392 5024
rect 215444 4972 215450 5024
rect 216214 4972 216220 5024
rect 216272 4972 216278 5024
rect 216769 5015 216827 5021
rect 216769 4981 216781 5015
rect 216815 5012 216827 5015
rect 216858 5012 216864 5024
rect 216815 4984 216864 5012
rect 216815 4981 216827 4984
rect 216769 4975 216827 4981
rect 216858 4972 216864 4984
rect 216916 4972 216922 5024
rect 221090 4972 221096 5024
rect 221148 5012 221154 5024
rect 295426 5012 295432 5024
rect 221148 4984 295432 5012
rect 221148 4972 221154 4984
rect 295426 4972 295432 4984
rect 295484 4972 295490 5024
rect 306006 4972 306012 5024
rect 306064 5012 306070 5024
rect 306193 5015 306251 5021
rect 306193 5012 306205 5015
rect 306064 4984 306205 5012
rect 306064 4972 306070 4984
rect 306193 4981 306205 4984
rect 306239 4981 306251 5015
rect 306193 4975 306251 4981
rect 306742 4972 306748 5024
rect 306800 4972 306806 5024
rect 307570 4972 307576 5024
rect 307628 4972 307634 5024
rect 307846 4972 307852 5024
rect 307904 5012 307910 5024
rect 308033 5015 308091 5021
rect 308033 5012 308045 5015
rect 307904 4984 308045 5012
rect 307904 4972 307910 4984
rect 308033 4981 308045 4984
rect 308079 4981 308091 5015
rect 308033 4975 308091 4981
rect 308582 4972 308588 5024
rect 308640 5012 308646 5024
rect 308677 5015 308735 5021
rect 308677 5012 308689 5015
rect 308640 4984 308689 5012
rect 308640 4972 308646 4984
rect 308677 4981 308689 4984
rect 308723 4981 308735 5015
rect 308677 4975 308735 4981
rect 357434 4972 357440 5024
rect 357492 5012 357498 5024
rect 402330 5012 402336 5024
rect 357492 4984 402336 5012
rect 357492 4972 357498 4984
rect 402330 4972 402336 4984
rect 402388 4972 402394 5024
rect 1104 4922 528816 4944
rect 1104 4870 66914 4922
rect 66966 4870 66978 4922
rect 67030 4870 67042 4922
rect 67094 4870 67106 4922
rect 67158 4870 67170 4922
rect 67222 4870 198842 4922
rect 198894 4870 198906 4922
rect 198958 4870 198970 4922
rect 199022 4870 199034 4922
rect 199086 4870 199098 4922
rect 199150 4870 330770 4922
rect 330822 4870 330834 4922
rect 330886 4870 330898 4922
rect 330950 4870 330962 4922
rect 331014 4870 331026 4922
rect 331078 4870 462698 4922
rect 462750 4870 462762 4922
rect 462814 4870 462826 4922
rect 462878 4870 462890 4922
rect 462942 4870 462954 4922
rect 463006 4870 528816 4922
rect 1104 4848 528816 4870
rect 63494 4768 63500 4820
rect 63552 4808 63558 4820
rect 156690 4808 156696 4820
rect 63552 4780 156696 4808
rect 63552 4768 63558 4780
rect 156690 4768 156696 4780
rect 156748 4768 156754 4820
rect 211522 4768 211528 4820
rect 211580 4808 211586 4820
rect 301130 4808 301136 4820
rect 211580 4780 301136 4808
rect 211580 4768 211586 4780
rect 301130 4768 301136 4780
rect 301188 4768 301194 4820
rect 308490 4768 308496 4820
rect 308548 4768 308554 4820
rect 350534 4768 350540 4820
rect 350592 4808 350598 4820
rect 403802 4808 403808 4820
rect 350592 4780 403808 4808
rect 350592 4768 350598 4780
rect 403802 4768 403808 4780
rect 403860 4768 403866 4820
rect 442810 4768 442816 4820
rect 442868 4808 442874 4820
rect 452654 4808 452660 4820
rect 442868 4780 452660 4808
rect 442868 4768 442874 4780
rect 452654 4768 452660 4780
rect 452712 4768 452718 4820
rect 131390 4700 131396 4752
rect 131448 4740 131454 4752
rect 224954 4740 224960 4752
rect 131448 4712 224960 4740
rect 131448 4700 131454 4712
rect 224954 4700 224960 4712
rect 225012 4700 225018 4752
rect 260006 4700 260012 4752
rect 260064 4740 260070 4752
rect 350718 4740 350724 4752
rect 260064 4712 350724 4740
rect 260064 4700 260070 4712
rect 350718 4700 350724 4712
rect 350776 4700 350782 4752
rect 353294 4700 353300 4752
rect 353352 4740 353358 4752
rect 407298 4740 407304 4752
rect 353352 4712 407304 4740
rect 353352 4700 353358 4712
rect 407298 4700 407304 4712
rect 407356 4700 407362 4752
rect 126422 4632 126428 4684
rect 126480 4672 126486 4684
rect 219894 4672 219900 4684
rect 126480 4644 219900 4672
rect 126480 4632 126486 4644
rect 219894 4632 219900 4644
rect 219952 4632 219958 4684
rect 220998 4632 221004 4684
rect 221056 4672 221062 4684
rect 314010 4672 314016 4684
rect 221056 4644 314016 4672
rect 221056 4632 221062 4644
rect 314010 4632 314016 4644
rect 314068 4632 314074 4684
rect 325326 4632 325332 4684
rect 325384 4672 325390 4684
rect 405274 4672 405280 4684
rect 325384 4644 405280 4672
rect 325384 4632 325390 4644
rect 405274 4632 405280 4644
rect 405332 4632 405338 4684
rect 28350 4564 28356 4616
rect 28408 4604 28414 4616
rect 120626 4604 120632 4616
rect 28408 4576 120632 4604
rect 28408 4564 28414 4576
rect 120626 4564 120632 4576
rect 120684 4564 120690 4616
rect 143902 4564 143908 4616
rect 143960 4604 143966 4616
rect 237742 4604 237748 4616
rect 143960 4576 237748 4604
rect 143960 4564 143966 4576
rect 237742 4564 237748 4576
rect 237800 4564 237806 4616
rect 307754 4564 307760 4616
rect 307812 4604 307818 4616
rect 308309 4607 308367 4613
rect 308309 4604 308321 4607
rect 307812 4576 308321 4604
rect 307812 4564 307818 4576
rect 308309 4573 308321 4576
rect 308355 4573 308367 4607
rect 308309 4567 308367 4573
rect 330018 4564 330024 4616
rect 330076 4604 330082 4616
rect 405918 4604 405924 4616
rect 330076 4576 405924 4604
rect 330076 4564 330082 4576
rect 405918 4564 405924 4576
rect 405976 4564 405982 4616
rect 23382 4496 23388 4548
rect 23440 4536 23446 4548
rect 58158 4536 58164 4548
rect 23440 4508 58164 4536
rect 23440 4496 23446 4508
rect 58158 4496 58164 4508
rect 58216 4496 58222 4548
rect 126606 4496 126612 4548
rect 126664 4536 126670 4548
rect 214466 4536 214472 4548
rect 126664 4508 214472 4536
rect 126664 4496 126670 4508
rect 214466 4496 214472 4508
rect 214524 4496 214530 4548
rect 215478 4496 215484 4548
rect 215536 4536 215542 4548
rect 215757 4539 215815 4545
rect 215757 4536 215769 4539
rect 215536 4508 215769 4536
rect 215536 4496 215542 4508
rect 215757 4505 215769 4508
rect 215803 4536 215815 4539
rect 217318 4536 217324 4548
rect 215803 4508 217324 4536
rect 215803 4505 215815 4508
rect 215757 4499 215815 4505
rect 217318 4496 217324 4508
rect 217376 4496 217382 4548
rect 287422 4496 287428 4548
rect 287480 4536 287486 4548
rect 381262 4536 381268 4548
rect 287480 4508 381268 4536
rect 287480 4496 287486 4508
rect 381262 4496 381268 4508
rect 381320 4496 381326 4548
rect 115477 4471 115535 4477
rect 115477 4437 115489 4471
rect 115523 4468 115535 4471
rect 115658 4468 115664 4480
rect 115523 4440 115664 4468
rect 115523 4437 115535 4440
rect 115477 4431 115535 4437
rect 115658 4428 115664 4440
rect 115716 4428 115722 4480
rect 116026 4428 116032 4480
rect 116084 4428 116090 4480
rect 116578 4428 116584 4480
rect 116636 4428 116642 4480
rect 117866 4428 117872 4480
rect 117924 4428 117930 4480
rect 118418 4428 118424 4480
rect 118476 4428 118482 4480
rect 118970 4428 118976 4480
rect 119028 4428 119034 4480
rect 119522 4428 119528 4480
rect 119580 4428 119586 4480
rect 120718 4428 120724 4480
rect 120776 4428 120782 4480
rect 121362 4428 121368 4480
rect 121420 4428 121426 4480
rect 122374 4428 122380 4480
rect 122432 4468 122438 4480
rect 122469 4471 122527 4477
rect 122469 4468 122481 4471
rect 122432 4440 122481 4468
rect 122432 4428 122438 4440
rect 122469 4437 122481 4440
rect 122515 4437 122527 4471
rect 122469 4431 122527 4437
rect 210418 4428 210424 4480
rect 210476 4428 210482 4480
rect 211062 4428 211068 4480
rect 211120 4428 211126 4480
rect 211617 4471 211675 4477
rect 211617 4437 211629 4471
rect 211663 4468 211675 4471
rect 211706 4468 211712 4480
rect 211663 4440 211712 4468
rect 211663 4437 211675 4440
rect 211617 4431 211675 4437
rect 211706 4428 211712 4440
rect 211764 4428 211770 4480
rect 212166 4428 212172 4480
rect 212224 4468 212230 4480
rect 212353 4471 212411 4477
rect 212353 4468 212365 4471
rect 212224 4440 212365 4468
rect 212224 4428 212230 4440
rect 212353 4437 212365 4440
rect 212399 4437 212411 4471
rect 212353 4431 212411 4437
rect 212997 4471 213055 4477
rect 212997 4437 213009 4471
rect 213043 4468 213055 4471
rect 213178 4468 213184 4480
rect 213043 4440 213184 4468
rect 213043 4437 213055 4440
rect 212997 4431 213055 4437
rect 213178 4428 213184 4440
rect 213236 4428 213242 4480
rect 213546 4428 213552 4480
rect 213604 4428 213610 4480
rect 213914 4428 213920 4480
rect 213972 4468 213978 4480
rect 214009 4471 214067 4477
rect 214009 4468 214021 4471
rect 213972 4440 214021 4468
rect 213972 4428 213978 4440
rect 214009 4437 214021 4440
rect 214055 4437 214067 4471
rect 214009 4431 214067 4437
rect 214653 4471 214711 4477
rect 214653 4437 214665 4471
rect 214699 4468 214711 4471
rect 215202 4468 215208 4480
rect 214699 4440 215208 4468
rect 214699 4437 214711 4440
rect 214653 4431 214711 4437
rect 215202 4428 215208 4440
rect 215260 4428 215266 4480
rect 216766 4428 216772 4480
rect 216824 4428 216830 4480
rect 217226 4428 217232 4480
rect 217284 4428 217290 4480
rect 217873 4471 217931 4477
rect 217873 4437 217885 4471
rect 217919 4468 217931 4471
rect 217962 4468 217968 4480
rect 217919 4440 217968 4468
rect 217919 4437 217931 4440
rect 217873 4431 217931 4437
rect 217962 4428 217968 4440
rect 218020 4428 218026 4480
rect 220078 4428 220084 4480
rect 220136 4468 220142 4480
rect 304166 4468 304172 4480
rect 220136 4440 304172 4468
rect 220136 4428 220142 4440
rect 304166 4428 304172 4440
rect 304224 4428 304230 4480
rect 305546 4428 305552 4480
rect 305604 4468 305610 4480
rect 305641 4471 305699 4477
rect 305641 4468 305653 4471
rect 305604 4440 305653 4468
rect 305604 4428 305610 4440
rect 305641 4437 305653 4440
rect 305687 4437 305699 4471
rect 305641 4431 305699 4437
rect 306190 4428 306196 4480
rect 306248 4428 306254 4480
rect 306374 4428 306380 4480
rect 306432 4468 306438 4480
rect 306745 4471 306803 4477
rect 306745 4468 306757 4471
rect 306432 4440 306757 4468
rect 306432 4428 306438 4440
rect 306745 4437 306757 4440
rect 306791 4437 306803 4471
rect 306745 4431 306803 4437
rect 306834 4428 306840 4480
rect 306892 4468 306898 4480
rect 307389 4471 307447 4477
rect 307389 4468 307401 4471
rect 306892 4440 307401 4468
rect 306892 4428 306898 4440
rect 307389 4437 307401 4440
rect 307435 4468 307447 4471
rect 307662 4468 307668 4480
rect 307435 4440 307668 4468
rect 307435 4437 307447 4440
rect 307389 4431 307447 4437
rect 307662 4428 307668 4440
rect 307720 4428 307726 4480
rect 309137 4471 309195 4477
rect 309137 4437 309149 4471
rect 309183 4468 309195 4471
rect 309226 4468 309232 4480
rect 309183 4440 309232 4468
rect 309183 4437 309195 4440
rect 309137 4431 309195 4437
rect 309226 4428 309232 4440
rect 309284 4428 309290 4480
rect 309594 4428 309600 4480
rect 309652 4428 309658 4480
rect 310422 4428 310428 4480
rect 310480 4428 310486 4480
rect 349798 4428 349804 4480
rect 349856 4468 349862 4480
rect 406194 4468 406200 4480
rect 349856 4440 406200 4468
rect 349856 4428 349862 4440
rect 406194 4428 406200 4440
rect 406252 4428 406258 4480
rect 1104 4378 528816 4400
rect 1104 4326 67574 4378
rect 67626 4326 67638 4378
rect 67690 4326 67702 4378
rect 67754 4326 67766 4378
rect 67818 4326 67830 4378
rect 67882 4326 199502 4378
rect 199554 4326 199566 4378
rect 199618 4326 199630 4378
rect 199682 4326 199694 4378
rect 199746 4326 199758 4378
rect 199810 4326 331430 4378
rect 331482 4326 331494 4378
rect 331546 4326 331558 4378
rect 331610 4326 331622 4378
rect 331674 4326 331686 4378
rect 331738 4326 463358 4378
rect 463410 4326 463422 4378
rect 463474 4326 463486 4378
rect 463538 4326 463550 4378
rect 463602 4326 463614 4378
rect 463666 4326 528816 4378
rect 1104 4304 528816 4326
rect 22922 4224 22928 4276
rect 22980 4264 22986 4276
rect 116302 4264 116308 4276
rect 22980 4236 116308 4264
rect 22980 4224 22986 4236
rect 116302 4224 116308 4236
rect 116360 4224 116366 4276
rect 208118 4224 208124 4276
rect 208176 4264 208182 4276
rect 211522 4264 211528 4276
rect 208176 4236 211528 4264
rect 208176 4224 208182 4236
rect 211522 4224 211528 4236
rect 211580 4224 211586 4276
rect 297358 4264 297364 4276
rect 211632 4236 297364 4264
rect 20990 4156 20996 4208
rect 21048 4196 21054 4208
rect 70394 4196 70400 4208
rect 21048 4168 70400 4196
rect 21048 4156 21054 4168
rect 70394 4156 70400 4168
rect 70452 4156 70458 4208
rect 98638 4156 98644 4208
rect 98696 4196 98702 4208
rect 192202 4196 192208 4208
rect 98696 4168 192208 4196
rect 98696 4156 98702 4168
rect 192202 4156 192208 4168
rect 192260 4156 192266 4208
rect 203886 4156 203892 4208
rect 203944 4196 203950 4208
rect 211632 4196 211660 4236
rect 297358 4224 297364 4236
rect 297416 4224 297422 4276
rect 317874 4224 317880 4276
rect 317932 4264 317938 4276
rect 403894 4264 403900 4276
rect 317932 4236 403900 4264
rect 317932 4224 317938 4236
rect 403894 4224 403900 4236
rect 403952 4224 403958 4276
rect 203944 4168 211660 4196
rect 211801 4199 211859 4205
rect 203944 4156 203950 4168
rect 211801 4165 211813 4199
rect 211847 4196 211859 4199
rect 220078 4196 220084 4208
rect 211847 4168 220084 4196
rect 211847 4165 211859 4168
rect 211801 4159 211859 4165
rect 220078 4156 220084 4168
rect 220136 4156 220142 4208
rect 273070 4156 273076 4208
rect 273128 4196 273134 4208
rect 367278 4196 367284 4208
rect 273128 4168 367284 4196
rect 273128 4156 273134 4168
rect 367278 4156 367284 4168
rect 367336 4156 367342 4208
rect 388438 4156 388444 4208
rect 388496 4196 388502 4208
rect 481634 4196 481640 4208
rect 388496 4168 481640 4196
rect 388496 4156 388502 4168
rect 481634 4156 481640 4168
rect 481692 4156 481698 4208
rect 115750 4088 115756 4140
rect 115808 4088 115814 4140
rect 116578 4128 116584 4140
rect 115860 4100 116584 4128
rect 20714 4020 20720 4072
rect 20772 4060 20778 4072
rect 115201 4063 115259 4069
rect 115201 4060 115213 4063
rect 20772 4032 115213 4060
rect 20772 4020 20778 4032
rect 115201 4029 115213 4032
rect 115247 4029 115259 4063
rect 115201 4023 115259 4029
rect 115860 3992 115888 4100
rect 116578 4088 116584 4100
rect 116636 4128 116642 4140
rect 116857 4131 116915 4137
rect 116857 4128 116869 4131
rect 116636 4100 116869 4128
rect 116636 4088 116642 4100
rect 116857 4097 116869 4100
rect 116903 4097 116915 4131
rect 116857 4091 116915 4097
rect 118697 4131 118755 4137
rect 118697 4097 118709 4131
rect 118743 4128 118755 4131
rect 118970 4128 118976 4140
rect 118743 4100 118976 4128
rect 118743 4097 118755 4100
rect 118697 4091 118755 4097
rect 118970 4088 118976 4100
rect 119028 4128 119034 4140
rect 120350 4128 120356 4140
rect 119028 4100 120356 4128
rect 119028 4088 119034 4100
rect 120350 4088 120356 4100
rect 120408 4088 120414 4140
rect 120626 4088 120632 4140
rect 120684 4128 120690 4140
rect 120721 4131 120779 4137
rect 120721 4128 120733 4131
rect 120684 4100 120733 4128
rect 120684 4088 120690 4100
rect 120721 4097 120733 4100
rect 120767 4097 120779 4131
rect 120721 4091 120779 4097
rect 121917 4131 121975 4137
rect 121917 4097 121929 4131
rect 121963 4097 121975 4131
rect 121917 4091 121975 4097
rect 117409 4063 117467 4069
rect 117409 4029 117421 4063
rect 117455 4029 117467 4063
rect 117409 4023 117467 4029
rect 103486 3964 115888 3992
rect 117424 3992 117452 4023
rect 118142 4020 118148 4072
rect 118200 4020 118206 4072
rect 121638 4020 121644 4072
rect 121696 4020 121702 4072
rect 121932 4060 121960 4091
rect 124490 4088 124496 4140
rect 124548 4088 124554 4140
rect 125134 4088 125140 4140
rect 125192 4088 125198 4140
rect 208946 4128 208952 4140
rect 128326 4100 132494 4128
rect 122561 4063 122619 4069
rect 122561 4060 122573 4063
rect 121932 4032 122573 4060
rect 122561 4029 122573 4032
rect 122607 4060 122619 4063
rect 122650 4060 122656 4072
rect 122607 4032 122656 4060
rect 122607 4029 122619 4032
rect 122561 4023 122619 4029
rect 122650 4020 122656 4032
rect 122708 4020 122714 4072
rect 123478 4020 123484 4072
rect 123536 4060 123542 4072
rect 126514 4060 126520 4072
rect 123536 4032 126520 4060
rect 123536 4020 123542 4032
rect 126514 4020 126520 4032
rect 126572 4020 126578 4072
rect 119154 3992 119160 4004
rect 117424 3964 119160 3992
rect 56502 3884 56508 3936
rect 56560 3924 56566 3936
rect 103486 3924 103514 3964
rect 119154 3952 119160 3964
rect 119212 3952 119218 4004
rect 128326 3992 128354 4100
rect 119264 3964 128354 3992
rect 132466 3992 132494 4100
rect 200086 4100 208952 4128
rect 200086 3992 200114 4100
rect 208946 4088 208952 4100
rect 209004 4088 209010 4140
rect 209038 4088 209044 4140
rect 209096 4088 209102 4140
rect 210145 4131 210203 4137
rect 210145 4097 210157 4131
rect 210191 4097 210203 4131
rect 210145 4091 210203 4097
rect 200942 4020 200948 4072
rect 201000 4060 201006 4072
rect 209593 4063 209651 4069
rect 209593 4060 209605 4063
rect 201000 4032 209605 4060
rect 201000 4020 201006 4032
rect 209593 4029 209605 4032
rect 209639 4029 209651 4063
rect 209593 4023 209651 4029
rect 210160 3992 210188 4091
rect 211062 4088 211068 4140
rect 211120 4128 211126 4140
rect 211249 4131 211307 4137
rect 211249 4128 211261 4131
rect 211120 4100 211261 4128
rect 211120 4088 211126 4100
rect 211249 4097 211261 4100
rect 211295 4097 211307 4131
rect 211249 4091 211307 4097
rect 212810 4088 212816 4140
rect 212868 4088 212874 4140
rect 213362 4088 213368 4140
rect 213420 4088 213426 4140
rect 213914 4088 213920 4140
rect 213972 4088 213978 4140
rect 215478 4088 215484 4140
rect 215536 4088 215542 4140
rect 216950 4088 216956 4140
rect 217008 4137 217014 4140
rect 217008 4131 217057 4137
rect 217008 4097 217011 4131
rect 217045 4097 217057 4131
rect 217008 4091 217057 4097
rect 217008 4088 217014 4091
rect 217318 4088 217324 4140
rect 217376 4128 217382 4140
rect 217376 4100 306374 4128
rect 217376 4088 217382 4100
rect 214926 4020 214932 4072
rect 214984 4020 214990 4072
rect 216674 4020 216680 4072
rect 216732 4020 216738 4072
rect 217612 4032 218100 4060
rect 210418 3992 210424 4004
rect 132466 3964 200114 3992
rect 200776 3964 209774 3992
rect 210160 3964 210424 3992
rect 56560 3896 103514 3924
rect 56560 3884 56566 3896
rect 116670 3884 116676 3936
rect 116728 3924 116734 3936
rect 119264 3924 119292 3964
rect 116728 3896 119292 3924
rect 116728 3884 116734 3896
rect 119338 3884 119344 3936
rect 119396 3884 119402 3936
rect 120261 3927 120319 3933
rect 120261 3893 120273 3927
rect 120307 3924 120319 3927
rect 120810 3924 120816 3936
rect 120307 3896 120816 3924
rect 120307 3893 120319 3896
rect 120261 3887 120319 3893
rect 120810 3884 120816 3896
rect 120868 3924 120874 3936
rect 200776 3924 200804 3964
rect 120868 3896 200804 3924
rect 120868 3884 120874 3896
rect 208394 3884 208400 3936
rect 208452 3884 208458 3936
rect 208486 3884 208492 3936
rect 208544 3924 208550 3936
rect 209590 3924 209596 3936
rect 208544 3896 209596 3924
rect 208544 3884 208550 3896
rect 209590 3884 209596 3896
rect 209648 3884 209654 3936
rect 209746 3924 209774 3964
rect 210418 3952 210424 3964
rect 210476 3992 210482 4004
rect 217612 3992 217640 4032
rect 210476 3964 217640 3992
rect 218072 3992 218100 4032
rect 218146 4020 218152 4072
rect 218204 4060 218210 4072
rect 218204 4032 301544 4060
rect 218204 4020 218210 4032
rect 301516 3992 301544 4032
rect 304166 4020 304172 4072
rect 304224 4020 304230 4072
rect 304810 4020 304816 4072
rect 304868 4020 304874 4072
rect 305178 4020 305184 4072
rect 305236 4060 305242 4072
rect 306193 4063 306251 4069
rect 306193 4060 306205 4063
rect 305236 4032 306205 4060
rect 305236 4020 305242 4032
rect 306193 4029 306205 4032
rect 306239 4029 306251 4063
rect 306346 4060 306374 4100
rect 306466 4088 306472 4140
rect 306524 4088 306530 4140
rect 306558 4088 306564 4140
rect 306616 4128 306622 4140
rect 307481 4131 307539 4137
rect 307481 4128 307493 4131
rect 306616 4100 307493 4128
rect 306616 4088 306622 4100
rect 307481 4097 307493 4100
rect 307527 4097 307539 4131
rect 307481 4091 307539 4097
rect 307662 4088 307668 4140
rect 307720 4128 307726 4140
rect 309137 4131 309195 4137
rect 307720 4100 308996 4128
rect 307720 4088 307726 4100
rect 308674 4060 308680 4072
rect 306346 4032 308680 4060
rect 306193 4023 306251 4029
rect 308674 4020 308680 4032
rect 308732 4020 308738 4072
rect 308861 4063 308919 4069
rect 308861 4029 308873 4063
rect 308907 4029 308919 4063
rect 308861 4023 308919 4029
rect 308876 3992 308904 4023
rect 218072 3964 224954 3992
rect 210476 3952 210482 3964
rect 212534 3924 212540 3936
rect 209746 3896 212540 3924
rect 212534 3884 212540 3896
rect 212592 3884 212598 3936
rect 216950 3884 216956 3936
rect 217008 3924 217014 3936
rect 217781 3927 217839 3933
rect 217781 3924 217793 3927
rect 217008 3896 217793 3924
rect 217008 3884 217014 3896
rect 217781 3893 217793 3896
rect 217827 3924 217839 3927
rect 218054 3924 218060 3936
rect 217827 3896 218060 3924
rect 217827 3893 217839 3896
rect 217781 3887 217839 3893
rect 218054 3884 218060 3896
rect 218112 3884 218118 3936
rect 218514 3884 218520 3936
rect 218572 3884 218578 3936
rect 219526 3884 219532 3936
rect 219584 3884 219590 3936
rect 219618 3884 219624 3936
rect 219676 3924 219682 3936
rect 220446 3924 220452 3936
rect 219676 3896 220452 3924
rect 219676 3884 219682 3896
rect 220446 3884 220452 3896
rect 220504 3884 220510 3936
rect 224926 3924 224954 3964
rect 229066 3964 296714 3992
rect 301516 3964 308904 3992
rect 308968 3992 308996 4100
rect 309137 4097 309149 4131
rect 309183 4128 309195 4131
rect 309686 4128 309692 4140
rect 309183 4100 309692 4128
rect 309183 4097 309195 4100
rect 309137 4091 309195 4097
rect 309686 4088 309692 4100
rect 309744 4088 309750 4140
rect 310422 4088 310428 4140
rect 310480 4128 310486 4140
rect 310517 4131 310575 4137
rect 310517 4128 310529 4131
rect 310480 4100 310529 4128
rect 310480 4088 310486 4100
rect 310517 4097 310529 4100
rect 310563 4097 310575 4131
rect 310517 4091 310575 4097
rect 310606 4088 310612 4140
rect 310664 4128 310670 4140
rect 311434 4128 311440 4140
rect 310664 4100 311440 4128
rect 310664 4088 310670 4100
rect 311434 4088 311440 4100
rect 311492 4088 311498 4140
rect 309226 4020 309232 4072
rect 309284 4060 309290 4072
rect 340046 4060 340052 4072
rect 309284 4032 340052 4060
rect 309284 4020 309290 4032
rect 340046 4020 340052 4032
rect 340104 4020 340110 4072
rect 310606 3992 310612 4004
rect 308968 3964 310612 3992
rect 229066 3924 229094 3964
rect 224926 3896 229094 3924
rect 296686 3924 296714 3964
rect 310606 3952 310612 3964
rect 310664 3952 310670 4004
rect 310698 3952 310704 4004
rect 310756 3952 310762 4004
rect 316770 3992 316776 4004
rect 310808 3964 316776 3992
rect 303982 3924 303988 3936
rect 296686 3896 303988 3924
rect 303982 3884 303988 3896
rect 304040 3884 304046 3936
rect 305454 3884 305460 3936
rect 305512 3884 305518 3936
rect 306466 3884 306472 3936
rect 306524 3924 306530 3936
rect 307018 3924 307024 3936
rect 306524 3896 307024 3924
rect 306524 3884 306530 3896
rect 307018 3884 307024 3896
rect 307076 3884 307082 3936
rect 307662 3884 307668 3936
rect 307720 3884 307726 3936
rect 309686 3884 309692 3936
rect 309744 3884 309750 3936
rect 309778 3884 309784 3936
rect 309836 3924 309842 3936
rect 310808 3924 310836 3964
rect 316770 3952 316776 3964
rect 316828 3952 316834 4004
rect 401502 3992 401508 4004
rect 321526 3964 401508 3992
rect 309836 3896 310836 3924
rect 309836 3884 309842 3896
rect 311342 3884 311348 3936
rect 311400 3884 311406 3936
rect 311434 3884 311440 3936
rect 311492 3924 311498 3936
rect 321526 3924 321554 3964
rect 401502 3952 401508 3964
rect 401560 3952 401566 4004
rect 311492 3896 321554 3924
rect 311492 3884 311498 3896
rect 1104 3834 528816 3856
rect 1104 3782 66914 3834
rect 66966 3782 66978 3834
rect 67030 3782 67042 3834
rect 67094 3782 67106 3834
rect 67158 3782 67170 3834
rect 67222 3782 198842 3834
rect 198894 3782 198906 3834
rect 198958 3782 198970 3834
rect 199022 3782 199034 3834
rect 199086 3782 199098 3834
rect 199150 3782 330770 3834
rect 330822 3782 330834 3834
rect 330886 3782 330898 3834
rect 330950 3782 330962 3834
rect 331014 3782 331026 3834
rect 331078 3782 462698 3834
rect 462750 3782 462762 3834
rect 462814 3782 462826 3834
rect 462878 3782 462890 3834
rect 462942 3782 462954 3834
rect 463006 3782 528816 3834
rect 1104 3760 528816 3782
rect 113821 3723 113879 3729
rect 113821 3689 113833 3723
rect 113867 3720 113879 3723
rect 114094 3720 114100 3732
rect 113867 3692 114100 3720
rect 113867 3689 113879 3692
rect 113821 3683 113879 3689
rect 114094 3680 114100 3692
rect 114152 3720 114158 3732
rect 117406 3720 117412 3732
rect 114152 3692 117412 3720
rect 114152 3680 114158 3692
rect 117406 3680 117412 3692
rect 117464 3680 117470 3732
rect 125870 3680 125876 3732
rect 125928 3680 125934 3732
rect 126422 3680 126428 3732
rect 126480 3680 126486 3732
rect 126514 3680 126520 3732
rect 126572 3720 126578 3732
rect 216582 3720 216588 3732
rect 126572 3692 216588 3720
rect 126572 3680 126578 3692
rect 216582 3680 216588 3692
rect 216640 3680 216646 3732
rect 220446 3680 220452 3732
rect 220504 3680 220510 3732
rect 220538 3680 220544 3732
rect 220596 3720 220602 3732
rect 310698 3720 310704 3732
rect 220596 3692 310704 3720
rect 220596 3680 220602 3692
rect 310698 3680 310704 3692
rect 310756 3680 310762 3732
rect 312722 3680 312728 3732
rect 312780 3720 312786 3732
rect 313185 3723 313243 3729
rect 313185 3720 313197 3723
rect 312780 3692 313197 3720
rect 312780 3680 312786 3692
rect 313185 3689 313197 3692
rect 313231 3720 313243 3723
rect 350534 3720 350540 3732
rect 313231 3692 350540 3720
rect 313231 3689 313243 3692
rect 313185 3683 313243 3689
rect 350534 3680 350540 3692
rect 350592 3680 350598 3732
rect 353938 3680 353944 3732
rect 353996 3720 354002 3732
rect 410242 3720 410248 3732
rect 353996 3692 410248 3720
rect 353996 3680 354002 3692
rect 410242 3680 410248 3692
rect 410300 3680 410306 3732
rect 116026 3612 116032 3664
rect 116084 3652 116090 3664
rect 200942 3652 200948 3664
rect 116084 3624 200948 3652
rect 116084 3612 116090 3624
rect 200942 3612 200948 3624
rect 201000 3612 201006 3664
rect 204272 3624 211660 3652
rect 108298 3544 108304 3596
rect 108356 3584 108362 3596
rect 114922 3584 114928 3596
rect 108356 3556 114928 3584
rect 108356 3544 108362 3556
rect 114922 3544 114928 3556
rect 114980 3544 114986 3596
rect 117314 3584 117320 3596
rect 115492 3556 117320 3584
rect 115492 3525 115520 3556
rect 117314 3544 117320 3556
rect 117372 3544 117378 3596
rect 118418 3584 118424 3596
rect 118160 3556 118424 3584
rect 114373 3519 114431 3525
rect 114373 3485 114385 3519
rect 114419 3516 114431 3519
rect 115477 3519 115535 3525
rect 115477 3516 115489 3519
rect 114419 3488 115489 3516
rect 114419 3485 114431 3488
rect 114373 3479 114431 3485
rect 115477 3485 115489 3488
rect 115523 3485 115535 3519
rect 115477 3479 115535 3485
rect 116670 3476 116676 3528
rect 116728 3476 116734 3528
rect 118160 3525 118188 3556
rect 118418 3544 118424 3556
rect 118476 3584 118482 3596
rect 204272 3584 204300 3624
rect 211632 3593 211660 3624
rect 211706 3612 211712 3664
rect 211764 3652 211770 3664
rect 219710 3652 219716 3664
rect 211764 3624 219716 3652
rect 211764 3612 211770 3624
rect 219710 3612 219716 3624
rect 219768 3612 219774 3664
rect 219820 3624 220308 3652
rect 211617 3587 211675 3593
rect 118476 3556 204300 3584
rect 204916 3556 211568 3584
rect 118476 3544 118482 3556
rect 118145 3519 118203 3525
rect 118145 3485 118157 3519
rect 118191 3485 118203 3519
rect 118145 3479 118203 3485
rect 118786 3476 118792 3528
rect 118844 3476 118850 3528
rect 119338 3476 119344 3528
rect 119396 3476 119402 3528
rect 120074 3476 120080 3528
rect 120132 3476 120138 3528
rect 120534 3476 120540 3528
rect 120592 3516 120598 3528
rect 120718 3516 120724 3528
rect 120592 3488 120724 3516
rect 120592 3476 120598 3488
rect 120718 3476 120724 3488
rect 120776 3476 120782 3528
rect 121273 3519 121331 3525
rect 121273 3485 121285 3519
rect 121319 3485 121331 3519
rect 121273 3479 121331 3485
rect 124309 3519 124367 3525
rect 124309 3485 124321 3519
rect 124355 3516 124367 3519
rect 125134 3516 125140 3528
rect 124355 3488 125140 3516
rect 124355 3485 124367 3488
rect 124309 3479 124367 3485
rect 22186 3408 22192 3460
rect 22244 3448 22250 3460
rect 114925 3451 114983 3457
rect 114925 3448 114937 3451
rect 22244 3420 114937 3448
rect 22244 3408 22250 3420
rect 114925 3417 114937 3420
rect 114971 3417 114983 3451
rect 114925 3411 114983 3417
rect 116118 3408 116124 3460
rect 116176 3408 116182 3460
rect 117590 3408 117596 3460
rect 117648 3408 117654 3460
rect 119154 3408 119160 3460
rect 119212 3448 119218 3460
rect 119982 3448 119988 3460
rect 119212 3420 119988 3448
rect 119212 3408 119218 3420
rect 119982 3408 119988 3420
rect 120040 3408 120046 3460
rect 120626 3408 120632 3460
rect 120684 3448 120690 3460
rect 121288 3448 121316 3479
rect 125134 3476 125140 3488
rect 125192 3476 125198 3528
rect 125321 3519 125379 3525
rect 125321 3485 125333 3519
rect 125367 3516 125379 3519
rect 125870 3516 125876 3528
rect 125367 3488 125876 3516
rect 125367 3485 125379 3488
rect 125321 3479 125379 3485
rect 125870 3476 125876 3488
rect 125928 3476 125934 3528
rect 204916 3516 204944 3556
rect 200086 3488 204944 3516
rect 208305 3519 208363 3525
rect 120684 3420 121316 3448
rect 120684 3408 120690 3420
rect 121822 3408 121828 3460
rect 121880 3408 121886 3460
rect 122374 3408 122380 3460
rect 122432 3448 122438 3460
rect 122432 3420 123340 3448
rect 122432 3408 122438 3420
rect 122558 3340 122564 3392
rect 122616 3340 122622 3392
rect 123202 3340 123208 3392
rect 123260 3340 123266 3392
rect 123312 3380 123340 3420
rect 123754 3408 123760 3460
rect 123812 3408 123818 3460
rect 125042 3408 125048 3460
rect 125100 3408 125106 3460
rect 125226 3408 125232 3460
rect 125284 3448 125290 3460
rect 126882 3448 126888 3460
rect 125284 3420 126888 3448
rect 125284 3408 125290 3420
rect 126882 3408 126888 3420
rect 126940 3408 126946 3460
rect 200086 3448 200114 3488
rect 208305 3485 208317 3519
rect 208351 3516 208363 3519
rect 208486 3516 208492 3528
rect 208351 3488 208492 3516
rect 208351 3485 208363 3488
rect 208305 3479 208363 3485
rect 208486 3476 208492 3488
rect 208544 3476 208550 3528
rect 208854 3476 208860 3528
rect 208912 3476 208918 3528
rect 209038 3476 209044 3528
rect 209096 3516 209102 3528
rect 209409 3519 209467 3525
rect 209409 3516 209421 3519
rect 209096 3488 209421 3516
rect 209096 3476 209102 3488
rect 209409 3485 209421 3488
rect 209455 3485 209467 3519
rect 209409 3479 209467 3485
rect 210973 3519 211031 3525
rect 210973 3485 210985 3519
rect 211019 3485 211031 3519
rect 211540 3516 211568 3556
rect 211617 3553 211629 3587
rect 211663 3553 211675 3587
rect 216493 3587 216551 3593
rect 216493 3584 216505 3587
rect 211617 3547 211675 3553
rect 212000 3556 216505 3584
rect 212000 3516 212028 3556
rect 216493 3553 216505 3556
rect 216539 3553 216551 3587
rect 219820 3584 219848 3624
rect 216493 3547 216551 3553
rect 216968 3556 219848 3584
rect 220280 3584 220308 3624
rect 220630 3612 220636 3664
rect 220688 3652 220694 3664
rect 308490 3652 308496 3664
rect 220688 3624 308496 3652
rect 220688 3612 220694 3624
rect 308490 3612 308496 3624
rect 308548 3612 308554 3664
rect 308674 3612 308680 3664
rect 308732 3652 308738 3664
rect 308732 3624 309180 3652
rect 308732 3612 308738 3624
rect 309045 3587 309103 3593
rect 309045 3584 309057 3587
rect 220280 3556 309057 3584
rect 211540 3488 212028 3516
rect 210973 3479 211031 3485
rect 128326 3420 200114 3448
rect 200592 3420 208348 3448
rect 128326 3380 128354 3420
rect 123312 3352 128354 3380
rect 164326 3340 164332 3392
rect 164384 3380 164390 3392
rect 200592 3380 200620 3420
rect 164384 3352 200620 3380
rect 208320 3380 208348 3420
rect 208946 3408 208952 3460
rect 209004 3448 209010 3460
rect 210421 3451 210479 3457
rect 210421 3448 210433 3451
rect 209004 3420 210433 3448
rect 209004 3408 209010 3420
rect 210421 3417 210433 3420
rect 210467 3417 210479 3451
rect 210988 3448 211016 3479
rect 212166 3476 212172 3528
rect 212224 3476 212230 3528
rect 212902 3476 212908 3528
rect 212960 3516 212966 3528
rect 213365 3519 213423 3525
rect 213365 3516 213377 3519
rect 212960 3488 213377 3516
rect 212960 3476 212966 3488
rect 213365 3485 213377 3488
rect 213411 3485 213423 3519
rect 213365 3479 213423 3485
rect 214561 3519 214619 3525
rect 214561 3485 214573 3519
rect 214607 3485 214619 3519
rect 214561 3479 214619 3485
rect 211706 3448 211712 3460
rect 210988 3420 211712 3448
rect 210421 3411 210479 3417
rect 211706 3408 211712 3420
rect 211764 3408 211770 3460
rect 212626 3408 212632 3460
rect 212684 3448 212690 3460
rect 212813 3451 212871 3457
rect 212813 3448 212825 3451
rect 212684 3420 212825 3448
rect 212684 3408 212690 3420
rect 212813 3417 212825 3420
rect 212859 3417 212871 3451
rect 212813 3411 212871 3417
rect 214006 3408 214012 3460
rect 214064 3408 214070 3460
rect 214576 3448 214604 3479
rect 215202 3476 215208 3528
rect 215260 3516 215266 3528
rect 215297 3519 215355 3525
rect 215297 3516 215309 3519
rect 215260 3488 215309 3516
rect 215260 3476 215266 3488
rect 215297 3485 215309 3488
rect 215343 3485 215355 3519
rect 216968 3516 216996 3556
rect 309045 3553 309057 3556
rect 309091 3553 309103 3587
rect 309152 3584 309180 3624
rect 309686 3612 309692 3664
rect 309744 3652 309750 3664
rect 319990 3652 319996 3664
rect 309744 3624 319996 3652
rect 309744 3612 309750 3624
rect 319990 3612 319996 3624
rect 320048 3612 320054 3664
rect 351914 3612 351920 3664
rect 351972 3652 351978 3664
rect 354030 3652 354036 3664
rect 351972 3624 354036 3652
rect 351972 3612 351978 3624
rect 354030 3612 354036 3624
rect 354088 3612 354094 3664
rect 355870 3612 355876 3664
rect 355928 3652 355934 3664
rect 401226 3652 401232 3664
rect 355928 3624 401232 3652
rect 355928 3612 355934 3624
rect 401226 3612 401232 3624
rect 401284 3612 401290 3664
rect 309965 3587 310023 3593
rect 309965 3584 309977 3587
rect 309152 3556 309977 3584
rect 309045 3547 309103 3553
rect 309965 3553 309977 3556
rect 310011 3553 310023 3587
rect 324498 3584 324504 3596
rect 309965 3547 310023 3553
rect 310256 3556 324504 3584
rect 215297 3479 215355 3485
rect 215404 3488 216996 3516
rect 217045 3519 217103 3525
rect 214834 3448 214840 3460
rect 214576 3420 214840 3448
rect 214834 3408 214840 3420
rect 214892 3448 214898 3460
rect 215404 3448 215432 3488
rect 217045 3485 217057 3519
rect 217091 3485 217103 3519
rect 217045 3479 217103 3485
rect 214892 3420 215432 3448
rect 214892 3408 214898 3420
rect 215846 3408 215852 3460
rect 215904 3408 215910 3460
rect 217060 3448 217088 3479
rect 217134 3476 217140 3528
rect 217192 3516 217198 3528
rect 217689 3519 217747 3525
rect 217689 3516 217701 3519
rect 217192 3488 217701 3516
rect 217192 3476 217198 3488
rect 217689 3485 217701 3488
rect 217735 3485 217747 3519
rect 217689 3479 217747 3485
rect 218241 3519 218299 3525
rect 218241 3485 218253 3519
rect 218287 3516 218299 3519
rect 218514 3516 218520 3528
rect 218287 3488 218520 3516
rect 218287 3485 218299 3488
rect 218241 3479 218299 3485
rect 218514 3476 218520 3488
rect 218572 3476 218578 3528
rect 218882 3476 218888 3528
rect 218940 3476 218946 3528
rect 219437 3519 219495 3525
rect 219437 3485 219449 3519
rect 219483 3516 219495 3519
rect 219618 3516 219624 3528
rect 219483 3488 219624 3516
rect 219483 3485 219495 3488
rect 219437 3479 219495 3485
rect 219618 3476 219624 3488
rect 219676 3476 219682 3528
rect 219710 3476 219716 3528
rect 219768 3516 219774 3528
rect 219768 3488 302924 3516
rect 219768 3476 219774 3488
rect 217226 3448 217232 3460
rect 217060 3420 217232 3448
rect 217226 3408 217232 3420
rect 217284 3448 217290 3460
rect 219986 3448 219992 3460
rect 217284 3420 219992 3448
rect 217284 3408 217290 3420
rect 219986 3408 219992 3420
rect 220044 3408 220050 3460
rect 220096 3420 229094 3448
rect 220096 3380 220124 3420
rect 208320 3352 220124 3380
rect 164384 3340 164390 3352
rect 220170 3340 220176 3392
rect 220228 3380 220234 3392
rect 220630 3380 220636 3392
rect 220228 3352 220636 3380
rect 220228 3340 220234 3352
rect 220630 3340 220636 3352
rect 220688 3340 220694 3392
rect 229066 3380 229094 3420
rect 300854 3408 300860 3460
rect 300912 3408 300918 3460
rect 259086 3380 259092 3392
rect 229066 3352 259092 3380
rect 259086 3340 259092 3352
rect 259144 3340 259150 3392
rect 300121 3383 300179 3389
rect 300121 3349 300133 3383
rect 300167 3380 300179 3383
rect 300302 3380 300308 3392
rect 300167 3352 300308 3380
rect 300167 3349 300179 3352
rect 300121 3343 300179 3349
rect 300302 3340 300308 3352
rect 300360 3340 300366 3392
rect 302786 3340 302792 3392
rect 302844 3340 302850 3392
rect 302896 3380 302924 3488
rect 303430 3476 303436 3528
rect 303488 3476 303494 3528
rect 303982 3476 303988 3528
rect 304040 3476 304046 3528
rect 304537 3519 304595 3525
rect 304537 3485 304549 3519
rect 304583 3516 304595 3519
rect 304810 3516 304816 3528
rect 304583 3488 304816 3516
rect 304583 3485 304595 3488
rect 304537 3479 304595 3485
rect 304810 3476 304816 3488
rect 304868 3476 304874 3528
rect 305270 3476 305276 3528
rect 305328 3476 305334 3528
rect 305546 3476 305552 3528
rect 305604 3476 305610 3528
rect 306098 3476 306104 3528
rect 306156 3516 306162 3528
rect 306193 3519 306251 3525
rect 306193 3516 306205 3519
rect 306156 3488 306205 3516
rect 306156 3476 306162 3488
rect 306193 3485 306205 3488
rect 306239 3485 306251 3519
rect 306193 3479 306251 3485
rect 306466 3476 306472 3528
rect 306524 3476 306530 3528
rect 307389 3519 307447 3525
rect 307389 3485 307401 3519
rect 307435 3485 307447 3519
rect 307389 3479 307447 3485
rect 307110 3408 307116 3460
rect 307168 3408 307174 3460
rect 307404 3448 307432 3479
rect 308122 3476 308128 3528
rect 308180 3476 308186 3528
rect 308401 3519 308459 3525
rect 308401 3485 308413 3519
rect 308447 3516 308459 3519
rect 309226 3516 309232 3528
rect 308447 3488 309232 3516
rect 308447 3485 308459 3488
rect 308401 3479 308459 3485
rect 309226 3476 309232 3488
rect 309284 3476 309290 3528
rect 309321 3519 309379 3525
rect 309321 3485 309333 3519
rect 309367 3516 309379 3519
rect 309594 3516 309600 3528
rect 309367 3488 309600 3516
rect 309367 3485 309379 3488
rect 309321 3479 309379 3485
rect 309594 3476 309600 3488
rect 309652 3516 309658 3528
rect 310256 3525 310284 3556
rect 324498 3544 324504 3556
rect 324556 3544 324562 3596
rect 331306 3584 331312 3596
rect 325666 3556 331312 3584
rect 310241 3519 310299 3525
rect 309652 3488 310192 3516
rect 309652 3476 309658 3488
rect 307570 3448 307576 3460
rect 307404 3420 307576 3448
rect 307570 3408 307576 3420
rect 307628 3448 307634 3460
rect 309778 3448 309784 3460
rect 307628 3420 309784 3448
rect 307628 3408 307634 3420
rect 309778 3408 309784 3420
rect 309836 3408 309842 3460
rect 310164 3448 310192 3488
rect 310241 3485 310253 3519
rect 310287 3485 310299 3519
rect 310241 3479 310299 3485
rect 310882 3476 310888 3528
rect 310940 3476 310946 3528
rect 311158 3476 311164 3528
rect 311216 3476 311222 3528
rect 325666 3516 325694 3556
rect 331306 3544 331312 3556
rect 331364 3544 331370 3596
rect 336366 3544 336372 3596
rect 336424 3584 336430 3596
rect 406470 3584 406476 3596
rect 336424 3556 406476 3584
rect 336424 3544 336430 3556
rect 406470 3544 406476 3556
rect 406528 3544 406534 3596
rect 311268 3488 325694 3516
rect 311268 3448 311296 3488
rect 348234 3476 348240 3528
rect 348292 3516 348298 3528
rect 399386 3516 399392 3528
rect 348292 3488 399392 3516
rect 348292 3476 348298 3488
rect 399386 3476 399392 3488
rect 399444 3476 399450 3528
rect 310164 3420 311296 3448
rect 311713 3451 311771 3457
rect 311713 3417 311725 3451
rect 311759 3448 311771 3451
rect 311759 3420 316724 3448
rect 311759 3417 311771 3420
rect 311713 3411 311771 3417
rect 307386 3380 307392 3392
rect 302896 3352 307392 3380
rect 307386 3340 307392 3352
rect 307444 3340 307450 3392
rect 309410 3340 309416 3392
rect 309468 3380 309474 3392
rect 311728 3380 311756 3411
rect 309468 3352 311756 3380
rect 309468 3340 309474 3352
rect 312262 3340 312268 3392
rect 312320 3340 312326 3392
rect 316696 3380 316724 3420
rect 316770 3408 316776 3460
rect 316828 3448 316834 3460
rect 344278 3448 344284 3460
rect 316828 3420 344284 3448
rect 316828 3408 316834 3420
rect 344278 3408 344284 3420
rect 344336 3408 344342 3460
rect 356974 3448 356980 3460
rect 344986 3420 356980 3448
rect 344986 3380 345014 3420
rect 356974 3408 356980 3420
rect 357032 3408 357038 3460
rect 409414 3448 409420 3460
rect 357084 3420 409420 3448
rect 316696 3352 345014 3380
rect 350442 3340 350448 3392
rect 350500 3380 350506 3392
rect 357084 3380 357112 3420
rect 409414 3408 409420 3420
rect 409472 3408 409478 3460
rect 350500 3352 357112 3380
rect 350500 3340 350506 3352
rect 357158 3340 357164 3392
rect 357216 3340 357222 3392
rect 393590 3340 393596 3392
rect 393648 3340 393654 3392
rect 394234 3340 394240 3392
rect 394292 3340 394298 3392
rect 394694 3340 394700 3392
rect 394752 3340 394758 3392
rect 396721 3383 396779 3389
rect 396721 3349 396733 3383
rect 396767 3380 396779 3383
rect 396902 3380 396908 3392
rect 396767 3352 396908 3380
rect 396767 3349 396779 3352
rect 396721 3343 396779 3349
rect 396902 3340 396908 3352
rect 396960 3340 396966 3392
rect 397362 3340 397368 3392
rect 397420 3380 397426 3392
rect 491294 3380 491300 3392
rect 397420 3352 491300 3380
rect 397420 3340 397426 3352
rect 491294 3340 491300 3352
rect 491352 3340 491358 3392
rect 1104 3290 528816 3312
rect 1104 3238 67574 3290
rect 67626 3238 67638 3290
rect 67690 3238 67702 3290
rect 67754 3238 67766 3290
rect 67818 3238 67830 3290
rect 67882 3238 199502 3290
rect 199554 3238 199566 3290
rect 199618 3238 199630 3290
rect 199682 3238 199694 3290
rect 199746 3238 199758 3290
rect 199810 3238 331430 3290
rect 331482 3238 331494 3290
rect 331546 3238 331558 3290
rect 331610 3238 331622 3290
rect 331674 3238 331686 3290
rect 331738 3238 463358 3290
rect 463410 3238 463422 3290
rect 463474 3238 463486 3290
rect 463538 3238 463550 3290
rect 463602 3238 463614 3290
rect 463666 3238 528816 3290
rect 1104 3216 528816 3238
rect 27614 3136 27620 3188
rect 27672 3176 27678 3188
rect 116118 3176 116124 3188
rect 27672 3148 116124 3176
rect 27672 3136 27678 3148
rect 116118 3136 116124 3148
rect 116176 3136 116182 3188
rect 117498 3176 117504 3188
rect 116872 3148 117504 3176
rect 22094 3068 22100 3120
rect 22152 3108 22158 3120
rect 115109 3111 115167 3117
rect 115109 3108 115121 3111
rect 22152 3080 113174 3108
rect 22152 3068 22158 3080
rect 108298 3040 108304 3052
rect 37476 3012 108304 3040
rect 24854 2932 24860 2984
rect 24912 2972 24918 2984
rect 37366 2972 37372 2984
rect 24912 2944 37372 2972
rect 24912 2932 24918 2944
rect 37366 2932 37372 2944
rect 37424 2932 37430 2984
rect 31754 2864 31760 2916
rect 31812 2904 31818 2916
rect 37476 2904 37504 3012
rect 108298 3000 108304 3012
rect 108356 3000 108362 3052
rect 113146 3040 113174 3080
rect 113468 3080 115121 3108
rect 113358 3040 113364 3052
rect 113146 3012 113364 3040
rect 113358 3000 113364 3012
rect 113416 3000 113422 3052
rect 37550 2932 37556 2984
rect 37608 2972 37614 2984
rect 113468 2972 113496 3080
rect 115109 3077 115121 3080
rect 115155 3077 115167 3111
rect 115109 3071 115167 3077
rect 116302 3068 116308 3120
rect 116360 3068 116366 3120
rect 114094 3000 114100 3052
rect 114152 3000 114158 3052
rect 115658 3000 115664 3052
rect 115716 3000 115722 3052
rect 116872 3049 116900 3148
rect 117498 3136 117504 3148
rect 117556 3176 117562 3188
rect 210234 3176 210240 3188
rect 117556 3148 210240 3176
rect 117556 3136 117562 3148
rect 210234 3136 210240 3148
rect 210292 3136 210298 3188
rect 215386 3176 215392 3188
rect 210344 3148 214236 3176
rect 118694 3068 118700 3120
rect 118752 3068 118758 3120
rect 120258 3068 120264 3120
rect 120316 3068 120322 3120
rect 120736 3080 123064 3108
rect 116857 3043 116915 3049
rect 116857 3009 116869 3043
rect 116903 3009 116915 3043
rect 116857 3003 116915 3009
rect 117866 3000 117872 3052
rect 117924 3040 117930 3052
rect 118053 3043 118111 3049
rect 118053 3040 118065 3043
rect 117924 3012 118065 3040
rect 117924 3000 117930 3012
rect 118053 3009 118065 3012
rect 118099 3040 118111 3043
rect 119249 3043 119307 3049
rect 118099 3012 118694 3040
rect 118099 3009 118111 3012
rect 118053 3003 118111 3009
rect 37608 2944 113496 2972
rect 113545 2975 113603 2981
rect 37608 2932 37614 2944
rect 113545 2941 113557 2975
rect 113591 2941 113603 2975
rect 113545 2935 113603 2941
rect 113560 2904 113588 2935
rect 117314 2932 117320 2984
rect 117372 2972 117378 2984
rect 117501 2975 117559 2981
rect 117501 2972 117513 2975
rect 117372 2944 117513 2972
rect 117372 2932 117378 2944
rect 117501 2941 117513 2944
rect 117547 2941 117559 2975
rect 117501 2935 117559 2941
rect 31812 2876 37504 2904
rect 37568 2876 113588 2904
rect 118666 2904 118694 3012
rect 119249 3009 119261 3043
rect 119295 3040 119307 3043
rect 119522 3040 119528 3052
rect 119295 3012 119528 3040
rect 119295 3009 119307 3012
rect 119249 3003 119307 3009
rect 119522 3000 119528 3012
rect 119580 3040 119586 3052
rect 120736 3040 120764 3080
rect 119580 3012 120764 3040
rect 120813 3043 120871 3049
rect 119580 3000 119586 3012
rect 120813 3009 120825 3043
rect 120859 3040 120871 3043
rect 121362 3040 121368 3052
rect 120859 3012 121368 3040
rect 120859 3009 120871 3012
rect 120813 3003 120871 3009
rect 121362 3000 121368 3012
rect 121420 3040 121426 3052
rect 122009 3043 122067 3049
rect 121420 3012 121960 3040
rect 121420 3000 121426 3012
rect 121546 2932 121552 2984
rect 121604 2932 121610 2984
rect 121730 2904 121736 2916
rect 118666 2876 121736 2904
rect 31812 2864 31818 2876
rect 28994 2796 29000 2848
rect 29052 2836 29058 2848
rect 37568 2836 37596 2876
rect 121730 2864 121736 2876
rect 121788 2864 121794 2916
rect 121932 2904 121960 3012
rect 122009 3009 122021 3043
rect 122055 3040 122067 3043
rect 122558 3040 122564 3052
rect 122055 3012 122564 3040
rect 122055 3009 122067 3012
rect 122009 3003 122067 3009
rect 122558 3000 122564 3012
rect 122616 3000 122622 3052
rect 122926 2932 122932 2984
rect 122984 2932 122990 2984
rect 123036 2972 123064 3080
rect 123846 3068 123852 3120
rect 123904 3068 123910 3120
rect 127253 3111 127311 3117
rect 127253 3108 127265 3111
rect 124416 3080 127265 3108
rect 123202 3000 123208 3052
rect 123260 3000 123266 3052
rect 124416 3049 124444 3080
rect 127253 3077 127265 3080
rect 127299 3108 127311 3111
rect 127342 3108 127348 3120
rect 127299 3080 127348 3108
rect 127299 3077 127311 3080
rect 127253 3071 127311 3077
rect 127342 3068 127348 3080
rect 127400 3068 127406 3120
rect 127434 3068 127440 3120
rect 127492 3108 127498 3120
rect 210344 3108 210372 3148
rect 214208 3117 214236 3148
rect 215266 3148 215392 3176
rect 212997 3111 213055 3117
rect 212997 3108 213009 3111
rect 127492 3080 210372 3108
rect 210712 3080 213009 3108
rect 127492 3068 127498 3080
rect 124401 3043 124459 3049
rect 124401 3009 124413 3043
rect 124447 3009 124459 3043
rect 124401 3003 124459 3009
rect 124582 3000 124588 3052
rect 124640 3040 124646 3052
rect 124640 3012 125364 3040
rect 124640 3000 124646 3012
rect 125226 2972 125232 2984
rect 123036 2944 125232 2972
rect 125226 2932 125232 2944
rect 125284 2932 125290 2984
rect 125336 2972 125364 3012
rect 125410 3000 125416 3052
rect 125468 3000 125474 3052
rect 125689 3043 125747 3049
rect 125689 3009 125701 3043
rect 125735 3040 125747 3043
rect 126238 3040 126244 3052
rect 125735 3012 126244 3040
rect 125735 3009 125747 3012
rect 125689 3003 125747 3009
rect 126238 3000 126244 3012
rect 126296 3000 126302 3052
rect 126348 3012 128354 3040
rect 126348 2972 126376 3012
rect 125336 2944 126376 2972
rect 128326 2972 128354 3012
rect 145834 3000 145840 3052
rect 145892 3000 145898 3052
rect 164326 3000 164332 3052
rect 164384 3000 164390 3052
rect 168006 3000 168012 3052
rect 168064 3040 168070 3052
rect 168653 3043 168711 3049
rect 168653 3040 168665 3043
rect 168064 3012 168665 3040
rect 168064 3000 168070 3012
rect 168653 3009 168665 3012
rect 168699 3009 168711 3043
rect 168653 3003 168711 3009
rect 168760 3012 171134 3040
rect 168760 2972 168788 3012
rect 128326 2944 168788 2972
rect 169202 2932 169208 2984
rect 169260 2932 169266 2984
rect 171106 2972 171134 3012
rect 201678 3000 201684 3052
rect 201736 3040 201742 3052
rect 202417 3043 202475 3049
rect 202417 3040 202429 3043
rect 201736 3012 202429 3040
rect 201736 3000 201742 3012
rect 202417 3009 202429 3012
rect 202463 3009 202475 3043
rect 202417 3003 202475 3009
rect 202782 3000 202788 3052
rect 202840 3000 202846 3052
rect 205453 3043 205511 3049
rect 204824 3012 205036 3040
rect 204824 2972 204852 3012
rect 171106 2944 204852 2972
rect 204898 2932 204904 2984
rect 204956 2932 204962 2984
rect 205008 2972 205036 3012
rect 205453 3009 205465 3043
rect 205499 3040 205511 3043
rect 206186 3040 206192 3052
rect 205499 3012 206192 3040
rect 205499 3009 205511 3012
rect 205453 3003 205511 3009
rect 206186 3000 206192 3012
rect 206244 3000 206250 3052
rect 206830 3000 206836 3052
rect 206888 3040 206894 3052
rect 207569 3043 207627 3049
rect 207569 3040 207581 3043
rect 206888 3012 207581 3040
rect 206888 3000 206894 3012
rect 207569 3009 207581 3012
rect 207615 3009 207627 3043
rect 207569 3003 207627 3009
rect 207676 3012 209176 3040
rect 207676 2972 207704 3012
rect 205008 2944 207704 2972
rect 208118 2932 208124 2984
rect 208176 2932 208182 2984
rect 208578 2932 208584 2984
rect 208636 2972 208642 2984
rect 209041 2975 209099 2981
rect 209041 2972 209053 2975
rect 208636 2944 209053 2972
rect 208636 2932 208642 2944
rect 209041 2941 209053 2944
rect 209087 2941 209099 2975
rect 209148 2972 209176 3012
rect 209590 3000 209596 3052
rect 209648 3000 209654 3052
rect 210712 3040 210740 3080
rect 212997 3077 213009 3080
rect 213043 3077 213055 3111
rect 212997 3071 213055 3077
rect 214193 3111 214251 3117
rect 214193 3077 214205 3111
rect 214239 3077 214251 3111
rect 214193 3071 214251 3077
rect 209746 3012 210740 3040
rect 209746 2972 209774 3012
rect 210786 3000 210792 3052
rect 210844 3000 210850 3052
rect 211985 3043 212043 3049
rect 211985 3009 211997 3043
rect 212031 3040 212043 3043
rect 213178 3040 213184 3052
rect 212031 3012 213184 3040
rect 212031 3009 212043 3012
rect 211985 3003 212043 3009
rect 213178 3000 213184 3012
rect 213236 3000 213242 3052
rect 213546 3000 213552 3052
rect 213604 3000 213610 3052
rect 214745 3043 214803 3049
rect 214745 3009 214757 3043
rect 214791 3040 214803 3043
rect 215266 3040 215294 3148
rect 215386 3136 215392 3148
rect 215444 3176 215450 3188
rect 220538 3176 220544 3188
rect 215444 3148 220544 3176
rect 215444 3136 215450 3148
rect 220538 3136 220544 3148
rect 220596 3136 220602 3188
rect 221090 3136 221096 3188
rect 221148 3136 221154 3188
rect 221182 3136 221188 3188
rect 221240 3176 221246 3188
rect 309137 3179 309195 3185
rect 309137 3176 309149 3179
rect 221240 3148 309149 3176
rect 221240 3136 221246 3148
rect 309137 3145 309149 3148
rect 309183 3145 309195 3179
rect 309137 3139 309195 3145
rect 311158 3136 311164 3188
rect 311216 3176 311222 3188
rect 314654 3176 314660 3188
rect 311216 3148 314660 3176
rect 311216 3136 311222 3148
rect 314654 3136 314660 3148
rect 314712 3136 314718 3188
rect 314746 3136 314752 3188
rect 314804 3136 314810 3188
rect 317874 3136 317880 3188
rect 317932 3136 317938 3188
rect 331306 3136 331312 3188
rect 331364 3136 331370 3188
rect 340046 3136 340052 3188
rect 340104 3136 340110 3188
rect 344278 3136 344284 3188
rect 344336 3136 344342 3188
rect 345017 3179 345075 3185
rect 345017 3176 345029 3179
rect 344388 3148 345029 3176
rect 216582 3068 216588 3120
rect 216640 3068 216646 3120
rect 217060 3080 218836 3108
rect 214791 3012 215294 3040
rect 215941 3043 215999 3049
rect 214791 3009 214803 3012
rect 214745 3003 214803 3009
rect 215941 3009 215953 3043
rect 215987 3040 215999 3043
rect 216214 3040 216220 3052
rect 215987 3012 216220 3040
rect 215987 3009 215999 3012
rect 215941 3003 215999 3009
rect 216214 3000 216220 3012
rect 216272 3040 216278 3052
rect 217060 3040 217088 3080
rect 216272 3012 217088 3040
rect 217137 3043 217195 3049
rect 216272 3000 216278 3012
rect 217137 3009 217149 3043
rect 217183 3040 217195 3043
rect 217962 3040 217968 3052
rect 217183 3012 217968 3040
rect 217183 3009 217195 3012
rect 217137 3003 217195 3009
rect 217962 3000 217968 3012
rect 218020 3040 218026 3052
rect 218020 3012 218652 3040
rect 218020 3000 218026 3012
rect 209148 2944 209774 2972
rect 209041 2935 209099 2941
rect 210234 2932 210240 2984
rect 210292 2932 210298 2984
rect 211430 2932 211436 2984
rect 211488 2932 211494 2984
rect 212534 2932 212540 2984
rect 212592 2972 212598 2984
rect 215389 2975 215447 2981
rect 215389 2972 215401 2975
rect 212592 2944 215401 2972
rect 212592 2932 212598 2944
rect 215389 2941 215401 2944
rect 215435 2941 215447 2975
rect 215389 2935 215447 2941
rect 121932 2876 125456 2904
rect 29052 2808 37596 2836
rect 29052 2796 29058 2808
rect 37642 2796 37648 2848
rect 37700 2796 37706 2848
rect 74537 2839 74595 2845
rect 74537 2805 74549 2839
rect 74583 2836 74595 2839
rect 74718 2836 74724 2848
rect 74583 2808 74724 2836
rect 74583 2805 74595 2808
rect 74537 2799 74595 2805
rect 74718 2796 74724 2808
rect 74776 2796 74782 2848
rect 74994 2796 75000 2848
rect 75052 2796 75058 2848
rect 108209 2839 108267 2845
rect 108209 2805 108221 2839
rect 108255 2836 108267 2839
rect 108390 2836 108396 2848
rect 108255 2808 108396 2836
rect 108255 2805 108267 2808
rect 108209 2799 108267 2805
rect 108390 2796 108396 2808
rect 108448 2796 108454 2848
rect 112165 2839 112223 2845
rect 112165 2805 112177 2839
rect 112211 2836 112223 2839
rect 112346 2836 112352 2848
rect 112211 2808 112352 2836
rect 112211 2805 112223 2808
rect 112165 2799 112223 2805
rect 112346 2796 112352 2808
rect 112404 2796 112410 2848
rect 112993 2839 113051 2845
rect 112993 2805 113005 2839
rect 113039 2836 113051 2839
rect 114186 2836 114192 2848
rect 113039 2808 114192 2836
rect 113039 2805 113051 2808
rect 112993 2799 113051 2805
rect 114186 2796 114192 2808
rect 114244 2796 114250 2848
rect 118050 2796 118056 2848
rect 118108 2836 118114 2848
rect 124582 2836 124588 2848
rect 118108 2808 124588 2836
rect 118108 2796 118114 2808
rect 124582 2796 124588 2808
rect 124640 2796 124646 2848
rect 125428 2836 125456 2876
rect 126054 2864 126060 2916
rect 126112 2904 126118 2916
rect 126701 2907 126759 2913
rect 126701 2904 126713 2907
rect 126112 2876 126713 2904
rect 126112 2864 126118 2876
rect 126701 2873 126713 2876
rect 126747 2873 126759 2907
rect 126701 2867 126759 2873
rect 126882 2864 126888 2916
rect 126940 2904 126946 2916
rect 214006 2904 214012 2916
rect 126940 2876 214012 2904
rect 126940 2864 126946 2876
rect 214006 2864 214012 2876
rect 214064 2864 214070 2916
rect 218624 2904 218652 3012
rect 218698 3000 218704 3052
rect 218756 3000 218762 3052
rect 218808 2972 218836 3080
rect 219894 3068 219900 3120
rect 219952 3068 219958 3120
rect 219253 3043 219311 3049
rect 219253 3009 219265 3043
rect 219299 3040 219311 3043
rect 219526 3040 219532 3052
rect 219299 3012 219532 3040
rect 219299 3009 219311 3012
rect 219253 3003 219311 3009
rect 219526 3000 219532 3012
rect 219584 3000 219590 3052
rect 220449 3043 220507 3049
rect 220449 3009 220461 3043
rect 220495 3040 220507 3043
rect 221108 3040 221136 3136
rect 220495 3012 221136 3040
rect 221200 3080 307340 3108
rect 220495 3009 220507 3012
rect 220449 3003 220507 3009
rect 221200 2972 221228 3080
rect 221366 3000 221372 3052
rect 221424 3040 221430 3052
rect 221424 3012 224954 3040
rect 221424 3000 221430 3012
rect 218808 2944 221228 2972
rect 221182 2904 221188 2916
rect 218624 2876 221188 2904
rect 221182 2864 221188 2876
rect 221240 2864 221246 2916
rect 224926 2904 224954 3012
rect 254026 3000 254032 3052
rect 254084 3000 254090 3052
rect 259086 3000 259092 3052
rect 259144 3000 259150 3052
rect 259641 3043 259699 3049
rect 259641 3009 259653 3043
rect 259687 3040 259699 3043
rect 260282 3040 260288 3052
rect 259687 3012 260288 3040
rect 259687 3009 259699 3012
rect 259641 3003 259699 3009
rect 260282 3000 260288 3012
rect 260340 3000 260346 3052
rect 296530 3000 296536 3052
rect 296588 3000 296594 3052
rect 297358 3000 297364 3052
rect 297416 3040 297422 3052
rect 298005 3043 298063 3049
rect 298005 3040 298017 3043
rect 297416 3012 298017 3040
rect 297416 3000 297422 3012
rect 298005 3009 298017 3012
rect 298051 3009 298063 3043
rect 298005 3003 298063 3009
rect 298646 3000 298652 3052
rect 298704 3000 298710 3052
rect 300210 3000 300216 3052
rect 300268 3000 300274 3052
rect 300581 3043 300639 3049
rect 300581 3009 300593 3043
rect 300627 3040 300639 3043
rect 300854 3040 300860 3052
rect 300627 3012 300860 3040
rect 300627 3009 300639 3012
rect 300581 3003 300639 3009
rect 300854 3000 300860 3012
rect 300912 3000 300918 3052
rect 301130 3000 301136 3052
rect 301188 3000 301194 3052
rect 301222 3000 301228 3052
rect 301280 3040 301286 3052
rect 303157 3043 303215 3049
rect 301280 3012 303108 3040
rect 301280 3000 301286 3012
rect 302881 2975 302939 2981
rect 302881 2972 302893 2975
rect 296686 2944 302893 2972
rect 296686 2904 296714 2944
rect 302881 2941 302893 2944
rect 302927 2941 302939 2975
rect 303080 2972 303108 3012
rect 303157 3009 303169 3043
rect 303203 3040 303215 3043
rect 303430 3040 303436 3052
rect 303203 3012 303436 3040
rect 303203 3009 303215 3012
rect 303157 3003 303215 3009
rect 303430 3000 303436 3012
rect 303488 3000 303494 3052
rect 303540 3012 304304 3040
rect 303540 2972 303568 3012
rect 303080 2944 303568 2972
rect 302881 2935 302939 2941
rect 303798 2932 303804 2984
rect 303856 2932 303862 2984
rect 304276 2972 304304 3012
rect 304350 3000 304356 3052
rect 304408 3000 304414 3052
rect 305825 3043 305883 3049
rect 304460 3012 305776 3040
rect 304460 2972 304488 3012
rect 304276 2944 304488 2972
rect 305362 2932 305368 2984
rect 305420 2972 305426 2984
rect 305549 2975 305607 2981
rect 305549 2972 305561 2975
rect 305420 2944 305561 2972
rect 305420 2932 305426 2944
rect 305549 2941 305561 2944
rect 305595 2941 305607 2975
rect 305748 2972 305776 3012
rect 305825 3009 305837 3043
rect 305871 3040 305883 3043
rect 306190 3040 306196 3052
rect 305871 3012 306196 3040
rect 305871 3009 305883 3012
rect 305825 3003 305883 3009
rect 306190 3000 306196 3012
rect 306248 3000 306254 3052
rect 306558 3040 306564 3052
rect 306346 3012 306564 3040
rect 306346 2972 306374 3012
rect 306558 3000 306564 3012
rect 306616 3000 306622 3052
rect 306653 3043 306711 3049
rect 306653 3009 306665 3043
rect 306699 3040 306711 3043
rect 306834 3040 306840 3052
rect 306699 3012 306840 3040
rect 306699 3009 306711 3012
rect 306653 3003 306711 3009
rect 306834 3000 306840 3012
rect 306892 3000 306898 3052
rect 305748 2944 306374 2972
rect 305549 2935 305607 2941
rect 224926 2876 296714 2904
rect 297545 2907 297603 2913
rect 297545 2873 297557 2907
rect 297591 2904 297603 2907
rect 301222 2904 301228 2916
rect 297591 2876 301228 2904
rect 297591 2873 297603 2876
rect 297545 2867 297603 2873
rect 301222 2864 301228 2876
rect 301280 2864 301286 2916
rect 301317 2907 301375 2913
rect 301317 2873 301329 2907
rect 301363 2904 301375 2907
rect 306469 2907 306527 2913
rect 301363 2876 306374 2904
rect 301363 2873 301375 2876
rect 301317 2867 301375 2873
rect 127434 2836 127440 2848
rect 125428 2808 127440 2836
rect 127434 2796 127440 2808
rect 127492 2796 127498 2848
rect 143166 2796 143172 2848
rect 143224 2796 143230 2848
rect 152182 2796 152188 2848
rect 152240 2836 152246 2848
rect 152277 2839 152335 2845
rect 152277 2836 152289 2839
rect 152240 2808 152289 2836
rect 152240 2796 152246 2808
rect 152277 2805 152289 2808
rect 152323 2805 152335 2839
rect 152277 2799 152335 2805
rect 164786 2796 164792 2848
rect 164844 2796 164850 2848
rect 168006 2796 168012 2848
rect 168064 2796 168070 2848
rect 201678 2796 201684 2848
rect 201736 2796 201742 2848
rect 206097 2839 206155 2845
rect 206097 2805 206109 2839
rect 206143 2836 206155 2839
rect 206186 2836 206192 2848
rect 206143 2808 206192 2836
rect 206143 2805 206155 2808
rect 206097 2799 206155 2805
rect 206186 2796 206192 2808
rect 206244 2796 206250 2848
rect 206830 2796 206836 2848
rect 206888 2796 206894 2848
rect 218149 2839 218207 2845
rect 218149 2805 218161 2839
rect 218195 2836 218207 2839
rect 218422 2836 218428 2848
rect 218195 2808 218428 2836
rect 218195 2805 218207 2808
rect 218149 2799 218207 2805
rect 218422 2796 218428 2808
rect 218480 2796 218486 2848
rect 221642 2796 221648 2848
rect 221700 2796 221706 2848
rect 247126 2796 247132 2848
rect 247184 2836 247190 2848
rect 247221 2839 247279 2845
rect 247221 2836 247233 2839
rect 247184 2808 247233 2836
rect 247184 2796 247190 2808
rect 247221 2805 247233 2808
rect 247267 2805 247279 2839
rect 247221 2799 247279 2805
rect 251545 2839 251603 2845
rect 251545 2805 251557 2839
rect 251591 2836 251603 2839
rect 251726 2836 251732 2848
rect 251591 2808 251732 2836
rect 251591 2805 251603 2808
rect 251545 2799 251603 2805
rect 251726 2796 251732 2808
rect 251784 2796 251790 2848
rect 260282 2796 260288 2848
rect 260340 2796 260346 2848
rect 295794 2796 295800 2848
rect 295852 2836 295858 2848
rect 295981 2839 296039 2845
rect 295981 2836 295993 2839
rect 295852 2808 295993 2836
rect 295852 2796 295858 2808
rect 295981 2805 295993 2808
rect 296027 2805 296039 2839
rect 295981 2799 296039 2805
rect 299566 2796 299572 2848
rect 299624 2796 299630 2848
rect 301130 2796 301136 2848
rect 301188 2836 301194 2848
rect 301777 2839 301835 2845
rect 301777 2836 301789 2839
rect 301188 2808 301789 2836
rect 301188 2796 301194 2808
rect 301777 2805 301789 2808
rect 301823 2805 301835 2839
rect 301777 2799 301835 2805
rect 304350 2796 304356 2848
rect 304408 2836 304414 2848
rect 305454 2836 305460 2848
rect 304408 2808 305460 2836
rect 304408 2796 304414 2808
rect 305454 2796 305460 2808
rect 305512 2796 305518 2848
rect 306346 2836 306374 2876
rect 306469 2873 306481 2907
rect 306515 2904 306527 2907
rect 306650 2904 306656 2916
rect 306515 2876 306656 2904
rect 306515 2873 306527 2876
rect 306469 2867 306527 2873
rect 306650 2864 306656 2876
rect 306708 2864 306714 2916
rect 307312 2904 307340 3080
rect 307386 3068 307392 3120
rect 307444 3068 307450 3120
rect 309410 3068 309416 3120
rect 309468 3068 309474 3120
rect 310698 3068 310704 3120
rect 310756 3068 310762 3120
rect 342162 3108 342168 3120
rect 310992 3080 321554 3108
rect 307665 3043 307723 3049
rect 307665 3009 307677 3043
rect 307711 3040 307723 3043
rect 307846 3040 307852 3052
rect 307711 3012 307852 3040
rect 307711 3009 307723 3012
rect 307665 3003 307723 3009
rect 307846 3000 307852 3012
rect 307904 3000 307910 3052
rect 308582 3000 308588 3052
rect 308640 3000 308646 3052
rect 310992 3049 311020 3080
rect 310977 3043 311035 3049
rect 310977 3009 310989 3043
rect 311023 3009 311035 3043
rect 311897 3043 311955 3049
rect 310977 3003 311035 3009
rect 311084 3012 311756 3040
rect 307386 2932 307392 2984
rect 307444 2972 307450 2984
rect 308309 2975 308367 2981
rect 308309 2972 308321 2975
rect 307444 2944 308321 2972
rect 307444 2932 307450 2944
rect 308309 2941 308321 2944
rect 308355 2941 308367 2975
rect 308309 2935 308367 2941
rect 308490 2932 308496 2984
rect 308548 2972 308554 2984
rect 311084 2972 311112 3012
rect 308548 2944 311112 2972
rect 311621 2975 311679 2981
rect 308548 2932 308554 2944
rect 311621 2941 311633 2975
rect 311667 2941 311679 2975
rect 311728 2972 311756 3012
rect 311897 3009 311909 3043
rect 311943 3040 311955 3043
rect 311943 3012 312676 3040
rect 311943 3009 311955 3012
rect 311897 3003 311955 3009
rect 312449 2975 312507 2981
rect 312449 2972 312461 2975
rect 311728 2944 312461 2972
rect 311621 2935 311679 2941
rect 312449 2941 312461 2944
rect 312495 2941 312507 2975
rect 312648 2972 312676 3012
rect 312722 3000 312728 3052
rect 312780 3000 312786 3052
rect 314010 3000 314016 3052
rect 314068 3040 314074 3052
rect 314565 3043 314623 3049
rect 314565 3040 314577 3043
rect 314068 3012 314577 3040
rect 314068 3000 314074 3012
rect 314565 3009 314577 3012
rect 314611 3009 314623 3043
rect 314565 3003 314623 3009
rect 317325 3043 317383 3049
rect 317325 3009 317337 3043
rect 317371 3040 317383 3043
rect 317874 3040 317880 3052
rect 317371 3012 317880 3040
rect 317371 3009 317383 3012
rect 317325 3003 317383 3009
rect 317874 3000 317880 3012
rect 317932 3000 317938 3052
rect 312648 2944 313872 2972
rect 312449 2935 312507 2941
rect 311636 2904 311664 2935
rect 313844 2904 313872 2944
rect 315758 2932 315764 2984
rect 315816 2932 315822 2984
rect 321526 2972 321554 3080
rect 325666 3080 342168 3108
rect 323394 2972 323400 2984
rect 321526 2944 323400 2972
rect 323394 2932 323400 2944
rect 323452 2932 323458 2984
rect 317141 2907 317199 2913
rect 317141 2904 317153 2907
rect 307312 2876 311664 2904
rect 311866 2876 313504 2904
rect 313844 2876 317153 2904
rect 307754 2836 307760 2848
rect 306346 2808 307760 2836
rect 307754 2796 307760 2808
rect 307812 2796 307818 2848
rect 309042 2796 309048 2848
rect 309100 2836 309106 2848
rect 311866 2836 311894 2876
rect 309100 2808 311894 2836
rect 309100 2796 309106 2808
rect 313366 2796 313372 2848
rect 313424 2796 313430 2848
rect 313476 2836 313504 2876
rect 317141 2873 317153 2876
rect 317187 2873 317199 2907
rect 325666 2904 325694 3080
rect 342162 3068 342168 3080
rect 342220 3068 342226 3120
rect 344388 3117 344416 3148
rect 345017 3145 345029 3148
rect 345063 3176 345075 3179
rect 348234 3176 348240 3188
rect 345063 3148 348240 3176
rect 345063 3145 345075 3148
rect 345017 3139 345075 3145
rect 348234 3136 348240 3148
rect 348292 3136 348298 3188
rect 350718 3136 350724 3188
rect 350776 3176 350782 3188
rect 353297 3179 353355 3185
rect 353297 3176 353309 3179
rect 350776 3148 353309 3176
rect 350776 3136 350782 3148
rect 353297 3145 353309 3148
rect 353343 3176 353355 3179
rect 353343 3148 353800 3176
rect 353343 3145 353355 3148
rect 353297 3139 353355 3145
rect 344373 3111 344431 3117
rect 344373 3077 344385 3111
rect 344419 3077 344431 3111
rect 344373 3071 344431 3077
rect 331401 3043 331459 3049
rect 331401 3009 331413 3043
rect 331447 3009 331459 3043
rect 331401 3003 331459 3009
rect 340141 3043 340199 3049
rect 340141 3009 340153 3043
rect 340187 3040 340199 3043
rect 340785 3043 340843 3049
rect 340785 3040 340797 3043
rect 340187 3012 340797 3040
rect 340187 3009 340199 3012
rect 340141 3003 340199 3009
rect 340785 3009 340797 3012
rect 340831 3040 340843 3043
rect 353294 3040 353300 3052
rect 340831 3012 353300 3040
rect 340831 3009 340843 3012
rect 340785 3003 340843 3009
rect 317141 2867 317199 2873
rect 317248 2876 325694 2904
rect 331416 2904 331444 3003
rect 353294 3000 353300 3012
rect 353352 3000 353358 3052
rect 353772 3049 353800 3148
rect 353938 3136 353944 3188
rect 353996 3136 354002 3188
rect 357529 3179 357587 3185
rect 357529 3145 357541 3179
rect 357575 3176 357587 3179
rect 357575 3148 364334 3176
rect 357575 3145 357587 3148
rect 357529 3139 357587 3145
rect 362218 3068 362224 3120
rect 362276 3068 362282 3120
rect 364306 3108 364334 3148
rect 382734 3136 382740 3188
rect 382792 3176 382798 3188
rect 478874 3176 478880 3188
rect 382792 3148 478880 3176
rect 382792 3136 382798 3148
rect 478874 3136 478880 3148
rect 478932 3136 478938 3188
rect 411070 3108 411076 3120
rect 364306 3080 411076 3108
rect 411070 3068 411076 3080
rect 411128 3068 411134 3120
rect 416314 3068 416320 3120
rect 416372 3068 416378 3120
rect 422570 3068 422576 3120
rect 422628 3108 422634 3120
rect 499758 3108 499764 3120
rect 422628 3080 499764 3108
rect 422628 3068 422634 3080
rect 499758 3068 499764 3080
rect 499816 3068 499822 3120
rect 353757 3043 353815 3049
rect 353757 3009 353769 3043
rect 353803 3009 353815 3043
rect 357158 3040 357164 3052
rect 353757 3003 353815 3009
rect 353864 3012 357164 3040
rect 340874 2932 340880 2984
rect 340932 2972 340938 2984
rect 340932 2944 349936 2972
rect 340932 2932 340938 2944
rect 332045 2907 332103 2913
rect 332045 2904 332057 2907
rect 331416 2876 332057 2904
rect 317248 2836 317276 2876
rect 332045 2873 332057 2876
rect 332091 2904 332103 2907
rect 349798 2904 349804 2916
rect 332091 2876 349804 2904
rect 332091 2873 332103 2876
rect 332045 2867 332103 2873
rect 349798 2864 349804 2876
rect 349856 2864 349862 2916
rect 349908 2904 349936 2944
rect 353864 2904 353892 3012
rect 357158 3000 357164 3012
rect 357216 3040 357222 3052
rect 357345 3043 357403 3049
rect 357345 3040 357357 3043
rect 357216 3012 357357 3040
rect 357216 3000 357222 3012
rect 357345 3009 357357 3012
rect 357391 3009 357403 3043
rect 357345 3003 357403 3009
rect 390186 3000 390192 3052
rect 390244 3000 390250 3052
rect 390554 3000 390560 3052
rect 390612 3000 390618 3052
rect 392949 3043 393007 3049
rect 392949 3040 392961 3043
rect 391032 3012 392961 3040
rect 354030 2932 354036 2984
rect 354088 2972 354094 2984
rect 391032 2972 391060 3012
rect 392949 3009 392961 3012
rect 392995 3009 393007 3043
rect 392949 3003 393007 3009
rect 393317 3043 393375 3049
rect 393317 3009 393329 3043
rect 393363 3009 393375 3043
rect 393317 3003 393375 3009
rect 354088 2944 391060 2972
rect 354088 2932 354094 2944
rect 391106 2932 391112 2984
rect 391164 2972 391170 2984
rect 391661 2975 391719 2981
rect 391661 2972 391673 2975
rect 391164 2944 391673 2972
rect 391164 2932 391170 2944
rect 391661 2941 391673 2944
rect 391707 2941 391719 2975
rect 393332 2972 393360 3003
rect 394234 3000 394240 3052
rect 394292 3040 394298 3052
rect 394418 3040 394424 3052
rect 394292 3012 394424 3040
rect 394292 3000 394298 3012
rect 394418 3000 394424 3012
rect 394476 3000 394482 3052
rect 396074 3040 396080 3052
rect 394528 3012 396080 3040
rect 393590 2972 393596 2984
rect 393332 2944 393596 2972
rect 391661 2935 391719 2941
rect 393590 2932 393596 2944
rect 393648 2972 393654 2984
rect 394528 2972 394556 3012
rect 396074 3000 396080 3012
rect 396132 3000 396138 3052
rect 396718 3000 396724 3052
rect 396776 3000 396782 3052
rect 397089 3043 397147 3049
rect 397089 3009 397101 3043
rect 397135 3040 397147 3043
rect 398101 3043 398159 3049
rect 398101 3040 398113 3043
rect 397135 3012 398113 3040
rect 397135 3009 397147 3012
rect 397089 3003 397147 3009
rect 398101 3009 398113 3012
rect 398147 3040 398159 3043
rect 401778 3040 401784 3052
rect 398147 3012 401784 3040
rect 398147 3009 398159 3012
rect 398101 3003 398159 3009
rect 401778 3000 401784 3012
rect 401836 3000 401842 3052
rect 452841 3043 452899 3049
rect 431926 3012 452792 3040
rect 393648 2944 394556 2972
rect 394973 2975 395031 2981
rect 393648 2932 393654 2944
rect 394973 2941 394985 2975
rect 395019 2972 395031 2975
rect 431926 2972 431954 3012
rect 452565 2975 452623 2981
rect 452565 2972 452577 2975
rect 395019 2944 431954 2972
rect 451246 2944 452577 2972
rect 395019 2941 395031 2944
rect 394973 2935 395031 2941
rect 349908 2876 353892 2904
rect 359550 2864 359556 2916
rect 359608 2904 359614 2916
rect 451246 2904 451274 2944
rect 452565 2941 452577 2944
rect 452611 2941 452623 2975
rect 452764 2972 452792 3012
rect 452841 3009 452853 3043
rect 452887 3040 452899 3043
rect 453393 3043 453451 3049
rect 453393 3040 453405 3043
rect 452887 3012 453405 3040
rect 452887 3009 452899 3012
rect 452841 3003 452899 3009
rect 453393 3009 453405 3012
rect 453439 3040 453451 3043
rect 484578 3040 484584 3052
rect 453439 3012 484584 3040
rect 453439 3009 453451 3012
rect 453393 3003 453451 3009
rect 484578 3000 484584 3012
rect 484636 3000 484642 3052
rect 488626 2972 488632 2984
rect 452764 2944 488632 2972
rect 452565 2935 452623 2941
rect 488626 2932 488632 2944
rect 488684 2932 488690 2984
rect 359608 2876 451274 2904
rect 359608 2864 359614 2876
rect 470410 2864 470416 2916
rect 470468 2864 470474 2916
rect 313476 2808 317276 2836
rect 318978 2796 318984 2848
rect 319036 2836 319042 2848
rect 319073 2839 319131 2845
rect 319073 2836 319085 2839
rect 319036 2808 319085 2836
rect 319036 2796 319042 2808
rect 319073 2805 319085 2808
rect 319119 2805 319131 2839
rect 319073 2799 319131 2805
rect 319438 2796 319444 2848
rect 319496 2836 319502 2848
rect 319625 2839 319683 2845
rect 319625 2836 319637 2839
rect 319496 2808 319637 2836
rect 319496 2796 319502 2808
rect 319625 2805 319637 2808
rect 319671 2805 319683 2839
rect 319625 2799 319683 2805
rect 323762 2796 323768 2848
rect 323820 2796 323826 2848
rect 324682 2796 324688 2848
rect 324740 2836 324746 2848
rect 324777 2839 324835 2845
rect 324777 2836 324789 2839
rect 324740 2808 324789 2836
rect 324740 2796 324746 2808
rect 324777 2805 324789 2808
rect 324823 2805 324835 2839
rect 324777 2799 324835 2805
rect 325142 2796 325148 2848
rect 325200 2836 325206 2848
rect 325329 2839 325387 2845
rect 325329 2836 325341 2839
rect 325200 2808 325341 2836
rect 325200 2796 325206 2808
rect 325329 2805 325341 2808
rect 325375 2805 325387 2839
rect 325329 2799 325387 2805
rect 332597 2839 332655 2845
rect 332597 2805 332609 2839
rect 332643 2836 332655 2839
rect 332778 2836 332784 2848
rect 332643 2808 332784 2836
rect 332643 2805 332655 2808
rect 332597 2799 332655 2805
rect 332778 2796 332784 2808
rect 332836 2796 332842 2848
rect 337286 2796 337292 2848
rect 337344 2836 337350 2848
rect 337473 2839 337531 2845
rect 337473 2836 337485 2839
rect 337344 2808 337485 2836
rect 337344 2796 337350 2808
rect 337473 2805 337485 2808
rect 337519 2805 337531 2839
rect 337473 2799 337531 2805
rect 337838 2796 337844 2848
rect 337896 2836 337902 2848
rect 338117 2839 338175 2845
rect 338117 2836 338129 2839
rect 337896 2808 338129 2836
rect 337896 2796 337902 2808
rect 338117 2805 338129 2808
rect 338163 2805 338175 2839
rect 338117 2799 338175 2805
rect 341518 2796 341524 2848
rect 341576 2796 341582 2848
rect 342070 2796 342076 2848
rect 342128 2796 342134 2848
rect 345566 2796 345572 2848
rect 345624 2796 345630 2848
rect 346670 2796 346676 2848
rect 346728 2796 346734 2848
rect 348418 2796 348424 2848
rect 348476 2836 348482 2848
rect 348605 2839 348663 2845
rect 348605 2836 348617 2839
rect 348476 2808 348617 2836
rect 348476 2796 348482 2808
rect 348605 2805 348617 2808
rect 348651 2805 348663 2839
rect 348605 2799 348663 2805
rect 349706 2796 349712 2848
rect 349764 2836 349770 2848
rect 349893 2839 349951 2845
rect 349893 2836 349905 2839
rect 349764 2808 349905 2836
rect 349764 2796 349770 2808
rect 349893 2805 349905 2808
rect 349939 2805 349951 2839
rect 349893 2799 349951 2805
rect 350537 2839 350595 2845
rect 350537 2805 350549 2839
rect 350583 2836 350595 2839
rect 350626 2836 350632 2848
rect 350583 2808 350632 2836
rect 350583 2805 350595 2808
rect 350537 2799 350595 2805
rect 350626 2796 350632 2808
rect 350684 2796 350690 2848
rect 352374 2796 352380 2848
rect 352432 2836 352438 2848
rect 352561 2839 352619 2845
rect 352561 2836 352573 2839
rect 352432 2808 352573 2836
rect 352432 2796 352438 2808
rect 352561 2805 352573 2808
rect 352607 2805 352619 2839
rect 352561 2799 352619 2805
rect 353662 2796 353668 2848
rect 353720 2836 353726 2848
rect 354490 2836 354496 2848
rect 353720 2808 354496 2836
rect 353720 2796 353726 2808
rect 354490 2796 354496 2808
rect 354548 2796 354554 2848
rect 356054 2796 356060 2848
rect 356112 2836 356118 2848
rect 356149 2839 356207 2845
rect 356149 2836 356161 2839
rect 356112 2808 356161 2836
rect 356112 2796 356118 2808
rect 356149 2805 356161 2808
rect 356195 2805 356207 2839
rect 356149 2799 356207 2805
rect 358170 2796 358176 2848
rect 358228 2796 358234 2848
rect 380894 2796 380900 2848
rect 380952 2796 380958 2848
rect 390554 2796 390560 2848
rect 390612 2836 390618 2848
rect 391201 2839 391259 2845
rect 391201 2836 391213 2839
rect 390612 2808 391213 2836
rect 390612 2796 390618 2808
rect 391201 2805 391213 2808
rect 391247 2836 391259 2839
rect 395982 2836 395988 2848
rect 391247 2808 395988 2836
rect 391247 2805 391259 2808
rect 391201 2799 391259 2805
rect 395982 2796 395988 2808
rect 396040 2796 396046 2848
rect 396166 2796 396172 2848
rect 396224 2796 396230 2848
rect 398926 2796 398932 2848
rect 398984 2796 398990 2848
rect 399846 2796 399852 2848
rect 399904 2836 399910 2848
rect 400033 2839 400091 2845
rect 400033 2836 400045 2839
rect 399904 2808 400045 2836
rect 399904 2796 399910 2808
rect 400033 2805 400045 2808
rect 400079 2805 400091 2839
rect 400033 2799 400091 2805
rect 400953 2839 401011 2845
rect 400953 2805 400965 2839
rect 400999 2836 401011 2839
rect 401134 2836 401140 2848
rect 400999 2808 401140 2836
rect 400999 2805 401011 2808
rect 400953 2799 401011 2805
rect 401134 2796 401140 2808
rect 401192 2796 401198 2848
rect 408494 2796 408500 2848
rect 408552 2796 408558 2848
rect 434990 2796 434996 2848
rect 435048 2796 435054 2848
rect 435726 2796 435732 2848
rect 435784 2836 435790 2848
rect 435821 2839 435879 2845
rect 435821 2836 435833 2839
rect 435784 2808 435833 2836
rect 435784 2796 435790 2808
rect 435821 2805 435833 2808
rect 435867 2805 435879 2839
rect 435821 2799 435879 2805
rect 1104 2746 528816 2768
rect 1104 2694 66914 2746
rect 66966 2694 66978 2746
rect 67030 2694 67042 2746
rect 67094 2694 67106 2746
rect 67158 2694 67170 2746
rect 67222 2694 198842 2746
rect 198894 2694 198906 2746
rect 198958 2694 198970 2746
rect 199022 2694 199034 2746
rect 199086 2694 199098 2746
rect 199150 2694 330770 2746
rect 330822 2694 330834 2746
rect 330886 2694 330898 2746
rect 330950 2694 330962 2746
rect 331014 2694 331026 2746
rect 331078 2694 462698 2746
rect 462750 2694 462762 2746
rect 462814 2694 462826 2746
rect 462878 2694 462890 2746
rect 462942 2694 462954 2746
rect 463006 2694 528816 2746
rect 1104 2672 528816 2694
rect 1854 2592 1860 2644
rect 1912 2592 1918 2644
rect 19886 2592 19892 2644
rect 19944 2592 19950 2644
rect 29178 2592 29184 2644
rect 29236 2632 29242 2644
rect 29236 2604 45554 2632
rect 29236 2592 29242 2604
rect 45526 2564 45554 2604
rect 53834 2592 53840 2644
rect 53892 2632 53898 2644
rect 55953 2635 56011 2641
rect 55953 2632 55965 2635
rect 53892 2604 55965 2632
rect 53892 2592 53898 2604
rect 55953 2601 55965 2604
rect 55999 2601 56011 2635
rect 55953 2595 56011 2601
rect 58158 2592 58164 2644
rect 58216 2592 58222 2644
rect 63586 2632 63592 2644
rect 58268 2604 63592 2632
rect 56502 2564 56508 2576
rect 45526 2536 56508 2564
rect 56502 2524 56508 2536
rect 56560 2524 56566 2576
rect 56689 2567 56747 2573
rect 56689 2533 56701 2567
rect 56735 2564 56747 2567
rect 58268 2564 58296 2604
rect 63586 2592 63592 2604
rect 63644 2592 63650 2644
rect 70394 2592 70400 2644
rect 70452 2632 70458 2644
rect 71038 2632 71044 2644
rect 70452 2604 71044 2632
rect 70452 2592 70458 2604
rect 71038 2592 71044 2604
rect 71096 2592 71102 2644
rect 73982 2592 73988 2644
rect 74040 2592 74046 2644
rect 74534 2592 74540 2644
rect 74592 2632 74598 2644
rect 164786 2632 164792 2644
rect 74592 2604 164792 2632
rect 74592 2592 74598 2604
rect 164786 2592 164792 2604
rect 164844 2592 164850 2644
rect 179414 2592 179420 2644
rect 179472 2632 179478 2644
rect 182177 2635 182235 2641
rect 182177 2632 182189 2635
rect 179472 2604 182189 2632
rect 179472 2592 179478 2604
rect 182177 2601 182189 2604
rect 182223 2601 182235 2635
rect 182177 2595 182235 2601
rect 211798 2592 211804 2644
rect 211856 2632 211862 2644
rect 211856 2604 301360 2632
rect 211856 2592 211862 2604
rect 143166 2564 143172 2576
rect 56735 2536 58296 2564
rect 58912 2536 143172 2564
rect 56735 2533 56747 2536
rect 56689 2527 56747 2533
rect 21910 2456 21916 2508
rect 21968 2496 21974 2508
rect 55858 2496 55864 2508
rect 21968 2468 55864 2496
rect 21968 2456 21974 2468
rect 55858 2456 55864 2468
rect 55916 2456 55922 2508
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2428 2099 2431
rect 20073 2431 20131 2437
rect 2087 2400 2636 2428
rect 2087 2397 2099 2400
rect 2041 2391 2099 2397
rect 2608 2304 2636 2400
rect 20073 2397 20085 2431
rect 20119 2428 20131 2431
rect 20625 2431 20683 2437
rect 20625 2428 20637 2431
rect 20119 2400 20637 2428
rect 20119 2397 20131 2400
rect 20073 2391 20131 2397
rect 20625 2397 20637 2400
rect 20671 2428 20683 2431
rect 31754 2428 31760 2440
rect 20671 2400 31760 2428
rect 20671 2397 20683 2400
rect 20625 2391 20683 2397
rect 31754 2388 31760 2400
rect 31812 2388 31818 2440
rect 35894 2388 35900 2440
rect 35952 2428 35958 2440
rect 36438 2431 36496 2437
rect 36438 2428 36450 2431
rect 35952 2400 36450 2428
rect 35952 2388 35958 2400
rect 36438 2397 36450 2400
rect 36484 2397 36496 2431
rect 36438 2391 36496 2397
rect 37642 2388 37648 2440
rect 37700 2428 37706 2440
rect 38105 2431 38163 2437
rect 38105 2428 38117 2431
rect 37700 2400 38117 2428
rect 37700 2388 37706 2400
rect 38105 2397 38117 2400
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 41966 2388 41972 2440
rect 42024 2428 42030 2440
rect 42613 2431 42671 2437
rect 42613 2428 42625 2431
rect 42024 2400 42625 2428
rect 42024 2388 42030 2400
rect 42613 2397 42625 2400
rect 42659 2397 42671 2431
rect 42613 2391 42671 2397
rect 48314 2388 48320 2440
rect 48372 2428 48378 2440
rect 48869 2431 48927 2437
rect 48869 2428 48881 2431
rect 48372 2400 48881 2428
rect 48372 2388 48378 2400
rect 48869 2397 48881 2400
rect 48915 2397 48927 2431
rect 53837 2431 53895 2437
rect 53837 2428 53849 2431
rect 48869 2391 48927 2397
rect 49068 2400 53849 2428
rect 24302 2320 24308 2372
rect 24360 2360 24366 2372
rect 24360 2332 36584 2360
rect 24360 2320 24366 2332
rect 2590 2252 2596 2304
rect 2648 2252 2654 2304
rect 26694 2252 26700 2304
rect 26752 2292 26758 2304
rect 35894 2292 35900 2304
rect 26752 2264 35900 2292
rect 26752 2252 26758 2264
rect 35894 2252 35900 2264
rect 35952 2252 35958 2304
rect 36556 2292 36584 2332
rect 36722 2320 36728 2372
rect 36780 2320 36786 2372
rect 36832 2332 42104 2360
rect 36832 2292 36860 2332
rect 36556 2264 36860 2292
rect 37918 2252 37924 2304
rect 37976 2252 37982 2304
rect 41966 2252 41972 2304
rect 42024 2252 42030 2304
rect 42076 2292 42104 2332
rect 42886 2320 42892 2372
rect 42944 2320 42950 2372
rect 49068 2360 49096 2400
rect 53837 2397 53849 2400
rect 53883 2428 53895 2431
rect 54389 2431 54447 2437
rect 54389 2428 54401 2431
rect 53883 2400 54401 2428
rect 53883 2397 53895 2400
rect 53837 2391 53895 2397
rect 54389 2397 54401 2400
rect 54435 2397 54447 2431
rect 54389 2391 54447 2397
rect 54662 2388 54668 2440
rect 54720 2388 54726 2440
rect 56137 2431 56195 2437
rect 56137 2397 56149 2431
rect 56183 2428 56195 2431
rect 56704 2428 56732 2527
rect 56183 2400 56732 2428
rect 56183 2397 56195 2400
rect 56137 2391 56195 2397
rect 58158 2388 58164 2440
rect 58216 2428 58222 2440
rect 58713 2431 58771 2437
rect 58713 2428 58725 2431
rect 58216 2400 58725 2428
rect 58216 2388 58222 2400
rect 58713 2397 58725 2400
rect 58759 2397 58771 2431
rect 58713 2391 58771 2397
rect 45526 2332 49096 2360
rect 49145 2363 49203 2369
rect 45526 2292 45554 2332
rect 49145 2329 49157 2363
rect 49191 2360 49203 2363
rect 58912 2360 58940 2536
rect 143166 2524 143172 2536
rect 143224 2524 143230 2576
rect 148226 2524 148232 2576
rect 148284 2524 148290 2576
rect 242897 2567 242955 2573
rect 242897 2564 242909 2567
rect 149348 2536 242909 2564
rect 71593 2499 71651 2505
rect 60706 2468 70900 2496
rect 49191 2332 58940 2360
rect 49191 2329 49203 2332
rect 49145 2323 49203 2329
rect 58986 2320 58992 2372
rect 59044 2320 59050 2372
rect 42076 2264 45554 2292
rect 48314 2252 48320 2304
rect 48372 2252 48378 2304
rect 55858 2252 55864 2304
rect 55916 2292 55922 2304
rect 60706 2292 60734 2468
rect 63221 2431 63279 2437
rect 63221 2428 63233 2431
rect 62592 2400 63233 2428
rect 62592 2304 62620 2400
rect 63221 2397 63233 2400
rect 63267 2397 63279 2431
rect 63221 2391 63279 2397
rect 63494 2388 63500 2440
rect 63552 2388 63558 2440
rect 66809 2431 66867 2437
rect 66809 2428 66821 2431
rect 66272 2400 66821 2428
rect 66272 2304 66300 2400
rect 66809 2397 66821 2400
rect 66855 2397 66867 2431
rect 66809 2391 66867 2397
rect 67085 2363 67143 2369
rect 67085 2329 67097 2363
rect 67131 2360 67143 2363
rect 70762 2360 70768 2372
rect 67131 2332 70768 2360
rect 67131 2329 67143 2332
rect 67085 2323 67143 2329
rect 70762 2320 70768 2332
rect 70820 2320 70826 2372
rect 70872 2360 70900 2468
rect 71593 2465 71605 2499
rect 71639 2496 71651 2499
rect 74534 2496 74540 2508
rect 71639 2468 74540 2496
rect 71639 2465 71651 2468
rect 71593 2459 71651 2465
rect 74534 2456 74540 2468
rect 74592 2456 74598 2508
rect 74994 2496 75000 2508
rect 74644 2468 75000 2496
rect 74644 2440 74672 2468
rect 74994 2456 75000 2468
rect 75052 2456 75058 2508
rect 110782 2496 110788 2508
rect 92216 2468 107424 2496
rect 71038 2388 71044 2440
rect 71096 2388 71102 2440
rect 74169 2431 74227 2437
rect 74169 2397 74181 2431
rect 74215 2428 74227 2431
rect 74626 2428 74632 2440
rect 74215 2400 74632 2428
rect 74215 2397 74227 2400
rect 74169 2391 74227 2397
rect 74626 2388 74632 2400
rect 74684 2388 74690 2440
rect 74718 2388 74724 2440
rect 74776 2388 74782 2440
rect 92014 2388 92020 2440
rect 92072 2388 92078 2440
rect 74736 2360 74764 2388
rect 70872 2332 74764 2360
rect 75270 2320 75276 2372
rect 75328 2320 75334 2372
rect 55916 2264 60734 2292
rect 55916 2252 55922 2264
rect 62574 2252 62580 2304
rect 62632 2252 62638 2304
rect 66254 2252 66260 2304
rect 66312 2252 66318 2304
rect 92216 2301 92244 2468
rect 92290 2388 92296 2440
rect 92348 2428 92354 2440
rect 92661 2431 92719 2437
rect 92661 2428 92673 2431
rect 92348 2400 92673 2428
rect 92348 2388 92354 2400
rect 92661 2397 92673 2400
rect 92707 2397 92719 2431
rect 92661 2391 92719 2397
rect 98089 2431 98147 2437
rect 98089 2397 98101 2431
rect 98135 2428 98147 2431
rect 98638 2428 98644 2440
rect 98135 2400 98644 2428
rect 98135 2397 98147 2400
rect 98089 2391 98147 2397
rect 98638 2388 98644 2400
rect 98696 2388 98702 2440
rect 103882 2388 103888 2440
rect 103940 2428 103946 2440
rect 107396 2437 107424 2468
rect 110248 2468 110788 2496
rect 104529 2431 104587 2437
rect 104529 2428 104541 2431
rect 103940 2400 104541 2428
rect 103940 2388 103946 2400
rect 104529 2397 104541 2400
rect 104575 2397 104587 2431
rect 104529 2391 104587 2397
rect 107381 2431 107439 2437
rect 107381 2397 107393 2431
rect 107427 2397 107439 2431
rect 107381 2391 107439 2397
rect 107654 2388 107660 2440
rect 107712 2388 107718 2440
rect 108390 2388 108396 2440
rect 108448 2388 108454 2440
rect 110248 2437 110276 2468
rect 110782 2456 110788 2468
rect 110840 2456 110846 2508
rect 113358 2456 113364 2508
rect 113416 2496 113422 2508
rect 113545 2499 113603 2505
rect 113545 2496 113557 2499
rect 113416 2468 113557 2496
rect 113416 2456 113422 2468
rect 113545 2465 113557 2468
rect 113591 2465 113603 2499
rect 113545 2459 113603 2465
rect 114922 2456 114928 2508
rect 114980 2456 114986 2508
rect 149348 2505 149376 2536
rect 242897 2533 242909 2536
rect 242943 2533 242955 2567
rect 301332 2564 301360 2604
rect 301406 2592 301412 2644
rect 301464 2632 301470 2644
rect 301501 2635 301559 2641
rect 301501 2632 301513 2635
rect 301464 2604 301513 2632
rect 301464 2592 301470 2604
rect 301501 2601 301513 2604
rect 301547 2601 301559 2635
rect 301501 2595 301559 2601
rect 302878 2592 302884 2644
rect 302936 2592 302942 2644
rect 304718 2592 304724 2644
rect 304776 2592 304782 2644
rect 308398 2592 308404 2644
rect 308456 2592 308462 2644
rect 308582 2592 308588 2644
rect 308640 2632 308646 2644
rect 308640 2604 314240 2632
rect 308640 2592 308646 2604
rect 302786 2564 302792 2576
rect 242897 2527 242955 2533
rect 249352 2536 301084 2564
rect 301332 2536 302792 2564
rect 116765 2499 116823 2505
rect 116765 2465 116777 2499
rect 116811 2496 116823 2499
rect 149333 2499 149391 2505
rect 116811 2468 142154 2496
rect 116811 2465 116823 2468
rect 116765 2459 116823 2465
rect 110233 2431 110291 2437
rect 110233 2397 110245 2431
rect 110279 2397 110291 2431
rect 110233 2391 110291 2397
rect 112346 2388 112352 2440
rect 112404 2388 112410 2440
rect 114097 2431 114155 2437
rect 114097 2397 114109 2431
rect 114143 2428 114155 2431
rect 114186 2428 114192 2440
rect 114143 2400 114192 2428
rect 114143 2397 114155 2400
rect 114097 2391 114155 2397
rect 114186 2388 114192 2400
rect 114244 2388 114250 2440
rect 116121 2431 116179 2437
rect 116121 2397 116133 2431
rect 116167 2428 116179 2431
rect 116210 2428 116216 2440
rect 116167 2400 116216 2428
rect 116167 2397 116179 2400
rect 116121 2391 116179 2397
rect 116210 2388 116216 2400
rect 116268 2428 116274 2440
rect 117866 2428 117872 2440
rect 116268 2400 117872 2428
rect 116268 2388 116274 2400
rect 117866 2388 117872 2400
rect 117924 2388 117930 2440
rect 118050 2388 118056 2440
rect 118108 2388 118114 2440
rect 119264 2437 119292 2468
rect 119249 2431 119307 2437
rect 119249 2397 119261 2431
rect 119295 2397 119307 2431
rect 119249 2391 119307 2397
rect 120626 2388 120632 2440
rect 120684 2388 120690 2440
rect 121825 2431 121883 2437
rect 121825 2397 121837 2431
rect 121871 2428 121883 2431
rect 122374 2428 122380 2440
rect 121871 2400 122380 2428
rect 121871 2397 121883 2400
rect 121825 2391 121883 2397
rect 122374 2388 122380 2400
rect 122432 2388 122438 2440
rect 123205 2431 123263 2437
rect 123205 2397 123217 2431
rect 123251 2428 123263 2431
rect 123478 2428 123484 2440
rect 123251 2400 123484 2428
rect 123251 2397 123263 2400
rect 123205 2391 123263 2397
rect 123478 2388 123484 2400
rect 123536 2388 123542 2440
rect 124401 2431 124459 2437
rect 124401 2397 124413 2431
rect 124447 2428 124459 2431
rect 124490 2428 124496 2440
rect 124447 2400 124496 2428
rect 124447 2397 124459 2400
rect 124401 2391 124459 2397
rect 124490 2388 124496 2400
rect 124548 2388 124554 2440
rect 125505 2431 125563 2437
rect 125505 2397 125517 2431
rect 125551 2397 125563 2431
rect 125505 2391 125563 2397
rect 96890 2320 96896 2372
rect 96948 2320 96954 2372
rect 105078 2320 105084 2372
rect 105136 2320 105142 2372
rect 108942 2320 108948 2372
rect 109000 2320 109006 2372
rect 112898 2320 112904 2372
rect 112956 2320 112962 2372
rect 117498 2320 117504 2372
rect 117556 2320 117562 2372
rect 118694 2320 118700 2372
rect 118752 2320 118758 2372
rect 120166 2320 120172 2372
rect 120224 2320 120230 2372
rect 121454 2320 121460 2372
rect 121512 2320 121518 2372
rect 122834 2320 122840 2372
rect 122892 2320 122898 2372
rect 123846 2320 123852 2372
rect 123904 2320 123910 2372
rect 125226 2320 125232 2372
rect 125284 2320 125290 2372
rect 125520 2360 125548 2391
rect 126054 2388 126060 2440
rect 126112 2388 126118 2440
rect 126606 2388 126612 2440
rect 126664 2388 126670 2440
rect 128265 2431 128323 2437
rect 128265 2397 128277 2431
rect 128311 2428 128323 2431
rect 130841 2431 130899 2437
rect 130841 2428 130853 2431
rect 128311 2400 128860 2428
rect 128311 2397 128323 2400
rect 128265 2391 128323 2397
rect 126422 2360 126428 2372
rect 125520 2332 126428 2360
rect 126422 2320 126428 2332
rect 126480 2320 126486 2372
rect 128832 2304 128860 2400
rect 130212 2400 130853 2428
rect 130212 2304 130240 2400
rect 130841 2397 130853 2400
rect 130887 2397 130899 2431
rect 130841 2391 130899 2397
rect 131390 2388 131396 2440
rect 131448 2388 131454 2440
rect 136729 2431 136787 2437
rect 136729 2428 136741 2431
rect 136100 2400 136741 2428
rect 136100 2304 136128 2400
rect 136729 2397 136741 2400
rect 136775 2397 136787 2431
rect 136729 2391 136787 2397
rect 137278 2388 137284 2440
rect 137336 2388 137342 2440
rect 142126 2360 142154 2468
rect 149333 2465 149345 2499
rect 149379 2465 149391 2499
rect 149333 2459 149391 2465
rect 151786 2468 211752 2496
rect 143166 2388 143172 2440
rect 143224 2428 143230 2440
rect 143353 2431 143411 2437
rect 143353 2428 143365 2431
rect 143224 2400 143365 2428
rect 143224 2388 143230 2400
rect 143353 2397 143365 2400
rect 143399 2397 143411 2431
rect 143353 2391 143411 2397
rect 143902 2388 143908 2440
rect 143960 2388 143966 2440
rect 145834 2388 145840 2440
rect 145892 2428 145898 2440
rect 146297 2431 146355 2437
rect 146297 2428 146309 2431
rect 145892 2400 146309 2428
rect 145892 2388 145898 2400
rect 146297 2397 146309 2400
rect 146343 2397 146355 2431
rect 146297 2391 146355 2397
rect 148226 2388 148232 2440
rect 148284 2428 148290 2440
rect 148873 2431 148931 2437
rect 148873 2428 148885 2431
rect 148284 2400 148885 2428
rect 148284 2388 148290 2400
rect 148873 2397 148885 2400
rect 148919 2397 148931 2431
rect 151786 2428 151814 2468
rect 148873 2391 148931 2397
rect 149532 2400 151814 2428
rect 149532 2360 149560 2400
rect 152182 2388 152188 2440
rect 152240 2388 152246 2440
rect 153473 2431 153531 2437
rect 153473 2428 153485 2431
rect 152752 2400 153485 2428
rect 142126 2332 149560 2360
rect 150986 2320 150992 2372
rect 151044 2320 151050 2372
rect 152752 2304 152780 2400
rect 153473 2397 153485 2400
rect 153519 2397 153531 2431
rect 153473 2391 153531 2397
rect 156690 2388 156696 2440
rect 156748 2428 156754 2440
rect 157337 2431 157395 2437
rect 157337 2428 157349 2431
rect 156748 2400 157349 2428
rect 156748 2388 156754 2400
rect 157337 2397 157349 2400
rect 157383 2397 157395 2431
rect 161293 2431 161351 2437
rect 161293 2428 161305 2431
rect 157337 2391 157395 2397
rect 160480 2400 161305 2428
rect 154022 2320 154028 2372
rect 154080 2320 154086 2372
rect 157886 2320 157892 2372
rect 157944 2320 157950 2372
rect 160480 2304 160508 2400
rect 161293 2397 161305 2400
rect 161339 2397 161351 2431
rect 161293 2391 161351 2397
rect 164326 2388 164332 2440
rect 164384 2388 164390 2440
rect 164786 2388 164792 2440
rect 164844 2428 164850 2440
rect 165065 2431 165123 2437
rect 165065 2428 165077 2431
rect 164844 2400 165077 2428
rect 164844 2388 164850 2400
rect 165065 2397 165077 2400
rect 165111 2397 165123 2431
rect 165065 2391 165123 2397
rect 170217 2431 170275 2437
rect 170217 2397 170229 2431
rect 170263 2397 170275 2431
rect 170217 2391 170275 2397
rect 182361 2431 182419 2437
rect 182361 2397 182373 2431
rect 182407 2428 182419 2431
rect 182407 2400 182956 2428
rect 182407 2397 182419 2400
rect 182361 2391 182419 2397
rect 161842 2320 161848 2372
rect 161900 2320 161906 2372
rect 165522 2320 165528 2372
rect 165580 2320 165586 2372
rect 169018 2320 169024 2372
rect 169076 2320 169082 2372
rect 92201 2295 92259 2301
rect 92201 2261 92213 2295
rect 92247 2261 92259 2295
rect 92201 2255 92259 2261
rect 110046 2252 110052 2304
rect 110104 2252 110110 2304
rect 126882 2252 126888 2304
rect 126940 2292 126946 2304
rect 128081 2295 128139 2301
rect 128081 2292 128093 2295
rect 126940 2264 128093 2292
rect 126940 2252 126946 2264
rect 128081 2261 128093 2264
rect 128127 2261 128139 2295
rect 128081 2255 128139 2261
rect 128814 2252 128820 2304
rect 128872 2252 128878 2304
rect 130194 2252 130200 2304
rect 130252 2252 130258 2304
rect 136082 2252 136088 2304
rect 136140 2252 136146 2304
rect 146110 2252 146116 2304
rect 146168 2252 146174 2304
rect 152734 2252 152740 2304
rect 152792 2252 152798 2304
rect 160462 2252 160468 2304
rect 160520 2252 160526 2304
rect 164142 2252 164148 2304
rect 164200 2252 164206 2304
rect 170232 2292 170260 2391
rect 182928 2304 182956 2400
rect 192202 2388 192208 2440
rect 192260 2388 192266 2440
rect 193033 2431 193091 2437
rect 193033 2397 193045 2431
rect 193079 2397 193091 2431
rect 198553 2431 198611 2437
rect 198553 2428 198565 2431
rect 193033 2391 193091 2397
rect 197924 2400 198565 2428
rect 170766 2292 170772 2304
rect 170232 2264 170772 2292
rect 170766 2252 170772 2264
rect 170824 2252 170830 2304
rect 182910 2252 182916 2304
rect 182968 2252 182974 2304
rect 193048 2292 193076 2391
rect 197924 2304 197952 2400
rect 198553 2397 198565 2400
rect 198599 2397 198611 2431
rect 198553 2391 198611 2397
rect 200206 2388 200212 2440
rect 200264 2428 200270 2440
rect 200853 2431 200911 2437
rect 200853 2428 200865 2431
rect 200264 2400 200865 2428
rect 200264 2388 200270 2400
rect 200853 2397 200865 2400
rect 200899 2397 200911 2431
rect 203337 2431 203395 2437
rect 203337 2428 203349 2431
rect 200853 2391 200911 2397
rect 202708 2400 203349 2428
rect 199105 2363 199163 2369
rect 199105 2329 199117 2363
rect 199151 2360 199163 2363
rect 199378 2360 199384 2372
rect 199151 2332 199384 2360
rect 199151 2329 199163 2332
rect 199105 2323 199163 2329
rect 199378 2320 199384 2332
rect 199436 2320 199442 2372
rect 202708 2304 202736 2400
rect 203337 2397 203349 2400
rect 203383 2397 203395 2431
rect 203337 2391 203395 2397
rect 203886 2388 203892 2440
rect 203944 2388 203950 2440
rect 205545 2431 205603 2437
rect 205545 2428 205557 2431
rect 204916 2400 205557 2428
rect 204916 2304 204944 2400
rect 205545 2397 205557 2400
rect 205591 2397 205603 2431
rect 205545 2391 205603 2397
rect 207658 2388 207664 2440
rect 207716 2388 207722 2440
rect 208213 2431 208271 2437
rect 208213 2397 208225 2431
rect 208259 2428 208271 2431
rect 208394 2428 208400 2440
rect 208259 2400 208400 2428
rect 208259 2397 208271 2400
rect 208213 2391 208271 2397
rect 208394 2388 208400 2400
rect 208452 2388 208458 2440
rect 209406 2428 209412 2440
rect 208688 2400 209412 2428
rect 206094 2320 206100 2372
rect 206152 2320 206158 2372
rect 206925 2363 206983 2369
rect 206925 2329 206937 2363
rect 206971 2360 206983 2363
rect 208688 2360 208716 2400
rect 209406 2388 209412 2400
rect 209464 2388 209470 2440
rect 211065 2431 211123 2437
rect 211065 2397 211077 2431
rect 211111 2397 211123 2431
rect 211065 2391 211123 2397
rect 206971 2332 208716 2360
rect 206971 2329 206983 2332
rect 206925 2323 206983 2329
rect 208854 2320 208860 2372
rect 208912 2320 208918 2372
rect 210234 2320 210240 2372
rect 210292 2320 210298 2372
rect 211080 2360 211108 2391
rect 211522 2388 211528 2440
rect 211580 2388 211586 2440
rect 211724 2428 211752 2468
rect 211798 2456 211804 2508
rect 211856 2456 211862 2508
rect 214926 2496 214932 2508
rect 211908 2468 214932 2496
rect 211908 2428 211936 2468
rect 214926 2456 214932 2468
rect 214984 2456 214990 2508
rect 216858 2496 216864 2508
rect 216692 2468 216864 2496
rect 216692 2440 216720 2468
rect 216858 2456 216864 2468
rect 216916 2456 216922 2508
rect 219158 2456 219164 2508
rect 219216 2456 219222 2508
rect 221642 2496 221648 2508
rect 219728 2468 221648 2496
rect 211724 2400 211936 2428
rect 213365 2431 213423 2437
rect 213365 2397 213377 2431
rect 213411 2428 213423 2431
rect 213638 2428 213644 2440
rect 213411 2400 213644 2428
rect 213411 2397 213423 2400
rect 213365 2391 213423 2397
rect 213638 2388 213644 2400
rect 213696 2388 213702 2440
rect 214282 2388 214288 2440
rect 214340 2428 214346 2440
rect 214561 2431 214619 2437
rect 214561 2428 214573 2431
rect 214340 2400 214573 2428
rect 214340 2388 214346 2400
rect 214561 2397 214573 2400
rect 214607 2397 214619 2431
rect 214561 2391 214619 2397
rect 215941 2431 215999 2437
rect 215941 2397 215953 2431
rect 215987 2428 215999 2431
rect 216674 2428 216680 2440
rect 215987 2400 216680 2428
rect 215987 2397 215999 2400
rect 215941 2391 215999 2397
rect 216674 2388 216680 2400
rect 216732 2388 216738 2440
rect 216766 2388 216772 2440
rect 216824 2428 216830 2440
rect 217137 2431 217195 2437
rect 217137 2428 217149 2431
rect 216824 2400 217149 2428
rect 216824 2388 216830 2400
rect 217137 2397 217149 2400
rect 217183 2428 217195 2431
rect 217183 2400 218376 2428
rect 217183 2397 217195 2400
rect 217137 2391 217195 2397
rect 211614 2360 211620 2372
rect 211080 2332 211620 2360
rect 211614 2320 211620 2332
rect 211672 2360 211678 2372
rect 212442 2360 212448 2372
rect 211672 2332 212448 2360
rect 211672 2320 211678 2332
rect 212442 2320 212448 2332
rect 212500 2320 212506 2372
rect 212810 2320 212816 2372
rect 212868 2320 212874 2372
rect 214006 2320 214012 2372
rect 214064 2320 214070 2372
rect 215386 2320 215392 2372
rect 215444 2320 215450 2372
rect 216582 2320 216588 2372
rect 216640 2320 216646 2372
rect 193582 2292 193588 2304
rect 193048 2264 193588 2292
rect 193582 2252 193588 2264
rect 193640 2252 193646 2304
rect 197906 2252 197912 2304
rect 197964 2252 197970 2304
rect 200390 2252 200396 2304
rect 200448 2252 200454 2304
rect 202690 2252 202696 2304
rect 202748 2252 202754 2304
rect 204898 2252 204904 2304
rect 204956 2252 204962 2304
rect 217962 2252 217968 2304
rect 218020 2292 218026 2304
rect 218241 2295 218299 2301
rect 218241 2292 218253 2295
rect 218020 2264 218253 2292
rect 218020 2252 218026 2264
rect 218241 2261 218253 2264
rect 218287 2261 218299 2295
rect 218348 2292 218376 2400
rect 218422 2388 218428 2440
rect 218480 2388 218486 2440
rect 219728 2437 219756 2468
rect 221642 2456 221648 2468
rect 221700 2496 221706 2508
rect 221700 2468 238754 2496
rect 221700 2456 221706 2468
rect 219713 2431 219771 2437
rect 219713 2397 219725 2431
rect 219759 2397 219771 2431
rect 219713 2391 219771 2397
rect 220354 2388 220360 2440
rect 220412 2428 220418 2440
rect 220449 2431 220507 2437
rect 220449 2428 220461 2431
rect 220412 2400 220461 2428
rect 220412 2388 220418 2400
rect 220449 2397 220461 2400
rect 220495 2397 220507 2431
rect 220449 2391 220507 2397
rect 220464 2360 220492 2391
rect 220998 2388 221004 2440
rect 221056 2388 221062 2440
rect 223577 2431 223635 2437
rect 223577 2397 223589 2431
rect 223623 2428 223635 2431
rect 223623 2400 224264 2428
rect 223623 2397 223635 2400
rect 223577 2391 223635 2397
rect 221553 2363 221611 2369
rect 221553 2360 221565 2363
rect 220464 2332 221565 2360
rect 221553 2329 221565 2332
rect 221599 2329 221611 2363
rect 221553 2323 221611 2329
rect 223022 2320 223028 2372
rect 223080 2320 223086 2372
rect 224236 2304 224264 2400
rect 224954 2388 224960 2440
rect 225012 2428 225018 2440
rect 225601 2431 225659 2437
rect 225601 2428 225613 2431
rect 225012 2400 225613 2428
rect 225012 2388 225018 2400
rect 225601 2397 225613 2400
rect 225647 2397 225659 2431
rect 225601 2391 225659 2397
rect 230750 2388 230756 2440
rect 230808 2428 230814 2440
rect 231397 2431 231455 2437
rect 231397 2428 231409 2431
rect 230808 2400 231409 2428
rect 230808 2388 230814 2400
rect 231397 2397 231409 2400
rect 231443 2397 231455 2431
rect 231397 2391 231455 2397
rect 236457 2431 236515 2437
rect 236457 2397 236469 2431
rect 236503 2428 236515 2431
rect 236503 2400 237052 2428
rect 236503 2397 236515 2400
rect 236457 2391 236515 2397
rect 226150 2320 226156 2372
rect 226208 2320 226214 2372
rect 231946 2320 231952 2372
rect 232004 2320 232010 2372
rect 237024 2304 237052 2400
rect 237742 2388 237748 2440
rect 237800 2428 237806 2440
rect 238481 2431 238539 2437
rect 238481 2428 238493 2431
rect 237800 2400 238493 2428
rect 237800 2388 237806 2400
rect 238481 2397 238493 2400
rect 238527 2397 238539 2431
rect 238481 2391 238539 2397
rect 238726 2360 238754 2468
rect 239030 2388 239036 2440
rect 239088 2388 239094 2440
rect 242912 2428 242940 2527
rect 243740 2468 249288 2496
rect 243633 2431 243691 2437
rect 243633 2428 243645 2431
rect 242912 2400 243645 2428
rect 243633 2397 243645 2400
rect 243679 2397 243691 2431
rect 243633 2391 243691 2397
rect 243740 2360 243768 2468
rect 247126 2388 247132 2440
rect 247184 2388 247190 2440
rect 248785 2431 248843 2437
rect 248785 2428 248797 2431
rect 248386 2400 248797 2428
rect 238726 2332 243768 2360
rect 244182 2320 244188 2372
rect 244240 2320 244246 2372
rect 246298 2320 246304 2372
rect 246356 2320 246362 2372
rect 221366 2292 221372 2304
rect 218348 2264 221372 2292
rect 218241 2255 218299 2261
rect 221366 2252 221372 2264
rect 221424 2252 221430 2304
rect 224218 2252 224224 2304
rect 224276 2252 224282 2304
rect 236270 2252 236276 2304
rect 236328 2252 236334 2304
rect 237006 2252 237012 2304
rect 237064 2252 237070 2304
rect 248046 2252 248052 2304
rect 248104 2292 248110 2304
rect 248386 2292 248414 2400
rect 248785 2397 248797 2400
rect 248831 2397 248843 2431
rect 248785 2391 248843 2397
rect 249260 2360 249288 2468
rect 249352 2437 249380 2536
rect 291102 2496 291108 2508
rect 249444 2468 289860 2496
rect 249337 2431 249395 2437
rect 249337 2397 249349 2431
rect 249383 2397 249395 2431
rect 249337 2391 249395 2397
rect 249444 2360 249472 2468
rect 251726 2388 251732 2440
rect 251784 2388 251790 2440
rect 254026 2388 254032 2440
rect 254084 2428 254090 2440
rect 254489 2431 254547 2437
rect 254489 2428 254501 2431
rect 254084 2400 254501 2428
rect 254084 2388 254090 2400
rect 254489 2397 254501 2400
rect 254535 2397 254547 2431
rect 254489 2391 254547 2397
rect 255774 2388 255780 2440
rect 255832 2428 255838 2440
rect 256513 2431 256571 2437
rect 256513 2428 256525 2431
rect 255832 2400 256525 2428
rect 255832 2388 255838 2400
rect 256513 2397 256525 2400
rect 256559 2397 256571 2431
rect 259457 2431 259515 2437
rect 259457 2428 259469 2431
rect 256513 2391 256571 2397
rect 258368 2400 259469 2428
rect 249260 2332 249472 2360
rect 252281 2363 252339 2369
rect 252281 2329 252293 2363
rect 252327 2360 252339 2363
rect 252327 2332 255912 2360
rect 252327 2329 252339 2332
rect 252281 2323 252339 2329
rect 248104 2264 248414 2292
rect 248104 2252 248110 2264
rect 254302 2252 254308 2304
rect 254360 2252 254366 2304
rect 255774 2252 255780 2304
rect 255832 2252 255838 2304
rect 255884 2292 255912 2332
rect 257062 2320 257068 2372
rect 257120 2320 257126 2372
rect 258368 2304 258396 2400
rect 259457 2397 259469 2400
rect 259503 2397 259515 2431
rect 259457 2391 259515 2397
rect 260006 2388 260012 2440
rect 260064 2388 260070 2440
rect 262306 2388 262312 2440
rect 262364 2428 262370 2440
rect 262953 2431 263011 2437
rect 262953 2428 262965 2431
rect 262364 2400 262965 2428
rect 262364 2388 262370 2400
rect 262953 2397 262965 2400
rect 262999 2397 263011 2431
rect 262953 2391 263011 2397
rect 263502 2388 263508 2440
rect 263560 2388 263566 2440
rect 265161 2431 265219 2437
rect 265161 2397 265173 2431
rect 265207 2397 265219 2431
rect 265161 2391 265219 2397
rect 272521 2431 272579 2437
rect 272521 2397 272533 2431
rect 272567 2428 272579 2431
rect 273070 2428 273076 2440
rect 272567 2400 273076 2428
rect 272567 2397 272579 2400
rect 272521 2391 272579 2397
rect 264330 2320 264336 2372
rect 264388 2320 264394 2372
rect 258258 2292 258264 2304
rect 255884 2264 258264 2292
rect 258258 2252 258264 2264
rect 258316 2252 258322 2304
rect 258350 2252 258356 2304
rect 258408 2252 258414 2304
rect 265176 2292 265204 2391
rect 273070 2388 273076 2400
rect 273128 2388 273134 2440
rect 277673 2431 277731 2437
rect 277673 2397 277685 2431
rect 277719 2428 277731 2431
rect 286505 2431 286563 2437
rect 277719 2400 278360 2428
rect 277719 2397 277731 2400
rect 277673 2391 277731 2397
rect 277118 2320 277124 2372
rect 277176 2320 277182 2372
rect 278332 2304 278360 2400
rect 286505 2397 286517 2431
rect 286551 2428 286563 2431
rect 287422 2428 287428 2440
rect 286551 2400 287428 2428
rect 286551 2397 286563 2400
rect 286505 2391 286563 2397
rect 287422 2388 287428 2400
rect 287480 2388 287486 2440
rect 285950 2320 285956 2372
rect 286008 2320 286014 2372
rect 289832 2360 289860 2468
rect 290568 2468 291108 2496
rect 290568 2437 290596 2468
rect 291102 2456 291108 2468
rect 291160 2456 291166 2508
rect 293770 2456 293776 2508
rect 293828 2456 293834 2508
rect 297729 2499 297787 2505
rect 297729 2496 297741 2499
rect 293880 2468 297741 2496
rect 290553 2431 290611 2437
rect 290553 2397 290565 2431
rect 290599 2397 290611 2431
rect 290553 2391 290611 2397
rect 292574 2388 292580 2440
rect 292632 2428 292638 2440
rect 293221 2431 293279 2437
rect 293221 2428 293233 2431
rect 292632 2400 293233 2428
rect 292632 2388 292638 2400
rect 293221 2397 293233 2400
rect 293267 2397 293279 2431
rect 293221 2391 293279 2397
rect 293880 2360 293908 2468
rect 297729 2465 297741 2468
rect 297775 2465 297787 2499
rect 297729 2459 297787 2465
rect 295426 2388 295432 2440
rect 295484 2388 295490 2440
rect 296441 2431 296499 2437
rect 296441 2397 296453 2431
rect 296487 2428 296499 2431
rect 296530 2428 296536 2440
rect 296487 2400 296536 2428
rect 296487 2397 296499 2400
rect 296441 2391 296499 2397
rect 296530 2388 296536 2400
rect 296588 2388 296594 2440
rect 296990 2388 296996 2440
rect 297048 2388 297054 2440
rect 298005 2431 298063 2437
rect 298005 2397 298017 2431
rect 298051 2428 298063 2431
rect 298646 2428 298652 2440
rect 298051 2400 298652 2428
rect 298051 2397 298063 2400
rect 298005 2391 298063 2397
rect 298646 2388 298652 2400
rect 298704 2388 298710 2440
rect 299566 2388 299572 2440
rect 299624 2388 299630 2440
rect 300302 2388 300308 2440
rect 300360 2388 300366 2440
rect 289832 2332 293908 2360
rect 295794 2320 295800 2372
rect 295852 2320 295858 2372
rect 299014 2320 299020 2372
rect 299072 2320 299078 2372
rect 300762 2320 300768 2372
rect 300820 2320 300826 2372
rect 301056 2360 301084 2536
rect 302786 2524 302792 2536
rect 302844 2524 302850 2576
rect 302896 2496 302924 2592
rect 309042 2564 309048 2576
rect 302206 2468 302924 2496
rect 303908 2536 309048 2564
rect 301777 2431 301835 2437
rect 301777 2397 301789 2431
rect 301823 2428 301835 2431
rect 302206 2428 302234 2468
rect 301823 2400 302234 2428
rect 301823 2397 301835 2400
rect 301777 2391 301835 2397
rect 302786 2388 302792 2440
rect 302844 2428 302850 2440
rect 303433 2431 303491 2437
rect 303433 2428 303445 2431
rect 302844 2400 303445 2428
rect 302844 2388 302850 2400
rect 303433 2397 303445 2400
rect 303479 2397 303491 2431
rect 303433 2391 303491 2397
rect 303908 2360 303936 2536
rect 309042 2524 309048 2536
rect 309100 2524 309106 2576
rect 312262 2564 312268 2576
rect 310992 2536 312268 2564
rect 305454 2456 305460 2508
rect 305512 2496 305518 2508
rect 310882 2496 310888 2508
rect 305512 2468 310888 2496
rect 305512 2456 305518 2468
rect 310882 2456 310888 2468
rect 310940 2456 310946 2508
rect 304166 2388 304172 2440
rect 304224 2428 304230 2440
rect 304537 2431 304595 2437
rect 304537 2428 304549 2431
rect 304224 2400 304549 2428
rect 304224 2388 304230 2400
rect 304537 2397 304549 2400
rect 304583 2397 304595 2431
rect 304537 2391 304595 2397
rect 306006 2388 306012 2440
rect 306064 2388 306070 2440
rect 306742 2388 306748 2440
rect 306800 2388 306806 2440
rect 309505 2431 309563 2437
rect 309505 2397 309517 2431
rect 309551 2428 309563 2431
rect 310606 2428 310612 2440
rect 309551 2400 310612 2428
rect 309551 2397 309563 2400
rect 309505 2391 309563 2397
rect 310606 2388 310612 2400
rect 310664 2388 310670 2440
rect 310698 2388 310704 2440
rect 310756 2388 310762 2440
rect 310992 2437 311020 2536
rect 312262 2524 312268 2536
rect 312320 2564 312326 2576
rect 313182 2564 313188 2576
rect 312320 2536 313188 2564
rect 312320 2524 312326 2536
rect 313182 2524 313188 2536
rect 313240 2524 313246 2576
rect 314212 2564 314240 2604
rect 314286 2592 314292 2644
rect 314344 2632 314350 2644
rect 314381 2635 314439 2641
rect 314381 2632 314393 2635
rect 314344 2604 314393 2632
rect 314344 2592 314350 2604
rect 314381 2601 314393 2604
rect 314427 2601 314439 2635
rect 314381 2595 314439 2601
rect 318334 2592 318340 2644
rect 318392 2592 318398 2644
rect 319622 2592 319628 2644
rect 319680 2592 319686 2644
rect 319714 2592 319720 2644
rect 319772 2632 319778 2644
rect 348329 2635 348387 2641
rect 348329 2632 348341 2635
rect 319772 2604 348341 2632
rect 319772 2592 319778 2604
rect 348329 2601 348341 2604
rect 348375 2601 348387 2635
rect 348329 2595 348387 2601
rect 350442 2592 350448 2644
rect 350500 2592 350506 2644
rect 355134 2592 355140 2644
rect 355192 2592 355198 2644
rect 355778 2592 355784 2644
rect 355836 2632 355842 2644
rect 355873 2635 355931 2641
rect 355873 2632 355885 2635
rect 355836 2604 355885 2632
rect 355836 2592 355842 2604
rect 355873 2601 355885 2604
rect 355919 2601 355931 2635
rect 355873 2595 355931 2601
rect 359550 2592 359556 2644
rect 359608 2592 359614 2644
rect 362494 2592 362500 2644
rect 362552 2592 362558 2644
rect 380526 2592 380532 2644
rect 380584 2592 380590 2644
rect 382734 2592 382740 2644
rect 382792 2592 382798 2644
rect 387150 2592 387156 2644
rect 387208 2592 387214 2644
rect 395614 2592 395620 2644
rect 395672 2592 395678 2644
rect 398558 2592 398564 2644
rect 398616 2592 398622 2644
rect 407850 2632 407856 2644
rect 398806 2604 407856 2632
rect 325234 2564 325240 2576
rect 314212 2536 325240 2564
rect 325234 2524 325240 2536
rect 325292 2524 325298 2576
rect 325326 2524 325332 2576
rect 325384 2524 325390 2576
rect 325418 2524 325424 2576
rect 325476 2564 325482 2576
rect 341429 2567 341487 2573
rect 341429 2564 341441 2567
rect 325476 2536 341441 2564
rect 325476 2524 325482 2536
rect 341429 2533 341441 2536
rect 341475 2533 341487 2567
rect 341429 2527 341487 2533
rect 342070 2524 342076 2576
rect 342128 2564 342134 2576
rect 398806 2564 398834 2604
rect 407850 2592 407856 2604
rect 407908 2592 407914 2644
rect 408494 2592 408500 2644
rect 408552 2632 408558 2644
rect 492674 2632 492680 2644
rect 408552 2604 492680 2632
rect 408552 2592 408558 2604
rect 492674 2592 492680 2604
rect 492732 2592 492738 2644
rect 342128 2536 398834 2564
rect 403636 2536 412634 2564
rect 342128 2524 342134 2536
rect 311158 2456 311164 2508
rect 311216 2496 311222 2508
rect 311216 2468 325280 2496
rect 311216 2456 311222 2468
rect 310977 2431 311035 2437
rect 310977 2397 310989 2431
rect 311023 2397 311035 2431
rect 312357 2431 312415 2437
rect 312357 2428 312369 2431
rect 310977 2391 311035 2397
rect 311176 2400 312369 2428
rect 301056 2332 303936 2360
rect 303982 2320 303988 2372
rect 304040 2320 304046 2372
rect 305454 2320 305460 2372
rect 305512 2320 305518 2372
rect 307294 2320 307300 2372
rect 307352 2320 307358 2372
rect 308493 2363 308551 2369
rect 308493 2329 308505 2363
rect 308539 2329 308551 2363
rect 308493 2323 308551 2329
rect 265710 2292 265716 2304
rect 265176 2264 265716 2292
rect 265710 2252 265716 2264
rect 265768 2252 265774 2304
rect 271782 2252 271788 2304
rect 271840 2292 271846 2304
rect 272337 2295 272395 2301
rect 272337 2292 272349 2295
rect 271840 2264 272349 2292
rect 271840 2252 271846 2264
rect 272337 2261 272349 2264
rect 272383 2261 272395 2295
rect 272337 2255 272395 2261
rect 278314 2252 278320 2304
rect 278372 2252 278378 2304
rect 288342 2252 288348 2304
rect 288400 2292 288406 2304
rect 290369 2295 290427 2301
rect 290369 2292 290381 2295
rect 288400 2264 290381 2292
rect 288400 2252 288406 2264
rect 290369 2261 290381 2264
rect 290415 2261 290427 2295
rect 290369 2255 290427 2261
rect 292574 2252 292580 2304
rect 292632 2252 292638 2304
rect 304994 2252 305000 2304
rect 305052 2292 305058 2304
rect 308508 2292 308536 2323
rect 309226 2320 309232 2372
rect 309284 2320 309290 2372
rect 311176 2360 311204 2400
rect 312357 2397 312369 2400
rect 312403 2397 312415 2431
rect 312357 2391 312415 2397
rect 313737 2431 313795 2437
rect 313737 2397 313749 2431
rect 313783 2428 313795 2431
rect 315669 2431 315727 2437
rect 315669 2428 315681 2431
rect 313783 2400 315681 2428
rect 313783 2397 313795 2400
rect 313737 2391 313795 2397
rect 315669 2397 315681 2400
rect 315715 2428 315727 2431
rect 315942 2428 315948 2440
rect 315715 2400 315948 2428
rect 315715 2397 315727 2400
rect 315669 2391 315727 2397
rect 315942 2388 315948 2400
rect 316000 2388 316006 2440
rect 316586 2388 316592 2440
rect 316644 2428 316650 2440
rect 317601 2431 317659 2437
rect 316644 2400 317184 2428
rect 316644 2388 316650 2400
rect 310532 2332 311204 2360
rect 311805 2363 311863 2369
rect 310532 2292 310560 2332
rect 311805 2329 311817 2363
rect 311851 2329 311863 2363
rect 311805 2323 311863 2329
rect 305052 2264 310560 2292
rect 305052 2252 305058 2264
rect 310606 2252 310612 2304
rect 310664 2292 310670 2304
rect 311342 2292 311348 2304
rect 310664 2264 311348 2292
rect 310664 2252 310670 2264
rect 311342 2252 311348 2264
rect 311400 2252 311406 2304
rect 311526 2252 311532 2304
rect 311584 2252 311590 2304
rect 311820 2292 311848 2323
rect 313274 2320 313280 2372
rect 313332 2320 313338 2372
rect 314657 2363 314715 2369
rect 314657 2329 314669 2363
rect 314703 2360 314715 2363
rect 315758 2360 315764 2372
rect 314703 2332 315764 2360
rect 314703 2329 314715 2332
rect 314657 2323 314715 2329
rect 315758 2320 315764 2332
rect 315816 2320 315822 2372
rect 317046 2320 317052 2372
rect 317104 2320 317110 2372
rect 317156 2360 317184 2400
rect 317601 2397 317613 2431
rect 317647 2428 317659 2431
rect 318334 2428 318340 2440
rect 317647 2400 318340 2428
rect 317647 2397 317659 2400
rect 317601 2391 317659 2397
rect 318334 2388 318340 2400
rect 318392 2388 318398 2440
rect 318978 2388 318984 2440
rect 319036 2388 319042 2440
rect 319438 2388 319444 2440
rect 319496 2388 319502 2440
rect 323581 2431 323639 2437
rect 323581 2397 323593 2431
rect 323627 2397 323639 2431
rect 323581 2391 323639 2397
rect 319714 2360 319720 2372
rect 317156 2332 319720 2360
rect 319714 2320 319720 2332
rect 319772 2320 319778 2372
rect 313366 2292 313372 2304
rect 311820 2264 313372 2292
rect 313366 2252 313372 2264
rect 313424 2252 313430 2304
rect 314746 2252 314752 2304
rect 314804 2292 314810 2304
rect 318797 2295 318855 2301
rect 318797 2292 318809 2295
rect 314804 2264 318809 2292
rect 314804 2252 314810 2264
rect 318797 2261 318809 2264
rect 318843 2261 318855 2295
rect 318797 2255 318855 2261
rect 323394 2252 323400 2304
rect 323452 2252 323458 2304
rect 323596 2292 323624 2391
rect 324682 2388 324688 2440
rect 324740 2388 324746 2440
rect 325142 2388 325148 2440
rect 325200 2388 325206 2440
rect 325252 2428 325280 2468
rect 325436 2468 357112 2496
rect 325252 2424 325372 2428
rect 325436 2424 325464 2468
rect 325252 2400 325464 2424
rect 325344 2396 325464 2400
rect 326617 2431 326675 2437
rect 326617 2397 326629 2431
rect 326663 2428 326675 2431
rect 327166 2428 327172 2440
rect 326663 2400 327172 2428
rect 326663 2397 326675 2400
rect 326617 2391 326675 2397
rect 327166 2388 327172 2400
rect 327224 2388 327230 2440
rect 329377 2431 329435 2437
rect 329377 2397 329389 2431
rect 329423 2428 329435 2431
rect 330018 2428 330024 2440
rect 329423 2400 330024 2428
rect 329423 2397 329435 2400
rect 329377 2391 329435 2397
rect 330018 2388 330024 2400
rect 330076 2388 330082 2440
rect 331769 2431 331827 2437
rect 331769 2397 331781 2431
rect 331815 2397 331827 2431
rect 331769 2391 331827 2397
rect 331214 2320 331220 2372
rect 331272 2320 331278 2372
rect 331784 2360 331812 2391
rect 332318 2388 332324 2440
rect 332376 2428 332382 2440
rect 333057 2431 333115 2437
rect 333057 2428 333069 2431
rect 332376 2400 333069 2428
rect 332376 2388 332382 2400
rect 333057 2397 333069 2400
rect 333103 2397 333115 2431
rect 333057 2391 333115 2397
rect 335449 2431 335507 2437
rect 335449 2397 335461 2431
rect 335495 2428 335507 2431
rect 336366 2428 336372 2440
rect 335495 2400 336372 2428
rect 335495 2397 335507 2400
rect 335449 2391 335507 2397
rect 336366 2388 336372 2400
rect 336424 2388 336430 2440
rect 337838 2388 337844 2440
rect 337896 2388 337902 2440
rect 340509 2431 340567 2437
rect 340509 2397 340521 2431
rect 340555 2428 340567 2431
rect 341518 2428 341524 2440
rect 340555 2400 341524 2428
rect 340555 2397 340567 2400
rect 340509 2391 340567 2397
rect 341518 2388 341524 2400
rect 341576 2388 341582 2440
rect 341613 2431 341671 2437
rect 341613 2397 341625 2431
rect 341659 2428 341671 2431
rect 342070 2428 342076 2440
rect 341659 2400 342076 2428
rect 341659 2397 341671 2400
rect 341613 2391 341671 2397
rect 342070 2388 342076 2400
rect 342128 2388 342134 2440
rect 342162 2388 342168 2440
rect 342220 2428 342226 2440
rect 342901 2431 342959 2437
rect 342901 2428 342913 2431
rect 342220 2400 342913 2428
rect 342220 2388 342226 2400
rect 342901 2397 342913 2400
rect 342947 2397 342959 2431
rect 342901 2391 342959 2397
rect 344649 2431 344707 2437
rect 344649 2397 344661 2431
rect 344695 2428 344707 2431
rect 345566 2428 345572 2440
rect 344695 2400 345572 2428
rect 344695 2397 344707 2400
rect 344649 2391 344707 2397
rect 345566 2388 345572 2400
rect 345624 2428 345630 2440
rect 346210 2428 346216 2440
rect 345624 2400 346216 2428
rect 345624 2388 345630 2400
rect 346210 2388 346216 2400
rect 346268 2388 346274 2440
rect 346578 2388 346584 2440
rect 346636 2428 346642 2440
rect 347317 2431 347375 2437
rect 347317 2428 347329 2431
rect 346636 2400 347329 2428
rect 346636 2388 346642 2400
rect 347317 2397 347329 2400
rect 347363 2397 347375 2431
rect 347317 2391 347375 2397
rect 350261 2431 350319 2437
rect 350261 2397 350273 2431
rect 350307 2428 350319 2431
rect 350626 2428 350632 2440
rect 350307 2400 350632 2428
rect 350307 2397 350319 2400
rect 350261 2391 350319 2397
rect 350626 2388 350632 2400
rect 350684 2388 350690 2440
rect 353662 2388 353668 2440
rect 353720 2388 353726 2440
rect 356054 2388 356060 2440
rect 356112 2388 356118 2440
rect 332778 2360 332784 2372
rect 331784 2332 332784 2360
rect 332778 2320 332784 2332
rect 332836 2320 332842 2372
rect 335262 2320 335268 2372
rect 335320 2320 335326 2372
rect 337286 2320 337292 2372
rect 337344 2320 337350 2372
rect 339954 2320 339960 2372
rect 340012 2320 340018 2372
rect 341978 2320 341984 2372
rect 342036 2360 342042 2372
rect 345753 2363 345811 2369
rect 342036 2332 344508 2360
rect 342036 2320 342042 2332
rect 323762 2292 323768 2304
rect 323596 2264 323768 2292
rect 323762 2252 323768 2264
rect 323820 2252 323826 2304
rect 324498 2252 324504 2304
rect 324556 2252 324562 2304
rect 326430 2252 326436 2304
rect 326488 2252 326494 2304
rect 329282 2252 329288 2304
rect 329340 2252 329346 2304
rect 332502 2252 332508 2304
rect 332560 2252 332566 2304
rect 337194 2252 337200 2304
rect 337252 2252 337258 2304
rect 338022 2252 338028 2304
rect 338080 2252 338086 2304
rect 342346 2252 342352 2304
rect 342404 2252 342410 2304
rect 344480 2301 344508 2332
rect 345753 2329 345765 2363
rect 345799 2360 345811 2363
rect 346670 2360 346676 2372
rect 345799 2332 346676 2360
rect 345799 2329 345811 2332
rect 345753 2323 345811 2329
rect 346670 2320 346676 2332
rect 346728 2320 346734 2372
rect 348418 2320 348424 2372
rect 348476 2320 348482 2372
rect 349706 2320 349712 2372
rect 349764 2320 349770 2372
rect 352374 2320 352380 2372
rect 352432 2320 352438 2372
rect 353294 2320 353300 2372
rect 353352 2320 353358 2372
rect 354493 2363 354551 2369
rect 354493 2329 354505 2363
rect 354539 2360 354551 2363
rect 355134 2360 355140 2372
rect 354539 2332 355140 2360
rect 354539 2329 354551 2332
rect 354493 2323 354551 2329
rect 355134 2320 355140 2332
rect 355192 2320 355198 2372
rect 344465 2295 344523 2301
rect 344465 2261 344477 2295
rect 344511 2261 344523 2295
rect 344465 2255 344523 2261
rect 345658 2252 345664 2304
rect 345716 2252 345722 2304
rect 346762 2252 346768 2304
rect 346820 2252 346826 2304
rect 349614 2252 349620 2304
rect 349672 2252 349678 2304
rect 352282 2252 352288 2304
rect 352340 2252 352346 2304
rect 354398 2252 354404 2304
rect 354456 2252 354462 2304
rect 357084 2301 357112 2468
rect 367278 2456 367284 2508
rect 367336 2456 367342 2508
rect 368477 2499 368535 2505
rect 368477 2496 368489 2499
rect 367848 2468 368489 2496
rect 357253 2431 357311 2437
rect 357253 2397 357265 2431
rect 357299 2428 357311 2431
rect 358170 2428 358176 2440
rect 357299 2400 358176 2428
rect 357299 2397 357311 2400
rect 357253 2391 357311 2397
rect 358170 2388 358176 2400
rect 358228 2388 358234 2440
rect 358449 2431 358507 2437
rect 358449 2397 358461 2431
rect 358495 2428 358507 2431
rect 359550 2428 359556 2440
rect 358495 2400 359556 2428
rect 358495 2397 358507 2400
rect 358449 2391 358507 2397
rect 359550 2388 359556 2400
rect 359608 2388 359614 2440
rect 362218 2388 362224 2440
rect 362276 2428 362282 2440
rect 367848 2437 367876 2468
rect 368477 2465 368489 2468
rect 368523 2496 368535 2499
rect 368523 2468 383654 2496
rect 368523 2465 368535 2468
rect 368477 2459 368535 2465
rect 362589 2431 362647 2437
rect 362589 2428 362601 2431
rect 362276 2400 362601 2428
rect 362276 2388 362282 2400
rect 362589 2397 362601 2400
rect 362635 2397 362647 2431
rect 362589 2391 362647 2397
rect 367833 2431 367891 2437
rect 367833 2397 367845 2431
rect 367879 2397 367891 2431
rect 367833 2391 367891 2397
rect 371697 2431 371755 2437
rect 371697 2397 371709 2431
rect 371743 2397 371755 2431
rect 371697 2391 371755 2397
rect 380713 2431 380771 2437
rect 380713 2397 380725 2431
rect 380759 2428 380771 2431
rect 380894 2428 380900 2440
rect 380759 2400 380900 2428
rect 380759 2397 380771 2400
rect 380713 2391 380771 2397
rect 357894 2320 357900 2372
rect 357952 2320 357958 2372
rect 371142 2320 371148 2372
rect 371200 2320 371206 2372
rect 371712 2360 371740 2391
rect 380894 2388 380900 2400
rect 380952 2388 380958 2440
rect 381262 2388 381268 2440
rect 381320 2388 381326 2440
rect 381817 2431 381875 2437
rect 381817 2397 381829 2431
rect 381863 2428 381875 2431
rect 382734 2428 382740 2440
rect 381863 2400 382740 2428
rect 381863 2397 381875 2400
rect 381817 2391 381875 2397
rect 382734 2388 382740 2400
rect 382792 2388 382798 2440
rect 383626 2428 383654 2468
rect 385310 2456 385316 2508
rect 385368 2456 385374 2508
rect 403636 2496 403664 2536
rect 385788 2468 403664 2496
rect 385788 2428 385816 2468
rect 403986 2456 403992 2508
rect 404044 2496 404050 2508
rect 404044 2468 404676 2496
rect 404044 2456 404050 2468
rect 383626 2400 385816 2428
rect 385865 2431 385923 2437
rect 385865 2397 385877 2431
rect 385911 2428 385923 2431
rect 385911 2400 386552 2428
rect 385911 2397 385923 2400
rect 385865 2391 385923 2397
rect 372430 2360 372436 2372
rect 371712 2332 372436 2360
rect 372430 2320 372436 2332
rect 372488 2320 372494 2372
rect 386524 2304 386552 2400
rect 387150 2388 387156 2440
rect 387208 2428 387214 2440
rect 387889 2431 387947 2437
rect 387889 2428 387901 2431
rect 387208 2400 387901 2428
rect 387208 2388 387214 2400
rect 387889 2397 387901 2400
rect 387935 2397 387947 2431
rect 387889 2391 387947 2397
rect 388438 2388 388444 2440
rect 388496 2388 388502 2440
rect 389545 2431 389603 2437
rect 389545 2397 389557 2431
rect 389591 2428 389603 2431
rect 389591 2400 390508 2428
rect 389591 2397 389603 2400
rect 389545 2391 389603 2397
rect 389266 2320 389272 2372
rect 389324 2320 389330 2372
rect 390480 2304 390508 2400
rect 391106 2388 391112 2440
rect 391164 2388 391170 2440
rect 394421 2431 394479 2437
rect 394421 2397 394433 2431
rect 394467 2428 394479 2431
rect 394694 2428 394700 2440
rect 394467 2400 394700 2428
rect 394467 2397 394479 2400
rect 394421 2391 394479 2397
rect 394694 2388 394700 2400
rect 394752 2388 394758 2440
rect 396902 2388 396908 2440
rect 396960 2388 396966 2440
rect 397362 2388 397368 2440
rect 397420 2388 397426 2440
rect 398745 2431 398803 2437
rect 398745 2397 398757 2431
rect 398791 2428 398803 2431
rect 398926 2428 398932 2440
rect 398791 2400 398932 2428
rect 398791 2397 398803 2400
rect 398745 2391 398803 2397
rect 398926 2388 398932 2400
rect 398984 2428 398990 2440
rect 398984 2400 399800 2428
rect 398984 2388 398990 2400
rect 391658 2320 391664 2372
rect 391716 2320 391722 2372
rect 393866 2320 393872 2372
rect 393924 2320 393930 2372
rect 395893 2363 395951 2369
rect 395893 2329 395905 2363
rect 395939 2360 395951 2363
rect 396166 2360 396172 2372
rect 395939 2332 396172 2360
rect 395939 2329 395951 2332
rect 395893 2323 395951 2329
rect 396166 2320 396172 2332
rect 396224 2360 396230 2372
rect 396224 2332 398696 2360
rect 396224 2320 396230 2332
rect 357069 2295 357127 2301
rect 357069 2261 357081 2295
rect 357115 2261 357127 2295
rect 357069 2255 357127 2261
rect 386506 2252 386512 2304
rect 386564 2252 386570 2304
rect 390462 2252 390468 2304
rect 390520 2252 390526 2304
rect 398668 2292 398696 2332
rect 399294 2320 399300 2372
rect 399352 2320 399358 2372
rect 399772 2360 399800 2400
rect 399846 2388 399852 2440
rect 399904 2388 399910 2440
rect 401134 2388 401140 2440
rect 401192 2388 401198 2440
rect 404648 2437 404676 2468
rect 407206 2456 407212 2508
rect 407264 2456 407270 2508
rect 408494 2496 408500 2508
rect 407776 2468 408500 2496
rect 407776 2437 407804 2468
rect 408494 2456 408500 2468
rect 408552 2456 408558 2508
rect 411806 2456 411812 2508
rect 411864 2456 411870 2508
rect 412606 2496 412634 2536
rect 422570 2524 422576 2576
rect 422628 2524 422634 2576
rect 434622 2524 434628 2576
rect 434680 2524 434686 2576
rect 434990 2524 434996 2576
rect 435048 2564 435054 2576
rect 505370 2564 505376 2576
rect 435048 2536 505376 2564
rect 435048 2524 435054 2536
rect 505370 2524 505376 2536
rect 505428 2524 505434 2576
rect 461029 2499 461087 2505
rect 461029 2496 461041 2499
rect 412606 2468 461041 2496
rect 461029 2465 461041 2468
rect 461075 2465 461087 2499
rect 461029 2459 461087 2465
rect 404633 2431 404691 2437
rect 404633 2397 404645 2431
rect 404679 2397 404691 2431
rect 404633 2391 404691 2397
rect 407761 2431 407819 2437
rect 407761 2397 407773 2431
rect 407807 2397 407819 2431
rect 407761 2391 407819 2397
rect 408310 2388 408316 2440
rect 408368 2428 408374 2440
rect 408405 2431 408463 2437
rect 408405 2428 408417 2431
rect 408368 2400 408417 2428
rect 408368 2388 408374 2400
rect 408405 2397 408417 2400
rect 408451 2428 408463 2431
rect 409325 2431 409383 2437
rect 409325 2428 409337 2431
rect 408451 2400 409337 2428
rect 408451 2397 408463 2400
rect 408405 2391 408463 2397
rect 409325 2397 409337 2400
rect 409371 2397 409383 2431
rect 409325 2391 409383 2397
rect 412361 2431 412419 2437
rect 412361 2397 412373 2431
rect 412407 2428 412419 2431
rect 412407 2400 412634 2428
rect 412407 2397 412419 2400
rect 412361 2391 412419 2397
rect 399772 2332 400996 2360
rect 400858 2292 400864 2304
rect 398668 2264 400864 2292
rect 400858 2252 400864 2264
rect 400916 2252 400922 2304
rect 400968 2292 400996 2332
rect 401502 2320 401508 2372
rect 401560 2320 401566 2372
rect 405182 2320 405188 2372
rect 405240 2320 405246 2372
rect 408681 2363 408739 2369
rect 408681 2329 408693 2363
rect 408727 2360 408739 2363
rect 409690 2360 409696 2372
rect 408727 2332 409696 2360
rect 408727 2329 408739 2332
rect 408681 2323 408739 2329
rect 409690 2320 409696 2332
rect 409748 2320 409754 2372
rect 407666 2292 407672 2304
rect 400968 2264 407672 2292
rect 407666 2252 407672 2264
rect 407724 2252 407730 2304
rect 412606 2292 412634 2400
rect 416314 2388 416320 2440
rect 416372 2428 416378 2440
rect 416777 2431 416835 2437
rect 416777 2428 416789 2431
rect 416372 2400 416789 2428
rect 416372 2388 416378 2400
rect 416777 2397 416789 2400
rect 416823 2397 416835 2431
rect 416777 2391 416835 2397
rect 421374 2388 421380 2440
rect 421432 2388 421438 2440
rect 421929 2431 421987 2437
rect 421929 2397 421941 2431
rect 421975 2428 421987 2431
rect 422570 2428 422576 2440
rect 421975 2400 422576 2428
rect 421975 2397 421987 2400
rect 421929 2391 421987 2397
rect 422570 2388 422576 2400
rect 422628 2388 422634 2440
rect 425701 2431 425759 2437
rect 425701 2397 425713 2431
rect 425747 2428 425759 2431
rect 434809 2431 434867 2437
rect 425747 2400 426572 2428
rect 425747 2397 425759 2400
rect 425701 2391 425759 2397
rect 425146 2320 425152 2372
rect 425204 2320 425210 2372
rect 426544 2304 426572 2400
rect 434809 2397 434821 2431
rect 434855 2428 434867 2431
rect 434990 2428 434996 2440
rect 434855 2400 434996 2428
rect 434855 2397 434867 2400
rect 434809 2391 434867 2397
rect 434990 2388 434996 2400
rect 435048 2388 435054 2440
rect 435726 2388 435732 2440
rect 435784 2388 435790 2440
rect 439961 2431 440019 2437
rect 439961 2397 439973 2431
rect 440007 2428 440019 2431
rect 448057 2431 448115 2437
rect 440007 2400 440648 2428
rect 440007 2397 440019 2400
rect 439961 2391 440019 2397
rect 435450 2320 435456 2372
rect 435508 2320 435514 2372
rect 439406 2320 439412 2372
rect 439464 2320 439470 2372
rect 440620 2304 440648 2400
rect 448057 2397 448069 2431
rect 448103 2428 448115 2431
rect 452841 2431 452899 2437
rect 448103 2400 448652 2428
rect 448103 2397 448115 2400
rect 448057 2391 448115 2397
rect 447778 2320 447784 2372
rect 447836 2320 447842 2372
rect 448624 2304 448652 2400
rect 452841 2397 452853 2431
rect 452887 2428 452899 2431
rect 461305 2431 461363 2437
rect 452887 2400 453436 2428
rect 452887 2397 452899 2400
rect 452841 2391 452899 2397
rect 453408 2304 453436 2400
rect 461305 2397 461317 2431
rect 461351 2428 461363 2431
rect 461351 2400 461900 2428
rect 461351 2397 461363 2400
rect 461305 2391 461363 2397
rect 461872 2304 461900 2400
rect 465718 2388 465724 2440
rect 465776 2388 465782 2440
rect 465997 2431 466055 2437
rect 465997 2397 466009 2431
rect 466043 2428 466055 2431
rect 466043 2400 466592 2428
rect 466043 2397 466055 2400
rect 465997 2391 466055 2397
rect 466564 2304 466592 2400
rect 470410 2388 470416 2440
rect 470468 2428 470474 2440
rect 470873 2431 470931 2437
rect 470873 2428 470885 2431
rect 470468 2400 470885 2428
rect 470468 2388 470474 2400
rect 470873 2397 470885 2400
rect 470919 2397 470931 2431
rect 470873 2391 470931 2397
rect 474645 2431 474703 2437
rect 474645 2397 474657 2431
rect 474691 2428 474703 2431
rect 479245 2431 479303 2437
rect 474691 2400 475516 2428
rect 474691 2397 474703 2400
rect 474645 2391 474703 2397
rect 474366 2320 474372 2372
rect 474424 2320 474430 2372
rect 475488 2304 475516 2400
rect 479245 2397 479257 2431
rect 479291 2428 479303 2431
rect 479291 2400 479840 2428
rect 479291 2397 479303 2400
rect 479245 2391 479303 2397
rect 478966 2320 478972 2372
rect 479024 2320 479030 2372
rect 479812 2304 479840 2400
rect 492401 2363 492459 2369
rect 492401 2329 492413 2363
rect 492447 2360 492459 2363
rect 492447 2332 493548 2360
rect 492447 2329 492459 2332
rect 492401 2323 492459 2329
rect 413002 2292 413008 2304
rect 412606 2264 413008 2292
rect 413002 2252 413008 2264
rect 413060 2252 413066 2304
rect 416590 2252 416596 2304
rect 416648 2252 416654 2304
rect 426526 2252 426532 2304
rect 426584 2252 426590 2304
rect 440602 2252 440608 2304
rect 440660 2252 440666 2304
rect 448606 2252 448612 2304
rect 448664 2252 448670 2304
rect 452654 2252 452660 2304
rect 452712 2252 452718 2304
rect 453390 2252 453396 2304
rect 453448 2252 453454 2304
rect 461854 2252 461860 2304
rect 461912 2252 461918 2304
rect 466546 2252 466552 2304
rect 466604 2252 466610 2304
rect 470686 2252 470692 2304
rect 470744 2252 470750 2304
rect 475470 2252 475476 2304
rect 475528 2252 475534 2304
rect 479794 2252 479800 2304
rect 479852 2252 479858 2304
rect 492122 2252 492128 2304
rect 492180 2252 492186 2304
rect 493520 2301 493548 2332
rect 493505 2295 493563 2301
rect 493505 2261 493517 2295
rect 493551 2292 493563 2295
rect 500862 2292 500868 2304
rect 493551 2264 500868 2292
rect 493551 2261 493563 2264
rect 493505 2255 493563 2261
rect 500862 2252 500868 2264
rect 500920 2252 500926 2304
rect 1104 2202 528816 2224
rect 1104 2150 67574 2202
rect 67626 2150 67638 2202
rect 67690 2150 67702 2202
rect 67754 2150 67766 2202
rect 67818 2150 67830 2202
rect 67882 2150 199502 2202
rect 199554 2150 199566 2202
rect 199618 2150 199630 2202
rect 199682 2150 199694 2202
rect 199746 2150 199758 2202
rect 199810 2150 331430 2202
rect 331482 2150 331494 2202
rect 331546 2150 331558 2202
rect 331610 2150 331622 2202
rect 331674 2150 331686 2202
rect 331738 2150 463358 2202
rect 463410 2150 463422 2202
rect 463474 2150 463486 2202
rect 463538 2150 463550 2202
rect 463602 2150 463614 2202
rect 463666 2150 528816 2202
rect 1104 2128 528816 2150
rect 26234 2048 26240 2100
rect 26292 2088 26298 2100
rect 31662 2088 31668 2100
rect 26292 2060 31668 2088
rect 26292 2048 26298 2060
rect 31662 2048 31668 2060
rect 31720 2048 31726 2100
rect 37918 2048 37924 2100
rect 37976 2088 37982 2100
rect 103882 2088 103888 2100
rect 37976 2060 103888 2088
rect 37976 2048 37982 2060
rect 103882 2048 103888 2060
rect 103940 2048 103946 2100
rect 108942 2048 108948 2100
rect 109000 2088 109006 2100
rect 202690 2088 202696 2100
rect 109000 2060 202696 2088
rect 109000 2048 109006 2060
rect 202690 2048 202696 2060
rect 202748 2048 202754 2100
rect 226150 2048 226156 2100
rect 226208 2088 226214 2100
rect 306190 2088 306196 2100
rect 226208 2060 306196 2088
rect 226208 2048 226214 2060
rect 306190 2048 306196 2060
rect 306248 2048 306254 2100
rect 307846 2048 307852 2100
rect 307904 2088 307910 2100
rect 316586 2088 316592 2100
rect 307904 2060 316592 2088
rect 307904 2048 307910 2060
rect 316586 2048 316592 2060
rect 316644 2048 316650 2100
rect 349614 2088 349620 2100
rect 316696 2060 349620 2088
rect 22646 1980 22652 2032
rect 22704 2020 22710 2032
rect 62574 2020 62580 2032
rect 22704 1992 62580 2020
rect 22704 1980 22710 1992
rect 62574 1980 62580 1992
rect 62632 1980 62638 2032
rect 70762 1980 70768 2032
rect 70820 2020 70826 2032
rect 120074 2020 120080 2032
rect 70820 1992 120080 2020
rect 70820 1980 70826 1992
rect 120074 1980 120080 1992
rect 120132 1980 120138 2032
rect 128814 1980 128820 2032
rect 128872 2020 128878 2032
rect 223022 2020 223028 2032
rect 128872 1992 223028 2020
rect 128872 1980 128878 1992
rect 223022 1980 223028 1992
rect 223080 1980 223086 2032
rect 231946 1980 231952 2032
rect 232004 2020 232010 2032
rect 306282 2020 306288 2032
rect 232004 1992 306288 2020
rect 232004 1980 232010 1992
rect 306282 1980 306288 1992
rect 306340 1980 306346 2032
rect 306466 1980 306472 2032
rect 306524 2020 306530 2032
rect 316696 2020 316724 2060
rect 349614 2048 349620 2060
rect 349672 2048 349678 2100
rect 386506 2048 386512 2100
rect 386564 2088 386570 2100
rect 478966 2088 478972 2100
rect 386564 2060 478972 2088
rect 386564 2048 386570 2060
rect 478966 2048 478972 2060
rect 479024 2048 479030 2100
rect 337194 2020 337200 2032
rect 306524 1992 316724 2020
rect 316788 1992 337200 2020
rect 306524 1980 306530 1992
rect 25958 1912 25964 1964
rect 26016 1952 26022 1964
rect 41966 1952 41972 1964
rect 26016 1924 41972 1952
rect 26016 1912 26022 1924
rect 41966 1912 41972 1924
rect 42024 1912 42030 1964
rect 42886 1912 42892 1964
rect 42944 1952 42950 1964
rect 136082 1952 136088 1964
rect 42944 1924 136088 1952
rect 42944 1912 42950 1924
rect 136082 1912 136088 1924
rect 136140 1912 136146 1964
rect 154022 1912 154028 1964
rect 154080 1952 154086 1964
rect 248046 1952 248052 1964
rect 154080 1924 248052 1952
rect 154080 1912 154086 1924
rect 248046 1912 248052 1924
rect 248104 1912 248110 1964
rect 316788 1952 316816 1992
rect 337194 1980 337200 1992
rect 337252 1980 337258 2032
rect 350534 1980 350540 2032
rect 350592 2020 350598 2032
rect 425146 2020 425152 2032
rect 350592 1992 425152 2020
rect 350592 1980 350598 1992
rect 425146 1980 425152 1992
rect 425204 1980 425210 2032
rect 426526 1980 426532 2032
rect 426584 2020 426590 2032
rect 494054 2020 494060 2032
rect 426584 1992 494060 2020
rect 426584 1980 426590 1992
rect 494054 1980 494060 1992
rect 494112 1980 494118 2032
rect 335262 1952 335268 1964
rect 311866 1924 316816 1952
rect 321526 1924 335268 1952
rect 21818 1844 21824 1896
rect 21876 1884 21882 1896
rect 66254 1884 66260 1896
rect 21876 1856 66260 1884
rect 21876 1844 21882 1856
rect 66254 1844 66260 1856
rect 66312 1844 66318 1896
rect 75270 1844 75276 1896
rect 75328 1884 75334 1896
rect 168006 1884 168012 1896
rect 75328 1856 168012 1884
rect 75328 1844 75334 1856
rect 168006 1844 168012 1856
rect 168064 1844 168070 1896
rect 200390 1844 200396 1896
rect 200448 1884 200454 1896
rect 211522 1884 211528 1896
rect 200448 1856 211528 1884
rect 200448 1844 200454 1856
rect 211522 1844 211528 1856
rect 211580 1844 211586 1896
rect 244182 1844 244188 1896
rect 244240 1884 244246 1896
rect 307754 1884 307760 1896
rect 244240 1856 307760 1884
rect 244240 1844 244246 1856
rect 307754 1844 307760 1856
rect 307812 1844 307818 1896
rect 24026 1776 24032 1828
rect 24084 1816 24090 1828
rect 31202 1816 31208 1828
rect 24084 1788 31208 1816
rect 24084 1776 24090 1788
rect 31202 1776 31208 1788
rect 31260 1776 31266 1828
rect 31404 1788 31616 1816
rect 27522 1708 27528 1760
rect 27580 1748 27586 1760
rect 31404 1748 31432 1788
rect 27580 1720 31432 1748
rect 31588 1748 31616 1788
rect 31662 1776 31668 1828
rect 31720 1816 31726 1828
rect 48314 1816 48320 1828
rect 31720 1788 48320 1816
rect 31720 1776 31726 1788
rect 48314 1776 48320 1788
rect 48372 1776 48378 1828
rect 74626 1776 74632 1828
rect 74684 1816 74690 1828
rect 111794 1816 111800 1828
rect 74684 1788 111800 1816
rect 74684 1776 74690 1788
rect 111794 1776 111800 1788
rect 111852 1776 111858 1828
rect 212166 1776 212172 1828
rect 212224 1816 212230 1828
rect 307110 1816 307116 1828
rect 212224 1788 307116 1816
rect 212224 1776 212230 1788
rect 307110 1776 307116 1788
rect 307168 1776 307174 1828
rect 311342 1776 311348 1828
rect 311400 1816 311406 1828
rect 311866 1816 311894 1924
rect 313182 1844 313188 1896
rect 313240 1884 313246 1896
rect 321526 1884 321554 1924
rect 335262 1912 335268 1924
rect 335320 1912 335326 1964
rect 349798 1912 349804 1964
rect 349856 1952 349862 1964
rect 371142 1952 371148 1964
rect 349856 1924 371148 1952
rect 349856 1912 349862 1924
rect 371142 1912 371148 1924
rect 371200 1912 371206 1964
rect 390462 1912 390468 1964
rect 390520 1952 390526 1964
rect 397822 1952 397828 1964
rect 390520 1924 397828 1952
rect 390520 1912 390526 1924
rect 397822 1912 397828 1924
rect 397880 1912 397886 1964
rect 440602 1912 440608 1964
rect 440660 1952 440666 1964
rect 488534 1952 488540 1964
rect 440660 1924 488540 1952
rect 440660 1912 440666 1924
rect 488534 1912 488540 1924
rect 488592 1912 488598 1964
rect 313240 1856 321554 1884
rect 313240 1844 313246 1856
rect 346302 1844 346308 1896
rect 346360 1884 346366 1896
rect 350626 1884 350632 1896
rect 346360 1856 350632 1884
rect 346360 1844 346366 1856
rect 350626 1844 350632 1856
rect 350684 1844 350690 1896
rect 389174 1844 389180 1896
rect 389232 1884 389238 1896
rect 399294 1884 399300 1896
rect 389232 1856 399300 1884
rect 389232 1844 389238 1856
rect 399294 1844 399300 1856
rect 399352 1844 399358 1896
rect 399478 1844 399484 1896
rect 399536 1884 399542 1896
rect 408034 1884 408040 1896
rect 399536 1856 408040 1884
rect 399536 1844 399542 1856
rect 408034 1844 408040 1856
rect 408092 1844 408098 1896
rect 448606 1844 448612 1896
rect 448664 1884 448670 1896
rect 485866 1884 485872 1896
rect 448664 1856 485872 1884
rect 448664 1844 448670 1856
rect 485866 1844 485872 1856
rect 485924 1844 485930 1896
rect 311400 1788 311894 1816
rect 311400 1776 311406 1788
rect 346670 1776 346676 1828
rect 346728 1816 346734 1828
rect 408310 1816 408316 1828
rect 346728 1788 408316 1816
rect 346728 1776 346734 1788
rect 408310 1776 408316 1788
rect 408368 1776 408374 1828
rect 453390 1776 453396 1828
rect 453448 1816 453454 1828
rect 484762 1816 484768 1828
rect 453448 1788 484768 1816
rect 453448 1776 453454 1788
rect 484762 1776 484768 1788
rect 484820 1776 484826 1828
rect 126054 1748 126060 1760
rect 31588 1720 126060 1748
rect 27580 1708 27586 1720
rect 126054 1708 126060 1720
rect 126112 1708 126118 1760
rect 127342 1708 127348 1760
rect 127400 1748 127406 1760
rect 216582 1748 216588 1760
rect 127400 1720 216588 1748
rect 127400 1708 127406 1720
rect 216582 1708 216588 1720
rect 216640 1708 216646 1760
rect 307018 1708 307024 1760
rect 307076 1748 307082 1760
rect 307076 1720 316724 1748
rect 307076 1708 307082 1720
rect 2590 1640 2596 1692
rect 2648 1680 2654 1692
rect 31386 1680 31392 1692
rect 2648 1652 31392 1680
rect 2648 1640 2654 1652
rect 31386 1640 31392 1652
rect 31444 1640 31450 1692
rect 31662 1640 31668 1692
rect 31720 1680 31726 1692
rect 96890 1680 96896 1692
rect 31720 1652 96896 1680
rect 31720 1640 31726 1652
rect 96890 1640 96896 1652
rect 96948 1640 96954 1692
rect 112898 1640 112904 1692
rect 112956 1680 112962 1692
rect 206830 1680 206836 1692
rect 112956 1652 206836 1680
rect 112956 1640 112962 1652
rect 206830 1640 206836 1652
rect 206888 1640 206894 1692
rect 208394 1640 208400 1692
rect 208452 1680 208458 1692
rect 246298 1680 246304 1692
rect 208452 1652 246304 1680
rect 208452 1640 208458 1652
rect 246298 1640 246304 1652
rect 246356 1640 246362 1692
rect 305546 1640 305552 1692
rect 305604 1680 305610 1692
rect 316696 1680 316724 1720
rect 319990 1708 319996 1760
rect 320048 1748 320054 1760
rect 329282 1748 329288 1760
rect 320048 1720 329288 1748
rect 320048 1708 320054 1720
rect 329282 1708 329288 1720
rect 329340 1708 329346 1760
rect 338022 1708 338028 1760
rect 338080 1748 338086 1760
rect 389266 1748 389272 1760
rect 338080 1720 389272 1748
rect 338080 1708 338086 1720
rect 389266 1708 389272 1720
rect 389324 1708 389330 1760
rect 399846 1708 399852 1760
rect 399904 1748 399910 1760
rect 408402 1748 408408 1760
rect 399904 1720 408408 1748
rect 399904 1708 399910 1720
rect 408402 1708 408408 1720
rect 408460 1708 408466 1760
rect 475470 1708 475476 1760
rect 475528 1748 475534 1760
rect 502334 1748 502340 1760
rect 475528 1720 502340 1748
rect 475528 1708 475534 1720
rect 502334 1708 502340 1720
rect 502392 1708 502398 1760
rect 345658 1680 345664 1692
rect 305604 1652 311894 1680
rect 316696 1652 345664 1680
rect 305604 1640 305610 1652
rect 21634 1572 21640 1624
rect 21692 1612 21698 1624
rect 24854 1612 24860 1624
rect 21692 1584 24860 1612
rect 21692 1572 21698 1584
rect 24854 1572 24860 1584
rect 24912 1572 24918 1624
rect 31478 1612 31484 1624
rect 28966 1584 31484 1612
rect 28258 1504 28264 1556
rect 28316 1544 28322 1556
rect 28966 1544 28994 1584
rect 31478 1572 31484 1584
rect 31536 1572 31542 1624
rect 115658 1572 115664 1624
rect 115716 1612 115722 1624
rect 208854 1612 208860 1624
rect 115716 1584 208860 1612
rect 115716 1572 115722 1584
rect 208854 1572 208860 1584
rect 208912 1572 208918 1624
rect 213178 1572 213184 1624
rect 213236 1612 213242 1624
rect 307386 1612 307392 1624
rect 213236 1584 307392 1612
rect 213236 1572 213242 1584
rect 307386 1572 307392 1584
rect 307444 1572 307450 1624
rect 311866 1612 311894 1652
rect 345658 1640 345664 1652
rect 345716 1640 345722 1692
rect 354490 1640 354496 1692
rect 354548 1680 354554 1692
rect 447778 1680 447784 1692
rect 354548 1652 447784 1680
rect 354548 1640 354554 1652
rect 447778 1640 447784 1652
rect 447836 1640 447842 1692
rect 466546 1640 466552 1692
rect 466604 1680 466610 1692
rect 489822 1680 489828 1692
rect 466604 1652 489828 1680
rect 466604 1640 466610 1652
rect 489822 1640 489828 1652
rect 489880 1640 489886 1692
rect 352282 1612 352288 1624
rect 311866 1584 352288 1612
rect 352282 1572 352288 1584
rect 352340 1572 352346 1624
rect 380894 1572 380900 1624
rect 380952 1612 380958 1624
rect 474366 1612 474372 1624
rect 380952 1584 474372 1612
rect 380952 1572 380958 1584
rect 474366 1572 474372 1584
rect 474424 1572 474430 1624
rect 479794 1572 479800 1624
rect 479852 1612 479858 1624
rect 496630 1612 496636 1624
rect 479852 1584 496636 1612
rect 479852 1572 479858 1584
rect 496630 1572 496636 1584
rect 496688 1572 496694 1624
rect 33686 1544 33692 1556
rect 28316 1516 28994 1544
rect 31404 1516 33692 1544
rect 28316 1504 28322 1516
rect 28074 1436 28080 1488
rect 28132 1476 28138 1488
rect 31404 1476 31432 1516
rect 33686 1504 33692 1516
rect 33744 1504 33750 1556
rect 58986 1504 58992 1556
rect 59044 1544 59050 1556
rect 152734 1544 152740 1556
rect 59044 1516 152740 1544
rect 59044 1504 59050 1516
rect 152734 1504 152740 1516
rect 152792 1504 152798 1556
rect 206094 1504 206100 1556
rect 206152 1544 206158 1556
rect 300302 1544 300308 1556
rect 206152 1516 300308 1544
rect 206152 1504 206158 1516
rect 300302 1504 300308 1516
rect 300360 1504 300366 1556
rect 306098 1504 306104 1556
rect 306156 1544 306162 1556
rect 354398 1544 354404 1556
rect 306156 1516 354404 1544
rect 306156 1504 306162 1516
rect 354398 1504 354404 1516
rect 354456 1504 354462 1556
rect 399570 1504 399576 1556
rect 399628 1544 399634 1556
rect 399628 1516 401272 1544
rect 399628 1504 399634 1516
rect 28132 1448 31432 1476
rect 28132 1436 28138 1448
rect 105078 1436 105084 1488
rect 105136 1476 105142 1488
rect 116118 1476 116124 1488
rect 105136 1448 116124 1476
rect 105136 1436 105142 1448
rect 116118 1436 116124 1448
rect 116176 1436 116182 1488
rect 120534 1436 120540 1488
rect 120592 1476 120598 1488
rect 212810 1476 212816 1488
rect 120592 1448 212816 1476
rect 120592 1436 120598 1448
rect 212810 1436 212816 1448
rect 212868 1436 212874 1488
rect 213914 1436 213920 1488
rect 213972 1476 213978 1488
rect 309226 1476 309232 1488
rect 213972 1448 309232 1476
rect 213972 1436 213978 1448
rect 309226 1436 309232 1448
rect 309284 1436 309290 1488
rect 332594 1436 332600 1488
rect 332652 1476 332658 1488
rect 401134 1476 401140 1488
rect 332652 1448 401140 1476
rect 332652 1436 332658 1448
rect 401134 1436 401140 1448
rect 401192 1436 401198 1488
rect 401244 1476 401272 1516
rect 401502 1504 401508 1556
rect 401560 1544 401566 1556
rect 407574 1544 407580 1556
rect 401560 1516 407580 1544
rect 401560 1504 401566 1516
rect 407574 1504 407580 1516
rect 407632 1504 407638 1556
rect 407666 1504 407672 1556
rect 407724 1544 407730 1556
rect 407724 1516 412634 1544
rect 407724 1504 407730 1516
rect 405090 1476 405096 1488
rect 401244 1448 405096 1476
rect 405090 1436 405096 1448
rect 405148 1436 405154 1488
rect 406930 1436 406936 1488
rect 406988 1476 406994 1488
rect 410518 1476 410524 1488
rect 406988 1448 410524 1476
rect 406988 1436 406994 1448
rect 410518 1436 410524 1448
rect 410576 1436 410582 1488
rect 28626 1368 28632 1420
rect 28684 1408 28690 1420
rect 28684 1380 31432 1408
rect 28684 1368 28690 1380
rect 23198 1300 23204 1352
rect 23256 1340 23262 1352
rect 26050 1340 26056 1352
rect 23256 1312 26056 1340
rect 23256 1300 23262 1312
rect 26050 1300 26056 1312
rect 26108 1300 26114 1352
rect 26142 1300 26148 1352
rect 26200 1340 26206 1352
rect 31018 1340 31024 1352
rect 26200 1312 31024 1340
rect 26200 1300 26206 1312
rect 31018 1300 31024 1312
rect 31076 1300 31082 1352
rect 31404 1340 31432 1380
rect 216674 1368 216680 1420
rect 216732 1408 216738 1420
rect 311526 1408 311532 1420
rect 216732 1380 311532 1408
rect 216732 1368 216738 1380
rect 311526 1368 311532 1380
rect 311584 1368 311590 1420
rect 400950 1368 400956 1420
rect 401008 1408 401014 1420
rect 402698 1408 402704 1420
rect 401008 1380 402704 1408
rect 401008 1368 401014 1380
rect 402698 1368 402704 1380
rect 402756 1368 402762 1420
rect 405182 1368 405188 1420
rect 405240 1408 405246 1420
rect 407206 1408 407212 1420
rect 405240 1380 407212 1408
rect 405240 1368 405246 1380
rect 407206 1368 407212 1380
rect 407264 1368 407270 1420
rect 412606 1408 412634 1516
rect 461854 1504 461860 1556
rect 461912 1544 461918 1556
rect 495618 1544 495624 1556
rect 461912 1516 495624 1544
rect 461912 1504 461918 1516
rect 495618 1504 495624 1516
rect 495676 1504 495682 1556
rect 480990 1476 480996 1488
rect 478708 1448 480996 1476
rect 478414 1408 478420 1420
rect 412606 1380 478420 1408
rect 478414 1368 478420 1380
rect 478472 1368 478478 1420
rect 32582 1340 32588 1352
rect 31404 1312 32588 1340
rect 32582 1300 32588 1312
rect 32640 1300 32646 1352
rect 33778 1300 33784 1352
rect 33836 1340 33842 1352
rect 117314 1340 117320 1352
rect 33836 1312 117320 1340
rect 33836 1300 33842 1312
rect 117314 1300 117320 1312
rect 117372 1300 117378 1352
rect 117866 1300 117872 1352
rect 117924 1340 117930 1352
rect 210234 1340 210240 1352
rect 117924 1312 210240 1340
rect 117924 1300 117930 1312
rect 210234 1300 210240 1312
rect 210292 1300 210298 1352
rect 306282 1300 306288 1352
rect 306340 1340 306346 1352
rect 325142 1340 325148 1352
rect 306340 1312 325148 1340
rect 306340 1300 306346 1312
rect 325142 1300 325148 1312
rect 325200 1300 325206 1352
rect 346210 1300 346216 1352
rect 346268 1340 346274 1352
rect 355962 1340 355968 1352
rect 346268 1312 355968 1340
rect 346268 1300 346274 1312
rect 355962 1300 355968 1312
rect 356020 1300 356026 1352
rect 358170 1300 358176 1352
rect 358228 1340 358234 1352
rect 407482 1340 407488 1352
rect 358228 1312 407488 1340
rect 358228 1300 358234 1312
rect 407482 1300 407488 1312
rect 407540 1300 407546 1352
rect 408402 1300 408408 1352
rect 408460 1340 408466 1352
rect 408460 1312 412634 1340
rect 408460 1300 408466 1312
rect 21910 1272 21916 1284
rect 20088 1244 21916 1272
rect 20088 864 20116 1244
rect 21910 1232 21916 1244
rect 21968 1232 21974 1284
rect 28994 1272 29000 1284
rect 22066 1244 29000 1272
rect 22066 1204 22094 1244
rect 28994 1232 29000 1244
rect 29052 1232 29058 1284
rect 30006 1232 30012 1284
rect 30064 1272 30070 1284
rect 31202 1272 31208 1284
rect 30064 1244 31208 1272
rect 30064 1232 30070 1244
rect 31202 1232 31208 1244
rect 31260 1232 31266 1284
rect 31570 1232 31576 1284
rect 31628 1272 31634 1284
rect 117498 1272 117504 1284
rect 31628 1244 117504 1272
rect 31628 1232 31634 1244
rect 117498 1232 117504 1244
rect 117556 1232 117562 1284
rect 121822 1232 121828 1284
rect 121880 1272 121886 1284
rect 215202 1272 215208 1284
rect 121880 1244 215208 1272
rect 121880 1232 121886 1244
rect 215202 1232 215208 1244
rect 215260 1232 215266 1284
rect 306006 1232 306012 1284
rect 306064 1272 306070 1284
rect 389174 1272 389180 1284
rect 306064 1244 389180 1272
rect 306064 1232 306070 1244
rect 389174 1232 389180 1244
rect 389232 1232 389238 1284
rect 394694 1232 394700 1284
rect 394752 1272 394758 1284
rect 398006 1272 398012 1284
rect 394752 1244 398012 1272
rect 394752 1232 394758 1244
rect 398006 1232 398012 1244
rect 398064 1232 398070 1284
rect 398098 1232 398104 1284
rect 398156 1272 398162 1284
rect 398156 1244 398972 1272
rect 398156 1232 398162 1244
rect 20364 1176 22094 1204
rect 22250 1176 23704 1204
rect 20364 864 20392 1176
rect 20622 1096 20628 1148
rect 20680 1096 20686 1148
rect 20624 864 20652 1096
rect 21726 932 21732 944
rect 20088 836 20208 864
rect 20364 836 20484 864
rect 20066 796 20122 800
rect 20180 796 20208 836
rect 20066 768 20208 796
rect 20338 796 20394 800
rect 20456 796 20484 836
rect 20338 768 20484 796
rect 20548 836 20652 864
rect 21284 904 21732 932
rect 20548 796 20576 836
rect 20610 796 20666 800
rect 20548 768 20666 796
rect 20066 0 20122 768
rect 20338 0 20394 768
rect 20610 0 20666 768
rect 20882 796 20938 800
rect 20990 796 20996 808
rect 20882 768 20996 796
rect 20882 0 20938 768
rect 20990 756 20996 768
rect 21048 756 21054 808
rect 21154 796 21210 800
rect 21284 796 21312 904
rect 21726 892 21732 904
rect 21784 892 21790 944
rect 22094 932 22100 944
rect 21836 904 22100 932
rect 21836 864 21864 904
rect 22094 892 22100 904
rect 22152 892 22158 944
rect 21560 836 21864 864
rect 22250 864 22278 1176
rect 23676 1068 23704 1176
rect 23750 1164 23756 1216
rect 23808 1204 23814 1216
rect 28258 1204 28264 1216
rect 23808 1176 28264 1204
rect 23808 1164 23814 1176
rect 28258 1164 28264 1176
rect 28316 1164 28322 1216
rect 31110 1204 31116 1216
rect 28644 1176 31116 1204
rect 24854 1096 24860 1148
rect 24912 1136 24918 1148
rect 28534 1136 28540 1148
rect 24912 1108 28540 1136
rect 24912 1096 24918 1108
rect 28534 1096 28540 1108
rect 28592 1096 28598 1148
rect 27614 1068 27620 1080
rect 23676 1040 27620 1068
rect 27614 1028 27620 1040
rect 27672 1028 27678 1080
rect 23382 1000 23388 1012
rect 23354 960 23388 1000
rect 23440 960 23446 1012
rect 23354 864 23382 960
rect 26234 932 26240 944
rect 22250 836 22324 864
rect 21154 768 21312 796
rect 21426 796 21482 800
rect 21560 796 21588 836
rect 21426 768 21588 796
rect 21698 796 21754 800
rect 21818 796 21824 808
rect 21698 768 21824 796
rect 21154 0 21210 768
rect 21426 0 21482 768
rect 21698 0 21754 768
rect 21818 756 21824 768
rect 21876 756 21882 808
rect 22296 800 22324 836
rect 23308 836 23382 864
rect 25148 904 26240 932
rect 21818 484 21824 536
rect 21876 524 21882 536
rect 21970 524 22026 800
rect 21876 496 22026 524
rect 21876 484 21882 496
rect 21970 0 22026 496
rect 22242 768 22324 800
rect 22514 796 22570 800
rect 22646 796 22652 808
rect 22514 768 22652 796
rect 22242 0 22298 768
rect 22514 0 22570 768
rect 22646 756 22652 768
rect 22704 756 22710 808
rect 23308 800 23336 836
rect 22786 728 22842 800
rect 22922 728 22928 740
rect 22786 700 22928 728
rect 22786 0 22842 700
rect 22922 688 22928 700
rect 22980 688 22986 740
rect 23058 728 23114 800
rect 23308 768 23386 800
rect 23198 728 23204 740
rect 23058 700 23204 728
rect 23058 0 23114 700
rect 23198 688 23204 700
rect 23256 688 23262 740
rect 23330 0 23386 768
rect 23602 796 23658 800
rect 23750 796 23756 808
rect 23602 768 23756 796
rect 23602 0 23658 768
rect 23750 756 23756 768
rect 23808 756 23814 808
rect 23874 728 23930 800
rect 24146 796 24202 800
rect 24302 796 24308 808
rect 24146 768 24308 796
rect 24026 728 24032 740
rect 23874 700 24032 728
rect 23874 0 23930 700
rect 24026 688 24032 700
rect 24084 688 24090 740
rect 24146 0 24202 768
rect 24302 756 24308 768
rect 24360 756 24366 808
rect 24418 796 24474 800
rect 24578 796 24584 808
rect 24418 768 24584 796
rect 24418 0 24474 768
rect 24578 756 24584 768
rect 24636 756 24642 808
rect 24690 796 24746 800
rect 24854 796 24860 808
rect 24690 768 24860 796
rect 24690 0 24746 768
rect 24854 756 24860 768
rect 24912 756 24918 808
rect 24962 796 25018 800
rect 25148 796 25176 904
rect 26234 892 26240 904
rect 26292 892 26298 944
rect 27614 932 27620 944
rect 26988 904 27620 932
rect 26418 864 26424 876
rect 25700 836 26424 864
rect 24962 768 25176 796
rect 25234 796 25290 800
rect 25406 796 25412 808
rect 25234 768 25412 796
rect 24962 0 25018 768
rect 25234 0 25290 768
rect 25406 756 25412 768
rect 25464 756 25470 808
rect 25506 796 25562 800
rect 25700 796 25728 836
rect 26418 824 26424 836
rect 26476 824 26482 876
rect 26988 864 27016 904
rect 27614 892 27620 904
rect 27672 892 27678 944
rect 28644 932 28672 1176
rect 31110 1164 31116 1176
rect 31168 1164 31174 1216
rect 36630 1164 36636 1216
rect 36688 1204 36694 1216
rect 108390 1204 108396 1216
rect 36688 1176 108396 1204
rect 36688 1164 36694 1176
rect 108390 1164 108396 1176
rect 108448 1164 108454 1216
rect 120074 1164 120080 1216
rect 120132 1204 120138 1216
rect 160462 1204 160468 1216
rect 120132 1176 160468 1204
rect 120132 1164 120138 1176
rect 160462 1164 160468 1176
rect 160520 1164 160526 1216
rect 161842 1164 161848 1216
rect 161900 1204 161906 1216
rect 255774 1204 255780 1216
rect 161900 1176 255780 1204
rect 161900 1164 161906 1176
rect 255774 1164 255780 1176
rect 255832 1164 255838 1216
rect 306190 1164 306196 1216
rect 306248 1204 306254 1216
rect 319438 1204 319444 1216
rect 306248 1176 319444 1204
rect 306248 1164 306254 1176
rect 319438 1164 319444 1176
rect 319496 1164 319502 1216
rect 323762 1164 323768 1216
rect 323820 1204 323826 1216
rect 398834 1204 398840 1216
rect 323820 1176 398840 1204
rect 323820 1164 323826 1176
rect 398834 1164 398840 1176
rect 398892 1164 398898 1216
rect 398944 1204 398972 1244
rect 399018 1232 399024 1284
rect 399076 1272 399082 1284
rect 412606 1272 412634 1312
rect 435726 1300 435732 1352
rect 435784 1340 435790 1352
rect 478708 1340 478736 1448
rect 480990 1436 480996 1448
rect 481048 1436 481054 1488
rect 478782 1368 478788 1420
rect 478840 1408 478846 1420
rect 492122 1408 492128 1420
rect 478840 1380 492128 1408
rect 478840 1368 478846 1380
rect 492122 1368 492128 1380
rect 492180 1368 492186 1420
rect 435784 1312 478736 1340
rect 435784 1300 435790 1312
rect 479610 1300 479616 1352
rect 479668 1340 479674 1352
rect 484670 1340 484676 1352
rect 479668 1312 484676 1340
rect 479668 1300 479674 1312
rect 484670 1300 484676 1312
rect 484728 1300 484734 1352
rect 484762 1300 484768 1352
rect 484820 1340 484826 1352
rect 484820 1312 489914 1340
rect 484820 1300 484826 1312
rect 480346 1272 480352 1284
rect 399076 1244 407528 1272
rect 412606 1244 480352 1272
rect 399076 1232 399082 1244
rect 401042 1204 401048 1216
rect 398944 1176 401048 1204
rect 401042 1164 401048 1176
rect 401100 1164 401106 1216
rect 401134 1164 401140 1216
rect 401192 1204 401198 1216
rect 407500 1204 407528 1244
rect 480346 1232 480352 1244
rect 480404 1232 480410 1284
rect 480898 1232 480904 1284
rect 480956 1272 480962 1284
rect 485774 1272 485780 1284
rect 480956 1244 485780 1272
rect 480956 1232 480962 1244
rect 485774 1232 485780 1244
rect 485832 1232 485838 1284
rect 485866 1232 485872 1284
rect 485924 1272 485930 1284
rect 488810 1272 488816 1284
rect 485924 1244 488816 1272
rect 485924 1232 485930 1244
rect 488810 1232 488816 1244
rect 488868 1232 488874 1284
rect 489886 1272 489914 1312
rect 494698 1300 494704 1352
rect 494756 1340 494762 1352
rect 494756 1312 508360 1340
rect 494756 1300 494762 1312
rect 489886 1244 507256 1272
rect 401192 1176 407068 1204
rect 407500 1176 412634 1204
rect 401192 1164 401198 1176
rect 31202 1136 31208 1148
rect 29334 1108 31208 1136
rect 29086 932 29092 944
rect 27724 904 28672 932
rect 28966 904 29092 932
rect 27724 864 27752 904
rect 28626 864 28632 876
rect 26528 836 27016 864
rect 27264 836 27752 864
rect 27816 836 28632 864
rect 25506 768 25728 796
rect 25778 796 25834 800
rect 25958 796 25964 808
rect 25778 768 25964 796
rect 25506 0 25562 768
rect 25778 0 25834 768
rect 25958 756 25964 768
rect 26016 756 26022 808
rect 26050 796 26106 800
rect 26142 796 26148 808
rect 26050 768 26148 796
rect 26050 0 26106 768
rect 26142 756 26148 768
rect 26200 756 26206 808
rect 26322 796 26378 800
rect 26528 796 26556 836
rect 26322 768 26556 796
rect 26594 796 26650 800
rect 26694 796 26700 808
rect 26594 768 26700 796
rect 26322 0 26378 768
rect 26594 0 26650 768
rect 26694 756 26700 768
rect 26752 756 26758 808
rect 26866 796 26922 800
rect 26970 796 26976 808
rect 26866 768 26976 796
rect 26866 0 26922 768
rect 26970 756 26976 768
rect 27028 756 27034 808
rect 27138 796 27194 800
rect 27264 796 27292 836
rect 27138 768 27292 796
rect 27410 796 27466 800
rect 27522 796 27528 808
rect 27410 768 27528 796
rect 27138 0 27194 768
rect 27410 0 27466 768
rect 27522 756 27528 768
rect 27580 756 27586 808
rect 27682 796 27738 800
rect 27816 796 27844 836
rect 28626 824 28632 836
rect 28684 824 28690 876
rect 27682 768 27844 796
rect 27954 796 28010 800
rect 28074 796 28080 808
rect 27954 768 28080 796
rect 27682 0 27738 768
rect 27954 0 28010 768
rect 28074 756 28080 768
rect 28132 756 28138 808
rect 28226 796 28282 800
rect 28350 796 28356 808
rect 28226 768 28356 796
rect 28226 0 28282 768
rect 28350 756 28356 768
rect 28408 756 28414 808
rect 28498 456 28554 800
rect 28770 660 28826 800
rect 28966 660 28994 904
rect 29086 892 29092 904
rect 29144 892 29150 944
rect 29334 864 29362 1108
rect 31202 1096 31208 1108
rect 31260 1096 31266 1148
rect 31478 1096 31484 1148
rect 31536 1136 31542 1148
rect 118142 1136 118148 1148
rect 31536 1108 118148 1136
rect 31536 1096 31542 1108
rect 118142 1096 118148 1108
rect 118200 1096 118206 1148
rect 182910 1096 182916 1148
rect 182968 1136 182974 1148
rect 277118 1136 277124 1148
rect 182968 1108 277124 1136
rect 182968 1096 182974 1108
rect 277118 1096 277124 1108
rect 277176 1096 277182 1148
rect 318978 1096 318984 1148
rect 319036 1136 319042 1148
rect 399662 1136 399668 1148
rect 319036 1108 399668 1136
rect 319036 1096 319042 1108
rect 399662 1096 399668 1108
rect 399720 1096 399726 1148
rect 402698 1096 402704 1148
rect 402756 1136 402762 1148
rect 406746 1136 406752 1148
rect 402756 1108 406752 1136
rect 402756 1096 402762 1108
rect 406746 1096 406752 1108
rect 406804 1096 406810 1148
rect 30006 1068 30012 1080
rect 29886 1040 30012 1068
rect 29886 864 29914 1040
rect 30006 1028 30012 1040
rect 30064 1028 30070 1080
rect 36814 1068 36820 1080
rect 30144 1040 36820 1068
rect 30144 864 30172 1040
rect 36814 1028 36820 1040
rect 36872 1028 36878 1080
rect 119982 1028 119988 1080
rect 120040 1068 120046 1080
rect 211062 1068 211068 1080
rect 120040 1040 211068 1068
rect 120040 1028 120046 1040
rect 211062 1028 211068 1040
rect 211120 1028 211126 1080
rect 237006 1028 237012 1080
rect 237064 1068 237070 1080
rect 331214 1068 331220 1080
rect 237064 1040 331220 1068
rect 237064 1028 237070 1040
rect 331214 1028 331220 1040
rect 331272 1028 331278 1080
rect 341518 1028 341524 1080
rect 341576 1068 341582 1080
rect 390554 1068 390560 1080
rect 341576 1040 390560 1068
rect 341576 1028 341582 1040
rect 390554 1028 390560 1040
rect 390612 1028 390618 1080
rect 397914 1028 397920 1080
rect 397972 1068 397978 1080
rect 399570 1068 399576 1080
rect 397972 1040 399576 1068
rect 397972 1028 397978 1040
rect 399570 1028 399576 1040
rect 399628 1028 399634 1080
rect 399754 1028 399760 1080
rect 399812 1068 399818 1080
rect 400950 1068 400956 1080
rect 399812 1040 400956 1068
rect 399812 1028 399818 1040
rect 400950 1028 400956 1040
rect 401008 1028 401014 1080
rect 406930 1068 406936 1080
rect 401244 1040 406936 1068
rect 30416 972 31708 1000
rect 30416 864 30444 972
rect 31680 932 31708 972
rect 31754 960 31760 1012
rect 31812 1000 31818 1012
rect 112346 1000 112352 1012
rect 31812 972 112352 1000
rect 31812 960 31818 972
rect 112346 960 112352 972
rect 112404 960 112410 1012
rect 116118 960 116124 1012
rect 116176 1000 116182 1012
rect 197906 1000 197912 1012
rect 116176 972 197912 1000
rect 116176 960 116182 972
rect 197906 960 197912 972
rect 197964 960 197970 1012
rect 199378 960 199384 1012
rect 199436 1000 199442 1012
rect 292574 1000 292580 1012
rect 199436 972 292580 1000
rect 199436 960 199442 972
rect 292574 960 292580 972
rect 292632 960 292638 1012
rect 299566 960 299572 1012
rect 299624 1000 299630 1012
rect 393866 1000 393872 1012
rect 299624 972 393872 1000
rect 299624 960 299630 972
rect 393866 960 393872 972
rect 393924 960 393930 1012
rect 401134 1000 401140 1012
rect 396046 972 401140 1000
rect 36446 932 36452 944
rect 29288 836 29362 864
rect 29840 836 29914 864
rect 30024 836 30172 864
rect 30300 836 30444 864
rect 30852 904 31616 932
rect 31680 904 36452 932
rect 28770 632 28994 660
rect 29042 796 29098 800
rect 29178 796 29184 808
rect 29042 768 29184 796
rect 28626 456 28632 468
rect 28498 428 28632 456
rect 28498 0 28554 428
rect 28626 416 28632 428
rect 28684 416 28690 468
rect 28770 0 28826 632
rect 29042 0 29098 768
rect 29178 756 29184 768
rect 29236 756 29242 808
rect 29288 800 29316 836
rect 29288 768 29370 800
rect 29314 0 29370 768
rect 29586 796 29642 800
rect 29730 796 29736 808
rect 29586 768 29736 796
rect 29586 0 29642 768
rect 29730 756 29736 768
rect 29788 756 29794 808
rect 29840 800 29868 836
rect 29840 768 29914 800
rect 30024 796 30052 836
rect 30130 796 30186 800
rect 30024 768 30186 796
rect 30300 796 30328 836
rect 30402 796 30458 800
rect 30300 768 30458 796
rect 29858 0 29914 768
rect 30130 0 30186 768
rect 30402 0 30458 768
rect 30674 796 30730 800
rect 30852 796 30880 904
rect 31294 864 31300 876
rect 31128 836 31300 864
rect 30674 768 30880 796
rect 30946 796 31002 800
rect 31128 796 31156 836
rect 31294 824 31300 836
rect 31352 824 31358 876
rect 30946 768 31156 796
rect 30674 0 30730 768
rect 30946 0 31002 768
rect 31218 116 31274 800
rect 31588 524 31616 904
rect 36446 892 36452 904
rect 36504 892 36510 944
rect 36538 892 36544 944
rect 36596 932 36602 944
rect 122834 932 122840 944
rect 36596 904 122840 932
rect 36596 892 36602 904
rect 122834 892 122840 904
rect 122892 892 122898 944
rect 210786 892 210792 944
rect 210844 932 210850 944
rect 305178 932 305184 944
rect 210844 904 305184 932
rect 210844 892 210850 904
rect 305178 892 305184 904
rect 305236 892 305242 944
rect 307754 892 307760 944
rect 307812 932 307818 944
rect 337838 932 337844 944
rect 307812 904 337844 932
rect 307812 892 307818 904
rect 337838 892 337844 904
rect 337896 892 337902 944
rect 391658 892 391664 944
rect 391716 932 391722 944
rect 396046 932 396074 972
rect 401134 960 401140 972
rect 401192 960 401198 1012
rect 391716 904 396074 932
rect 391716 892 391722 904
rect 398006 892 398012 944
rect 398064 932 398070 944
rect 401244 932 401272 1040
rect 406930 1028 406936 1040
rect 406988 1028 406994 1080
rect 401428 972 406516 1000
rect 398064 904 401272 932
rect 398064 892 398070 904
rect 401318 892 401324 944
rect 401376 932 401382 944
rect 401428 932 401456 972
rect 406378 932 406384 944
rect 401376 904 401456 932
rect 401520 904 406384 932
rect 401376 892 401382 904
rect 31662 824 31668 876
rect 31720 864 31726 876
rect 31754 864 31760 876
rect 31720 836 31760 864
rect 31720 824 31726 836
rect 31754 824 31760 836
rect 31812 824 31818 876
rect 31846 824 31852 876
rect 31904 864 31910 876
rect 121638 864 121644 876
rect 31904 836 121644 864
rect 31904 824 31910 836
rect 121638 824 121644 836
rect 121696 824 121702 876
rect 157886 824 157892 876
rect 157944 864 157950 876
rect 251726 864 251732 876
rect 157944 836 251732 864
rect 157944 824 157950 836
rect 251726 824 251732 836
rect 251784 824 251790 876
rect 254302 824 254308 876
rect 254360 864 254366 876
rect 306742 864 306748 876
rect 254360 836 306748 864
rect 254360 824 254366 836
rect 306742 824 306748 836
rect 306800 824 306806 876
rect 313366 824 313372 876
rect 313424 864 313430 876
rect 313424 836 393314 864
rect 313424 824 313430 836
rect 36814 756 36820 808
rect 36872 796 36878 808
rect 123846 796 123852 808
rect 36872 768 123852 796
rect 36872 756 36878 768
rect 123846 756 123852 768
rect 123904 756 123910 808
rect 165522 756 165528 808
rect 165580 796 165586 808
rect 258350 796 258356 808
rect 165580 768 258356 796
rect 165580 756 165586 768
rect 258350 756 258356 768
rect 258408 756 258414 808
rect 265710 756 265716 808
rect 265768 796 265774 808
rect 357894 796 357900 808
rect 265768 768 357900 796
rect 265768 756 265774 768
rect 357894 756 357900 768
rect 357952 756 357958 808
rect 111794 688 111800 740
rect 111852 728 111858 740
rect 169018 728 169024 740
rect 111852 700 169024 728
rect 111852 688 111858 700
rect 169018 688 169024 700
rect 169076 688 169082 740
rect 257062 688 257068 740
rect 257120 728 257126 740
rect 346302 728 346308 740
rect 257120 700 346308 728
rect 257120 688 257126 700
rect 346302 688 346308 700
rect 346360 688 346366 740
rect 393286 728 393314 836
rect 398190 824 398196 876
rect 398248 864 398254 876
rect 401520 864 401548 904
rect 406378 892 406384 904
rect 406436 892 406442 944
rect 398248 836 401548 864
rect 398248 824 398254 836
rect 401594 824 401600 876
rect 401652 864 401658 876
rect 406488 864 406516 972
rect 407040 932 407068 1176
rect 407482 1096 407488 1148
rect 407540 1136 407546 1148
rect 408862 1136 408868 1148
rect 407540 1108 408868 1136
rect 407540 1096 407546 1108
rect 408862 1096 408868 1108
rect 408920 1096 408926 1148
rect 411438 1068 411444 1080
rect 407500 1040 411444 1068
rect 407206 960 407212 1012
rect 407264 1000 407270 1012
rect 407500 1000 407528 1040
rect 411438 1028 411444 1040
rect 411496 1028 411502 1080
rect 412606 1068 412634 1176
rect 413002 1164 413008 1216
rect 413060 1204 413066 1216
rect 486878 1204 486884 1216
rect 413060 1176 486884 1204
rect 413060 1164 413066 1176
rect 486878 1164 486884 1176
rect 486936 1164 486942 1216
rect 488534 1164 488540 1216
rect 488592 1204 488598 1216
rect 500126 1204 500132 1216
rect 488592 1176 500132 1204
rect 488592 1164 488598 1176
rect 500126 1164 500132 1176
rect 500184 1164 500190 1216
rect 416590 1096 416596 1148
rect 416648 1136 416654 1148
rect 416648 1108 499574 1136
rect 416648 1096 416654 1108
rect 480898 1068 480904 1080
rect 412606 1040 480904 1068
rect 480898 1028 480904 1040
rect 480956 1028 480962 1080
rect 480990 1028 480996 1080
rect 481048 1068 481054 1080
rect 482554 1068 482560 1080
rect 481048 1040 482560 1068
rect 481048 1028 481054 1040
rect 482554 1028 482560 1040
rect 482612 1028 482618 1080
rect 482646 1028 482652 1080
rect 482704 1068 482710 1080
rect 494698 1068 494704 1080
rect 482704 1040 494704 1068
rect 482704 1028 482710 1040
rect 494698 1028 494704 1040
rect 494756 1028 494762 1080
rect 499546 1068 499574 1108
rect 499546 1040 505094 1068
rect 407264 972 407528 1000
rect 407264 960 407270 972
rect 407574 960 407580 1012
rect 407632 1000 407638 1012
rect 494514 1000 494520 1012
rect 407632 972 494520 1000
rect 407632 960 407638 972
rect 494514 960 494520 972
rect 494572 960 494578 1012
rect 494900 972 499574 1000
rect 479610 932 479616 944
rect 407040 904 479616 932
rect 479610 892 479616 904
rect 479668 892 479674 944
rect 479702 892 479708 944
rect 479760 932 479766 944
rect 494900 932 494928 972
rect 499546 932 499574 972
rect 479760 904 494928 932
rect 495084 904 495204 932
rect 499546 904 500816 932
rect 479760 892 479766 904
rect 401652 836 401916 864
rect 406488 836 409184 864
rect 401652 824 401658 836
rect 397822 756 397828 808
rect 397880 796 397886 808
rect 400050 796 400106 800
rect 397880 768 400106 796
rect 397880 756 397886 768
rect 399294 728 399300 740
rect 393286 700 399300 728
rect 399294 688 399300 700
rect 399352 688 399358 740
rect 32858 620 32864 672
rect 32916 660 32922 672
rect 117590 660 117596 672
rect 32916 632 117596 660
rect 32916 620 32922 632
rect 117590 620 117596 632
rect 117648 620 117654 672
rect 120350 620 120356 672
rect 120408 660 120414 672
rect 211430 660 211436 672
rect 120408 632 211436 660
rect 120408 620 120414 632
rect 211430 620 211436 632
rect 211488 620 211494 672
rect 212442 620 212448 672
rect 212500 660 212506 672
rect 305454 660 305460 672
rect 212500 632 305460 660
rect 212500 620 212506 632
rect 305454 620 305460 632
rect 305512 620 305518 672
rect 307294 620 307300 672
rect 307352 660 307358 672
rect 332594 660 332600 672
rect 307352 632 332600 660
rect 307352 620 307358 632
rect 332594 620 332600 632
rect 332652 620 332658 672
rect 332778 620 332784 672
rect 332836 660 332842 672
rect 350534 660 350540 672
rect 332836 632 350540 660
rect 332836 620 332842 632
rect 350534 620 350540 632
rect 350592 620 350598 672
rect 395982 620 395988 672
rect 396040 660 396046 672
rect 399938 660 399944 672
rect 396040 632 399944 660
rect 396040 620 396046 632
rect 399938 620 399944 632
rect 399996 620 400002 672
rect 36446 552 36452 604
rect 36504 592 36510 604
rect 125042 592 125048 604
rect 36504 564 125048 592
rect 36504 552 36510 564
rect 125042 552 125048 564
rect 125100 552 125106 604
rect 146110 552 146116 604
rect 146168 592 146174 604
rect 204898 592 204904 604
rect 146168 564 204904 592
rect 146168 552 146174 564
rect 204898 552 204904 564
rect 204956 552 204962 604
rect 206186 552 206192 604
rect 206244 592 206250 604
rect 299014 592 299020 604
rect 206244 564 299020 592
rect 206244 552 206250 564
rect 299014 552 299020 564
rect 299072 552 299078 604
rect 324682 552 324688 604
rect 324740 592 324746 604
rect 397914 592 397920 604
rect 324740 564 397920 592
rect 324740 552 324746 564
rect 397914 552 397920 564
rect 397972 552 397978 604
rect 36630 524 36636 536
rect 31588 496 36636 524
rect 36630 484 36636 496
rect 36688 484 36694 536
rect 193582 484 193588 536
rect 193640 524 193646 536
rect 285950 524 285956 536
rect 193640 496 285956 524
rect 193640 484 193646 496
rect 285950 484 285956 496
rect 286008 484 286014 536
rect 295794 484 295800 536
rect 295852 524 295858 536
rect 338022 524 338028 536
rect 295852 496 338028 524
rect 295852 484 295858 496
rect 338022 484 338028 496
rect 338080 484 338086 536
rect 33686 416 33692 468
rect 33744 456 33750 468
rect 121454 456 121460 468
rect 33744 428 121460 456
rect 33744 416 33750 428
rect 121454 416 121460 428
rect 121512 416 121518 468
rect 152182 416 152188 468
rect 152240 456 152246 468
rect 208394 456 208400 468
rect 152240 428 208400 456
rect 152240 416 152246 428
rect 208394 416 208400 428
rect 208452 416 208458 468
rect 258258 416 258264 468
rect 258316 456 258322 468
rect 346578 456 346584 468
rect 258316 428 346584 456
rect 258316 416 258322 428
rect 346578 416 346584 428
rect 346636 416 346642 468
rect 356054 416 356060 468
rect 356112 456 356118 468
rect 398006 456 398012 468
rect 356112 428 398012 456
rect 356112 416 356118 428
rect 398006 416 398012 428
rect 398064 416 398070 468
rect 170766 348 170772 400
rect 170824 388 170830 400
rect 264330 388 264336 400
rect 170824 360 264336 388
rect 170824 348 170830 360
rect 264330 348 264336 360
rect 264388 348 264394 400
rect 278314 348 278320 400
rect 278372 388 278378 400
rect 349798 388 349804 400
rect 278372 360 349804 388
rect 278372 348 278378 360
rect 349798 348 349804 360
rect 349856 348 349862 400
rect 352374 348 352380 400
rect 352432 388 352438 400
rect 398190 388 398196 400
rect 352432 360 398196 388
rect 352432 348 352438 360
rect 398190 348 398196 360
rect 398248 348 398254 400
rect 32582 280 32588 332
rect 32640 320 32646 332
rect 121546 320 121552 332
rect 32640 292 121552 320
rect 32640 280 32646 292
rect 121546 280 121552 292
rect 121604 280 121610 332
rect 121730 280 121736 332
rect 121788 320 121794 332
rect 212626 320 212632 332
rect 121788 292 212632 320
rect 121788 280 121794 292
rect 212626 280 212632 292
rect 212684 280 212690 332
rect 247126 280 247132 332
rect 247184 320 247190 332
rect 339954 320 339960 332
rect 247184 292 339960 320
rect 247184 280 247190 292
rect 339954 280 339960 292
rect 340012 280 340018 332
rect 349706 280 349712 332
rect 349764 320 349770 332
rect 398098 320 398104 332
rect 349764 292 398104 320
rect 349764 280 349770 292
rect 398098 280 398104 292
rect 398156 280 398162 332
rect 31386 212 31392 264
rect 31444 252 31450 264
rect 118694 252 118700 264
rect 31444 224 118700 252
rect 31444 212 31450 224
rect 118694 212 118700 224
rect 118752 212 118758 264
rect 218422 212 218428 264
rect 218480 252 218486 264
rect 313274 252 313280 264
rect 218480 224 313280 252
rect 218480 212 218486 224
rect 313274 212 313280 224
rect 313332 212 313338 264
rect 348418 212 348424 264
rect 348476 252 348482 264
rect 399846 252 399852 264
rect 348476 224 399852 252
rect 348476 212 348482 224
rect 399846 212 399852 224
rect 399904 212 399910 264
rect 31570 144 31576 196
rect 31628 184 31634 196
rect 120166 184 120172 196
rect 31628 156 120172 184
rect 31628 144 31634 156
rect 120166 144 120172 156
rect 120224 144 120230 196
rect 215846 144 215852 196
rect 215904 184 215910 196
rect 310422 184 310428 196
rect 215904 156 310428 184
rect 215904 144 215910 156
rect 310422 144 310428 156
rect 310480 144 310486 196
rect 346762 144 346768 196
rect 346820 184 346826 196
rect 399478 184 399484 196
rect 346820 156 399484 184
rect 346820 144 346826 156
rect 399478 144 399484 156
rect 399536 144 399542 196
rect 125226 116 125232 128
rect 31218 88 125232 116
rect 31218 0 31274 88
rect 125226 76 125232 88
rect 125284 76 125290 128
rect 337286 76 337292 128
rect 337344 116 337350 128
rect 399754 116 399760 128
rect 337344 88 399760 116
rect 337344 76 337350 88
rect 399754 76 399760 88
rect 399812 76 399818 128
rect 31754 8 31760 60
rect 31812 48 31818 60
rect 123754 48 123760 60
rect 31812 20 123760 48
rect 31812 8 31818 20
rect 123754 8 123760 20
rect 123812 8 123818 60
rect 315758 8 315764 60
rect 315816 48 315822 60
rect 399938 48 399944 60
rect 315816 20 399944 48
rect 315816 8 315822 20
rect 399938 8 399944 20
rect 399996 8 400002 60
rect 400050 0 400106 768
rect 400214 620 400220 672
rect 400272 660 400278 672
rect 400322 660 400378 800
rect 400272 632 400378 660
rect 400272 620 400278 632
rect 400322 0 400378 632
rect 400490 416 400496 468
rect 400548 456 400554 468
rect 400594 456 400650 800
rect 400766 756 400772 808
rect 400824 796 400830 808
rect 400866 796 400922 800
rect 400824 768 400922 796
rect 400824 756 400830 768
rect 400548 428 400650 456
rect 400548 416 400554 428
rect 400594 0 400650 428
rect 400866 0 400922 768
rect 400950 756 400956 808
rect 401008 796 401014 808
rect 401138 796 401194 800
rect 401008 768 401194 796
rect 401008 756 401014 768
rect 401138 0 401194 768
rect 401318 756 401324 808
rect 401376 796 401382 808
rect 401410 796 401466 800
rect 401376 768 401466 796
rect 401376 756 401382 768
rect 401410 0 401466 768
rect 401682 796 401738 800
rect 401778 796 401784 808
rect 401682 768 401784 796
rect 401682 0 401738 768
rect 401778 756 401784 768
rect 401836 756 401842 808
rect 401888 796 401916 836
rect 401954 796 402010 800
rect 401888 768 402010 796
rect 401954 0 402010 768
rect 402054 756 402060 808
rect 402112 796 402118 808
rect 402226 796 402282 800
rect 402112 768 402282 796
rect 402112 756 402118 768
rect 402226 0 402282 768
rect 402330 756 402336 808
rect 402388 796 402394 808
rect 402498 796 402554 800
rect 402388 768 402554 796
rect 402388 756 402394 768
rect 402498 0 402554 768
rect 402606 756 402612 808
rect 402664 796 402670 808
rect 402770 796 402826 800
rect 402664 768 402826 796
rect 402664 756 402670 768
rect 402770 0 402826 768
rect 403042 796 403098 800
rect 403158 796 403164 808
rect 403042 768 403164 796
rect 403042 0 403098 768
rect 403158 756 403164 768
rect 403216 756 403222 808
rect 403314 660 403370 800
rect 403434 660 403440 672
rect 403314 632 403440 660
rect 403314 0 403370 632
rect 403434 620 403440 632
rect 403492 620 403498 672
rect 403434 484 403440 536
rect 403492 524 403498 536
rect 403586 524 403642 800
rect 403710 756 403716 808
rect 403768 796 403774 808
rect 403858 796 403914 800
rect 403768 768 403914 796
rect 403768 756 403774 768
rect 403492 496 403642 524
rect 403492 484 403498 496
rect 403586 0 403642 496
rect 403858 0 403914 768
rect 403986 756 403992 808
rect 404044 796 404050 808
rect 404130 796 404186 800
rect 404044 768 404186 796
rect 404044 756 404050 768
rect 404130 0 404186 768
rect 404262 756 404268 808
rect 404320 796 404326 808
rect 404402 796 404458 800
rect 404320 768 404458 796
rect 404320 756 404326 768
rect 404402 0 404458 768
rect 404538 756 404544 808
rect 404596 796 404602 808
rect 404674 796 404730 800
rect 404596 768 404730 796
rect 404596 756 404602 768
rect 404674 0 404730 768
rect 404814 756 404820 808
rect 404872 796 404878 808
rect 404946 796 405002 800
rect 404872 768 405002 796
rect 404872 756 404878 768
rect 404946 0 405002 768
rect 405090 756 405096 808
rect 405148 796 405154 808
rect 405218 796 405274 800
rect 405148 768 405274 796
rect 405148 756 405154 768
rect 405218 0 405274 768
rect 405366 756 405372 808
rect 405424 796 405430 808
rect 405490 796 405546 800
rect 405424 768 405546 796
rect 405424 756 405430 768
rect 405490 0 405546 768
rect 405762 796 405818 800
rect 405918 796 405924 808
rect 405762 768 405924 796
rect 405762 0 405818 768
rect 405918 756 405924 768
rect 405976 756 405982 808
rect 406034 524 406090 800
rect 406194 756 406200 808
rect 406252 796 406258 808
rect 406306 796 406362 800
rect 406252 768 406362 796
rect 406252 756 406258 768
rect 406194 524 406200 536
rect 406034 496 406200 524
rect 406034 0 406090 496
rect 406194 484 406200 496
rect 406252 484 406258 536
rect 406306 0 406362 768
rect 406470 756 406476 808
rect 406528 796 406534 808
rect 406578 796 406634 800
rect 406528 768 406634 796
rect 406528 756 406534 768
rect 406578 0 406634 768
rect 406746 756 406752 808
rect 406804 796 406810 808
rect 406850 796 406906 800
rect 406804 768 406906 796
rect 406804 756 406810 768
rect 406850 0 406906 768
rect 407122 796 407178 800
rect 407206 796 407212 808
rect 407122 768 407212 796
rect 407122 0 407178 768
rect 407206 756 407212 768
rect 407264 756 407270 808
rect 407298 756 407304 808
rect 407356 796 407362 808
rect 407394 796 407450 800
rect 407356 768 407450 796
rect 407356 756 407362 768
rect 407394 0 407450 768
rect 407666 660 407722 800
rect 407758 756 407764 808
rect 407816 796 407822 808
rect 407938 796 407994 800
rect 407816 768 407994 796
rect 407816 756 407822 768
rect 407758 660 407764 672
rect 407666 632 407764 660
rect 407666 0 407722 632
rect 407758 620 407764 632
rect 407816 620 407822 672
rect 407938 0 407994 768
rect 408034 756 408040 808
rect 408092 796 408098 808
rect 408210 796 408266 800
rect 408092 768 408266 796
rect 408092 756 408098 768
rect 408210 0 408266 768
rect 408310 756 408316 808
rect 408368 796 408374 808
rect 408482 796 408538 800
rect 408368 768 408538 796
rect 408368 756 408374 768
rect 408482 0 408538 768
rect 408586 756 408592 808
rect 408644 796 408650 808
rect 408754 796 408810 800
rect 408644 768 408810 796
rect 408644 756 408650 768
rect 408754 0 408810 768
rect 408862 756 408868 808
rect 408920 796 408926 808
rect 409026 796 409082 800
rect 408920 768 409082 796
rect 409156 796 409184 836
rect 409690 824 409696 876
rect 409748 864 409754 876
rect 409748 836 411392 864
rect 409748 824 409754 836
rect 409298 796 409354 800
rect 409156 768 409354 796
rect 408920 756 408926 768
rect 409026 0 409082 768
rect 409298 0 409354 768
rect 409414 756 409420 808
rect 409472 796 409478 808
rect 409570 796 409626 800
rect 409472 768 409626 796
rect 409472 756 409478 768
rect 409570 0 409626 768
rect 409690 484 409696 536
rect 409748 524 409754 536
rect 409842 524 409898 800
rect 409966 756 409972 808
rect 410024 796 410030 808
rect 410114 796 410170 800
rect 410024 768 410170 796
rect 410024 756 410030 768
rect 409748 496 409898 524
rect 409748 484 409754 496
rect 409842 0 409898 496
rect 410114 0 410170 768
rect 410242 756 410248 808
rect 410300 796 410306 808
rect 410386 796 410442 800
rect 410300 768 410442 796
rect 410300 756 410306 768
rect 410386 0 410442 768
rect 410518 756 410524 808
rect 410576 796 410582 808
rect 410658 796 410714 800
rect 410576 768 410714 796
rect 410576 756 410582 768
rect 410658 0 410714 768
rect 410794 756 410800 808
rect 410852 796 410858 808
rect 410930 796 410986 800
rect 410852 768 410986 796
rect 410852 756 410858 768
rect 410930 0 410986 768
rect 411070 756 411076 808
rect 411128 796 411134 808
rect 411202 796 411258 800
rect 411128 768 411258 796
rect 411128 756 411134 768
rect 411202 0 411258 768
rect 411364 592 411392 836
rect 411438 824 411444 876
rect 411496 864 411502 876
rect 495084 864 495112 904
rect 411496 836 495112 864
rect 495176 864 495204 904
rect 495176 836 497780 864
rect 411496 824 411502 836
rect 478874 756 478880 808
rect 478932 796 478938 808
rect 480018 796 480074 800
rect 478932 768 480074 796
rect 478932 756 478938 768
rect 479702 592 479708 604
rect 411364 564 479708 592
rect 479702 552 479708 564
rect 479760 552 479766 604
rect 470686 8 470692 60
rect 470744 48 470750 60
rect 479702 48 479708 60
rect 470744 20 479708 48
rect 470744 8 470750 20
rect 479702 8 479708 20
rect 479760 8 479766 60
rect 480018 0 480074 768
rect 480346 756 480352 808
rect 480404 796 480410 808
rect 481106 796 481162 800
rect 480404 768 481162 796
rect 480404 756 480410 768
rect 481106 0 481162 768
rect 481634 756 481640 808
rect 481692 796 481698 808
rect 482194 796 482250 800
rect 481692 768 482250 796
rect 481692 756 481698 768
rect 482194 0 482250 768
rect 482554 756 482560 808
rect 482612 796 482618 808
rect 483282 796 483338 800
rect 482612 768 483338 796
rect 482612 756 482618 768
rect 483282 0 483338 768
rect 484370 796 484426 800
rect 484578 796 484584 808
rect 484370 768 484584 796
rect 484370 0 484426 768
rect 484578 756 484584 768
rect 484636 756 484642 808
rect 484670 756 484676 808
rect 484728 796 484734 808
rect 485458 796 485514 800
rect 484728 768 485514 796
rect 484728 756 484734 768
rect 485458 0 485514 768
rect 485774 756 485780 808
rect 485832 796 485838 808
rect 486546 796 486602 800
rect 485832 768 486602 796
rect 485832 756 485838 768
rect 486546 0 486602 768
rect 486878 756 486884 808
rect 486936 796 486942 808
rect 487634 796 487690 800
rect 486936 768 487690 796
rect 486936 756 486942 768
rect 487634 0 487690 768
rect 488626 756 488632 808
rect 488684 796 488690 808
rect 488722 796 488778 800
rect 488684 768 488778 796
rect 488684 756 488690 768
rect 488722 0 488778 768
rect 488810 756 488816 808
rect 488868 796 488874 808
rect 489810 796 489866 800
rect 488868 768 489866 796
rect 488868 756 488874 768
rect 489810 0 489866 768
rect 489914 756 489920 808
rect 489972 796 489978 808
rect 490898 796 490954 800
rect 489972 768 490954 796
rect 489972 756 489978 768
rect 490898 0 490954 768
rect 491294 756 491300 808
rect 491352 796 491358 808
rect 491986 796 492042 800
rect 491352 768 492042 796
rect 491352 756 491358 768
rect 491986 0 492042 768
rect 492674 756 492680 808
rect 492732 796 492738 808
rect 493074 796 493130 800
rect 492732 768 493130 796
rect 492732 756 492738 768
rect 493074 0 493130 768
rect 494054 756 494060 808
rect 494112 796 494118 808
rect 494162 796 494218 800
rect 494112 768 494218 796
rect 494112 756 494118 768
rect 494162 0 494218 768
rect 494514 688 494520 740
rect 494572 728 494578 740
rect 495250 728 495306 800
rect 495618 756 495624 808
rect 495676 796 495682 808
rect 496338 796 496394 800
rect 495676 768 496394 796
rect 495676 756 495682 768
rect 494572 700 495306 728
rect 494572 688 494578 700
rect 495250 0 495306 700
rect 496338 0 496394 768
rect 496630 756 496636 808
rect 496688 796 496694 808
rect 497426 796 497482 800
rect 496688 768 497482 796
rect 497752 796 497780 836
rect 498514 796 498570 800
rect 497752 768 498570 796
rect 496688 756 496694 768
rect 497426 0 497482 768
rect 498514 0 498570 768
rect 499602 796 499658 800
rect 499758 796 499764 808
rect 499602 768 499764 796
rect 499602 0 499658 768
rect 499758 756 499764 768
rect 499816 756 499822 808
rect 500126 756 500132 808
rect 500184 796 500190 808
rect 500690 796 500746 800
rect 500184 768 500746 796
rect 500788 796 500816 904
rect 500862 824 500868 876
rect 500920 864 500926 876
rect 505066 864 505094 1040
rect 507228 864 507256 1244
rect 508332 864 508360 1312
rect 500920 836 503208 864
rect 500920 824 500926 836
rect 501778 796 501834 800
rect 500788 768 501834 796
rect 500184 756 500190 768
rect 500690 0 500746 768
rect 501778 0 501834 768
rect 502334 756 502340 808
rect 502392 796 502398 808
rect 502866 796 502922 800
rect 502392 768 502922 796
rect 503180 796 503208 836
rect 505020 836 505094 864
rect 507136 836 507256 864
rect 508240 836 508360 864
rect 505020 800 505048 836
rect 503954 796 504010 800
rect 503180 768 504010 796
rect 505020 768 505098 800
rect 502392 756 502398 768
rect 502866 0 502922 768
rect 503954 0 504010 768
rect 505042 0 505098 768
rect 505370 756 505376 808
rect 505428 796 505434 808
rect 506130 796 506186 800
rect 505428 768 506186 796
rect 507136 796 507164 836
rect 507218 796 507274 800
rect 507136 768 507274 796
rect 508240 796 508268 836
rect 508306 796 508362 800
rect 508240 768 508362 796
rect 505428 756 505434 768
rect 506130 0 506186 768
rect 507218 0 507274 768
rect 508306 0 508362 768
<< via1 >>
rect 1860 9188 1912 9240
rect 34428 9188 34480 9240
rect 52368 9188 52420 9240
rect 68928 9188 68980 9240
rect 102232 9188 102284 9240
rect 119988 9188 120040 9240
rect 136548 9188 136600 9240
rect 17868 8848 17920 8900
rect 187608 9188 187660 9240
rect 204168 9188 204220 9240
rect 222108 9188 222160 9240
rect 153108 8916 153160 8968
rect 273168 9188 273220 9240
rect 289452 9188 289504 9240
rect 340788 9188 340840 9240
rect 357256 9188 357308 9240
rect 375288 9188 375340 9240
rect 171048 8916 171100 8968
rect 238668 8916 238720 8968
rect 85488 8848 85540 8900
rect 426348 9188 426400 9240
rect 442908 9188 442960 9240
rect 306288 8916 306340 8968
rect 324228 8916 324280 8968
rect 391848 8916 391900 8968
rect 408408 8916 408460 8968
rect 255228 8848 255280 8900
rect 302884 8440 302936 8492
rect 395620 8440 395672 8492
rect 293776 8372 293828 8424
rect 387156 8372 387208 8424
rect 308404 8304 308456 8356
rect 403992 8304 404044 8356
rect 362500 7692 362552 7744
rect 408316 7692 408368 7744
rect 67574 7590 67626 7642
rect 67638 7590 67690 7642
rect 67702 7590 67754 7642
rect 67766 7590 67818 7642
rect 67830 7590 67882 7642
rect 199502 7590 199554 7642
rect 199566 7590 199618 7642
rect 199630 7590 199682 7642
rect 199694 7590 199746 7642
rect 199758 7590 199810 7642
rect 331430 7590 331482 7642
rect 331494 7590 331546 7642
rect 331558 7590 331610 7642
rect 331622 7590 331674 7642
rect 331686 7590 331738 7642
rect 463358 7590 463410 7642
rect 463422 7590 463474 7642
rect 463486 7590 463538 7642
rect 463550 7590 463602 7642
rect 463614 7590 463666 7642
rect 319628 7488 319680 7540
rect 404544 7488 404596 7540
rect 218520 7420 218572 7472
rect 306656 7420 306708 7472
rect 314752 7420 314804 7472
rect 403716 7420 403768 7472
rect 219532 7352 219584 7404
rect 300216 7352 300268 7404
rect 315948 7352 316000 7404
rect 407212 7352 407264 7404
rect 220452 7284 220504 7336
rect 301412 7284 301464 7336
rect 310704 7284 310756 7336
rect 403072 7284 403124 7336
rect 202788 7216 202840 7268
rect 296536 7216 296588 7268
rect 303436 7216 303488 7268
rect 396724 7216 396776 7268
rect 31300 7148 31352 7200
rect 125416 7148 125468 7200
rect 125876 7148 125928 7200
rect 218704 7148 218756 7200
rect 291108 7148 291160 7200
rect 385316 7148 385368 7200
rect 66914 7046 66966 7098
rect 66978 7046 67030 7098
rect 67042 7046 67094 7098
rect 67106 7046 67158 7098
rect 67170 7046 67222 7098
rect 198842 7046 198894 7098
rect 198906 7046 198958 7098
rect 198970 7046 199022 7098
rect 199034 7046 199086 7098
rect 199098 7046 199150 7098
rect 330770 7046 330822 7098
rect 330834 7046 330886 7098
rect 330898 7046 330950 7098
rect 330962 7046 331014 7098
rect 331026 7046 331078 7098
rect 462698 7046 462750 7098
rect 462762 7046 462814 7098
rect 462826 7046 462878 7098
rect 462890 7046 462942 7098
rect 462954 7046 463006 7098
rect 125140 6944 125192 6996
rect 217140 6944 217192 6996
rect 218060 6944 218112 6996
rect 314292 6944 314344 6996
rect 318340 6944 318392 6996
rect 411812 6944 411864 6996
rect 124496 6876 124548 6928
rect 218888 6876 218940 6928
rect 304724 6876 304776 6928
rect 402060 6876 402112 6928
rect 17868 6808 17920 6860
rect 19892 6808 19944 6860
rect 34428 6808 34480 6860
rect 37648 6808 37700 6860
rect 52368 6808 52420 6860
rect 53840 6808 53892 6860
rect 68928 6808 68980 6860
rect 73988 6808 74040 6860
rect 85488 6808 85540 6860
rect 92020 6808 92072 6860
rect 119988 6808 120040 6860
rect 126796 6808 126848 6860
rect 67574 6502 67626 6554
rect 67638 6502 67690 6554
rect 67702 6502 67754 6554
rect 67766 6502 67818 6554
rect 67830 6502 67882 6554
rect 199502 6502 199554 6554
rect 199566 6502 199618 6554
rect 199630 6502 199682 6554
rect 199694 6502 199746 6554
rect 199758 6502 199810 6554
rect 331430 6502 331482 6554
rect 331494 6502 331546 6554
rect 331558 6502 331610 6554
rect 331622 6502 331674 6554
rect 331686 6502 331738 6554
rect 463358 6502 463410 6554
rect 463422 6502 463474 6554
rect 463486 6502 463538 6554
rect 463550 6502 463602 6554
rect 463614 6502 463666 6554
rect 300860 6264 300912 6316
rect 351920 6264 351972 6316
rect 114192 6196 114244 6248
rect 208584 6196 208636 6248
rect 209412 6196 209464 6248
rect 306104 6196 306156 6248
rect 324228 6196 324280 6248
rect 341984 6196 342036 6248
rect 357256 6196 357308 6248
rect 380532 6196 380584 6248
rect 391848 6196 391900 6248
rect 416320 6196 416372 6248
rect 426348 6196 426400 6248
rect 442816 6196 442868 6248
rect 102232 6128 102284 6180
rect 110052 6128 110104 6180
rect 136548 6128 136600 6180
rect 145840 6128 145892 6180
rect 153108 6128 153160 6180
rect 164148 6128 164200 6180
rect 171048 6128 171100 6180
rect 179420 6128 179472 6180
rect 187608 6128 187660 6180
rect 200212 6128 200264 6180
rect 204168 6128 204220 6180
rect 217416 6128 217468 6180
rect 222108 6128 222160 6180
rect 236276 6128 236328 6180
rect 238668 6128 238720 6180
rect 254032 6128 254084 6180
rect 255228 6128 255280 6180
rect 271788 6128 271840 6180
rect 273168 6128 273220 6180
rect 288348 6128 288400 6180
rect 289452 6128 289504 6180
rect 305000 6128 305052 6180
rect 306288 6128 306340 6180
rect 326436 6128 326488 6180
rect 340788 6128 340840 6180
rect 362224 6128 362276 6180
rect 375288 6128 375340 6180
rect 398564 6128 398616 6180
rect 408408 6128 408460 6180
rect 434628 6128 434680 6180
rect 442908 6128 442960 6180
rect 470416 6128 470468 6180
rect 27712 6060 27764 6112
rect 120264 6060 120316 6112
rect 126244 6060 126296 6112
rect 219164 6060 219216 6112
rect 304816 6060 304868 6112
rect 355784 6060 355836 6112
rect 66914 5958 66966 6010
rect 66978 5958 67030 6010
rect 67042 5958 67094 6010
rect 67106 5958 67158 6010
rect 67170 5958 67222 6010
rect 198842 5958 198894 6010
rect 198906 5958 198958 6010
rect 198970 5958 199022 6010
rect 199034 5958 199086 6010
rect 199098 5958 199150 6010
rect 330770 5958 330822 6010
rect 330834 5958 330886 6010
rect 330898 5958 330950 6010
rect 330962 5958 331014 6010
rect 331026 5958 331078 6010
rect 462698 5958 462750 6010
rect 462762 5958 462814 6010
rect 462826 5958 462878 6010
rect 462890 5958 462942 6010
rect 462954 5958 463006 6010
rect 29736 5856 29788 5908
rect 123852 5856 123904 5908
rect 169208 5856 169260 5908
rect 262312 5856 262364 5908
rect 263508 5856 263560 5908
rect 340880 5856 340932 5908
rect 355140 5856 355192 5908
rect 409972 5856 410024 5908
rect 117320 5788 117372 5840
rect 207664 5788 207716 5840
rect 209044 5788 209096 5840
rect 303804 5788 303856 5840
rect 342352 5788 342404 5840
rect 407764 5788 407816 5840
rect 26424 5720 26476 5772
rect 120080 5720 120132 5772
rect 212816 5720 212868 5772
rect 308128 5720 308180 5772
rect 338028 5720 338080 5772
rect 407120 5720 407172 5772
rect 117412 5652 117464 5704
rect 208860 5652 208912 5704
rect 209596 5652 209648 5704
rect 305276 5652 305328 5704
rect 332508 5652 332560 5704
rect 406108 5652 406160 5704
rect 24584 5584 24636 5636
rect 118792 5584 118844 5636
rect 119344 5584 119396 5636
rect 213368 5584 213420 5636
rect 298652 5584 298704 5636
rect 390192 5584 390244 5636
rect 25412 5516 25464 5568
rect 118700 5516 118752 5568
rect 208400 5516 208452 5568
rect 305368 5516 305420 5568
rect 327172 5516 327224 5568
rect 421380 5516 421432 5568
rect 67574 5414 67626 5466
rect 67638 5414 67690 5466
rect 67702 5414 67754 5466
rect 67766 5414 67818 5466
rect 67830 5414 67882 5466
rect 199502 5414 199554 5466
rect 199566 5414 199618 5466
rect 199630 5414 199682 5466
rect 199694 5414 199746 5466
rect 199758 5414 199810 5466
rect 331430 5414 331482 5466
rect 331494 5414 331546 5466
rect 331558 5414 331610 5466
rect 331622 5414 331674 5466
rect 331686 5414 331738 5466
rect 463358 5414 463410 5466
rect 463422 5414 463474 5466
rect 463486 5414 463538 5466
rect 463550 5414 463602 5466
rect 463614 5414 463666 5466
rect 110788 5176 110840 5228
rect 204904 5176 204956 5228
rect 213644 5219 213696 5228
rect 213644 5185 213653 5219
rect 213653 5185 213687 5219
rect 213687 5185 213696 5219
rect 213644 5176 213696 5185
rect 218152 5176 218204 5228
rect 63592 5108 63644 5160
rect 150992 5108 151044 5160
rect 214472 5108 214524 5160
rect 220360 5108 220412 5160
rect 239036 5108 239088 5160
rect 332324 5108 332376 5160
rect 137284 5040 137336 5092
rect 230756 5040 230808 5092
rect 308496 5040 308548 5092
rect 355876 5040 355928 5092
rect 116216 5015 116268 5024
rect 116216 4981 116225 5015
rect 116225 4981 116259 5015
rect 116259 4981 116268 5015
rect 116216 4972 116268 4981
rect 116676 4972 116728 5024
rect 117504 5015 117556 5024
rect 117504 4981 117513 5015
rect 117513 4981 117547 5015
rect 117547 4981 117556 5015
rect 117504 4972 117556 4981
rect 118056 4972 118108 5024
rect 210792 4972 210844 5024
rect 211620 5015 211672 5024
rect 211620 4981 211629 5015
rect 211629 4981 211663 5015
rect 211663 4981 211672 5015
rect 211620 4972 211672 4981
rect 214288 5015 214340 5024
rect 214288 4981 214297 5015
rect 214297 4981 214331 5015
rect 214331 4981 214340 5015
rect 214288 4972 214340 4981
rect 214840 5015 214892 5024
rect 214840 4981 214849 5015
rect 214849 4981 214883 5015
rect 214883 4981 214892 5015
rect 214840 4972 214892 4981
rect 215392 5015 215444 5024
rect 215392 4981 215401 5015
rect 215401 4981 215435 5015
rect 215435 4981 215444 5015
rect 215392 4972 215444 4981
rect 216220 5015 216272 5024
rect 216220 4981 216229 5015
rect 216229 4981 216263 5015
rect 216263 4981 216272 5015
rect 216220 4972 216272 4981
rect 216864 4972 216916 5024
rect 221096 4972 221148 5024
rect 295432 4972 295484 5024
rect 306012 4972 306064 5024
rect 306748 5015 306800 5024
rect 306748 4981 306757 5015
rect 306757 4981 306791 5015
rect 306791 4981 306800 5015
rect 306748 4972 306800 4981
rect 307576 5015 307628 5024
rect 307576 4981 307585 5015
rect 307585 4981 307619 5015
rect 307619 4981 307628 5015
rect 307576 4972 307628 4981
rect 307852 4972 307904 5024
rect 308588 4972 308640 5024
rect 357440 4972 357492 5024
rect 402336 4972 402388 5024
rect 66914 4870 66966 4922
rect 66978 4870 67030 4922
rect 67042 4870 67094 4922
rect 67106 4870 67158 4922
rect 67170 4870 67222 4922
rect 198842 4870 198894 4922
rect 198906 4870 198958 4922
rect 198970 4870 199022 4922
rect 199034 4870 199086 4922
rect 199098 4870 199150 4922
rect 330770 4870 330822 4922
rect 330834 4870 330886 4922
rect 330898 4870 330950 4922
rect 330962 4870 331014 4922
rect 331026 4870 331078 4922
rect 462698 4870 462750 4922
rect 462762 4870 462814 4922
rect 462826 4870 462878 4922
rect 462890 4870 462942 4922
rect 462954 4870 463006 4922
rect 63500 4768 63552 4820
rect 156696 4768 156748 4820
rect 211528 4768 211580 4820
rect 301136 4768 301188 4820
rect 308496 4811 308548 4820
rect 308496 4777 308505 4811
rect 308505 4777 308539 4811
rect 308539 4777 308548 4811
rect 308496 4768 308548 4777
rect 350540 4768 350592 4820
rect 403808 4768 403860 4820
rect 442816 4768 442868 4820
rect 452660 4768 452712 4820
rect 131396 4700 131448 4752
rect 224960 4700 225012 4752
rect 260012 4700 260064 4752
rect 350724 4700 350776 4752
rect 353300 4700 353352 4752
rect 407304 4700 407356 4752
rect 126428 4632 126480 4684
rect 219900 4632 219952 4684
rect 221004 4632 221056 4684
rect 314016 4632 314068 4684
rect 325332 4632 325384 4684
rect 405280 4632 405332 4684
rect 28356 4564 28408 4616
rect 120632 4564 120684 4616
rect 143908 4564 143960 4616
rect 237748 4564 237800 4616
rect 307760 4564 307812 4616
rect 330024 4564 330076 4616
rect 405924 4564 405976 4616
rect 23388 4496 23440 4548
rect 58164 4496 58216 4548
rect 126612 4496 126664 4548
rect 214472 4496 214524 4548
rect 215484 4496 215536 4548
rect 217324 4496 217376 4548
rect 287428 4496 287480 4548
rect 381268 4496 381320 4548
rect 115664 4428 115716 4480
rect 116032 4471 116084 4480
rect 116032 4437 116041 4471
rect 116041 4437 116075 4471
rect 116075 4437 116084 4471
rect 116032 4428 116084 4437
rect 116584 4471 116636 4480
rect 116584 4437 116593 4471
rect 116593 4437 116627 4471
rect 116627 4437 116636 4471
rect 116584 4428 116636 4437
rect 117872 4471 117924 4480
rect 117872 4437 117881 4471
rect 117881 4437 117915 4471
rect 117915 4437 117924 4471
rect 117872 4428 117924 4437
rect 118424 4471 118476 4480
rect 118424 4437 118433 4471
rect 118433 4437 118467 4471
rect 118467 4437 118476 4471
rect 118424 4428 118476 4437
rect 118976 4471 119028 4480
rect 118976 4437 118985 4471
rect 118985 4437 119019 4471
rect 119019 4437 119028 4471
rect 118976 4428 119028 4437
rect 119528 4471 119580 4480
rect 119528 4437 119537 4471
rect 119537 4437 119571 4471
rect 119571 4437 119580 4471
rect 119528 4428 119580 4437
rect 120724 4471 120776 4480
rect 120724 4437 120733 4471
rect 120733 4437 120767 4471
rect 120767 4437 120776 4471
rect 120724 4428 120776 4437
rect 121368 4471 121420 4480
rect 121368 4437 121377 4471
rect 121377 4437 121411 4471
rect 121411 4437 121420 4471
rect 121368 4428 121420 4437
rect 122380 4428 122432 4480
rect 210424 4471 210476 4480
rect 210424 4437 210433 4471
rect 210433 4437 210467 4471
rect 210467 4437 210476 4471
rect 210424 4428 210476 4437
rect 211068 4471 211120 4480
rect 211068 4437 211077 4471
rect 211077 4437 211111 4471
rect 211111 4437 211120 4471
rect 211068 4428 211120 4437
rect 211712 4428 211764 4480
rect 212172 4428 212224 4480
rect 213184 4428 213236 4480
rect 213552 4471 213604 4480
rect 213552 4437 213561 4471
rect 213561 4437 213595 4471
rect 213595 4437 213604 4471
rect 213552 4428 213604 4437
rect 213920 4428 213972 4480
rect 215208 4428 215260 4480
rect 216772 4471 216824 4480
rect 216772 4437 216781 4471
rect 216781 4437 216815 4471
rect 216815 4437 216824 4471
rect 216772 4428 216824 4437
rect 217232 4471 217284 4480
rect 217232 4437 217241 4471
rect 217241 4437 217275 4471
rect 217275 4437 217284 4471
rect 217232 4428 217284 4437
rect 217968 4428 218020 4480
rect 220084 4428 220136 4480
rect 304172 4428 304224 4480
rect 305552 4428 305604 4480
rect 306196 4471 306248 4480
rect 306196 4437 306205 4471
rect 306205 4437 306239 4471
rect 306239 4437 306248 4471
rect 306196 4428 306248 4437
rect 306380 4428 306432 4480
rect 306840 4428 306892 4480
rect 307668 4428 307720 4480
rect 309232 4428 309284 4480
rect 309600 4471 309652 4480
rect 309600 4437 309609 4471
rect 309609 4437 309643 4471
rect 309643 4437 309652 4471
rect 309600 4428 309652 4437
rect 310428 4471 310480 4480
rect 310428 4437 310437 4471
rect 310437 4437 310471 4471
rect 310471 4437 310480 4471
rect 310428 4428 310480 4437
rect 349804 4428 349856 4480
rect 406200 4428 406252 4480
rect 67574 4326 67626 4378
rect 67638 4326 67690 4378
rect 67702 4326 67754 4378
rect 67766 4326 67818 4378
rect 67830 4326 67882 4378
rect 199502 4326 199554 4378
rect 199566 4326 199618 4378
rect 199630 4326 199682 4378
rect 199694 4326 199746 4378
rect 199758 4326 199810 4378
rect 331430 4326 331482 4378
rect 331494 4326 331546 4378
rect 331558 4326 331610 4378
rect 331622 4326 331674 4378
rect 331686 4326 331738 4378
rect 463358 4326 463410 4378
rect 463422 4326 463474 4378
rect 463486 4326 463538 4378
rect 463550 4326 463602 4378
rect 463614 4326 463666 4378
rect 22928 4224 22980 4276
rect 116308 4224 116360 4276
rect 208124 4224 208176 4276
rect 211528 4224 211580 4276
rect 20996 4156 21048 4208
rect 70400 4156 70452 4208
rect 98644 4156 98696 4208
rect 192208 4156 192260 4208
rect 203892 4156 203944 4208
rect 297364 4224 297416 4276
rect 317880 4224 317932 4276
rect 403900 4224 403952 4276
rect 220084 4156 220136 4208
rect 273076 4156 273128 4208
rect 367284 4156 367336 4208
rect 388444 4156 388496 4208
rect 481640 4156 481692 4208
rect 115756 4131 115808 4140
rect 115756 4097 115765 4131
rect 115765 4097 115799 4131
rect 115799 4097 115808 4131
rect 115756 4088 115808 4097
rect 20720 4020 20772 4072
rect 116584 4088 116636 4140
rect 118976 4088 119028 4140
rect 120356 4088 120408 4140
rect 120632 4088 120684 4140
rect 118148 4063 118200 4072
rect 118148 4029 118157 4063
rect 118157 4029 118191 4063
rect 118191 4029 118200 4063
rect 118148 4020 118200 4029
rect 121644 4063 121696 4072
rect 121644 4029 121653 4063
rect 121653 4029 121687 4063
rect 121687 4029 121696 4063
rect 121644 4020 121696 4029
rect 124496 4131 124548 4140
rect 124496 4097 124505 4131
rect 124505 4097 124539 4131
rect 124539 4097 124548 4131
rect 124496 4088 124548 4097
rect 125140 4131 125192 4140
rect 125140 4097 125149 4131
rect 125149 4097 125183 4131
rect 125183 4097 125192 4131
rect 125140 4088 125192 4097
rect 122656 4020 122708 4072
rect 123484 4063 123536 4072
rect 123484 4029 123493 4063
rect 123493 4029 123527 4063
rect 123527 4029 123536 4063
rect 123484 4020 123536 4029
rect 126520 4020 126572 4072
rect 56508 3884 56560 3936
rect 119160 3952 119212 4004
rect 208952 4088 209004 4140
rect 209044 4131 209096 4140
rect 209044 4097 209053 4131
rect 209053 4097 209087 4131
rect 209087 4097 209096 4131
rect 209044 4088 209096 4097
rect 200948 4020 201000 4072
rect 211068 4088 211120 4140
rect 212816 4131 212868 4140
rect 212816 4097 212825 4131
rect 212825 4097 212859 4131
rect 212859 4097 212868 4131
rect 212816 4088 212868 4097
rect 213368 4131 213420 4140
rect 213368 4097 213377 4131
rect 213377 4097 213411 4131
rect 213411 4097 213420 4131
rect 213368 4088 213420 4097
rect 213920 4131 213972 4140
rect 213920 4097 213929 4131
rect 213929 4097 213963 4131
rect 213963 4097 213972 4131
rect 213920 4088 213972 4097
rect 215484 4131 215536 4140
rect 215484 4097 215493 4131
rect 215493 4097 215527 4131
rect 215527 4097 215536 4131
rect 215484 4088 215536 4097
rect 216956 4088 217008 4140
rect 217324 4088 217376 4140
rect 214932 4063 214984 4072
rect 214932 4029 214941 4063
rect 214941 4029 214975 4063
rect 214975 4029 214984 4063
rect 214932 4020 214984 4029
rect 216680 4063 216732 4072
rect 216680 4029 216689 4063
rect 216689 4029 216723 4063
rect 216723 4029 216732 4063
rect 216680 4020 216732 4029
rect 116676 3884 116728 3936
rect 119344 3927 119396 3936
rect 119344 3893 119353 3927
rect 119353 3893 119387 3927
rect 119387 3893 119396 3927
rect 119344 3884 119396 3893
rect 120816 3884 120868 3936
rect 208400 3927 208452 3936
rect 208400 3893 208409 3927
rect 208409 3893 208443 3927
rect 208443 3893 208452 3927
rect 208400 3884 208452 3893
rect 208492 3884 208544 3936
rect 209596 3884 209648 3936
rect 210424 3952 210476 4004
rect 218152 4020 218204 4072
rect 304172 4063 304224 4072
rect 304172 4029 304181 4063
rect 304181 4029 304215 4063
rect 304215 4029 304224 4063
rect 304172 4020 304224 4029
rect 304816 4063 304868 4072
rect 304816 4029 304825 4063
rect 304825 4029 304859 4063
rect 304859 4029 304868 4063
rect 304816 4020 304868 4029
rect 305184 4020 305236 4072
rect 306472 4131 306524 4140
rect 306472 4097 306481 4131
rect 306481 4097 306515 4131
rect 306515 4097 306524 4131
rect 306472 4088 306524 4097
rect 306564 4088 306616 4140
rect 307668 4088 307720 4140
rect 308680 4020 308732 4072
rect 212540 3884 212592 3936
rect 216956 3884 217008 3936
rect 218060 3884 218112 3936
rect 218520 3927 218572 3936
rect 218520 3893 218529 3927
rect 218529 3893 218563 3927
rect 218563 3893 218572 3927
rect 218520 3884 218572 3893
rect 219532 3927 219584 3936
rect 219532 3893 219541 3927
rect 219541 3893 219575 3927
rect 219575 3893 219584 3927
rect 219532 3884 219584 3893
rect 219624 3884 219676 3936
rect 220452 3884 220504 3936
rect 309692 4088 309744 4140
rect 310428 4088 310480 4140
rect 310612 4088 310664 4140
rect 311440 4088 311492 4140
rect 309232 4020 309284 4072
rect 340052 4020 340104 4072
rect 310612 3952 310664 4004
rect 310704 3995 310756 4004
rect 310704 3961 310713 3995
rect 310713 3961 310747 3995
rect 310747 3961 310756 3995
rect 310704 3952 310756 3961
rect 303988 3884 304040 3936
rect 305460 3927 305512 3936
rect 305460 3893 305469 3927
rect 305469 3893 305503 3927
rect 305503 3893 305512 3927
rect 305460 3884 305512 3893
rect 306472 3884 306524 3936
rect 307024 3927 307076 3936
rect 307024 3893 307033 3927
rect 307033 3893 307067 3927
rect 307067 3893 307076 3927
rect 307024 3884 307076 3893
rect 307668 3927 307720 3936
rect 307668 3893 307677 3927
rect 307677 3893 307711 3927
rect 307711 3893 307720 3927
rect 307668 3884 307720 3893
rect 309692 3927 309744 3936
rect 309692 3893 309701 3927
rect 309701 3893 309735 3927
rect 309735 3893 309744 3927
rect 309692 3884 309744 3893
rect 309784 3884 309836 3936
rect 316776 3952 316828 4004
rect 311348 3927 311400 3936
rect 311348 3893 311357 3927
rect 311357 3893 311391 3927
rect 311391 3893 311400 3927
rect 311348 3884 311400 3893
rect 311440 3884 311492 3936
rect 401508 3952 401560 4004
rect 66914 3782 66966 3834
rect 66978 3782 67030 3834
rect 67042 3782 67094 3834
rect 67106 3782 67158 3834
rect 67170 3782 67222 3834
rect 198842 3782 198894 3834
rect 198906 3782 198958 3834
rect 198970 3782 199022 3834
rect 199034 3782 199086 3834
rect 199098 3782 199150 3834
rect 330770 3782 330822 3834
rect 330834 3782 330886 3834
rect 330898 3782 330950 3834
rect 330962 3782 331014 3834
rect 331026 3782 331078 3834
rect 462698 3782 462750 3834
rect 462762 3782 462814 3834
rect 462826 3782 462878 3834
rect 462890 3782 462942 3834
rect 462954 3782 463006 3834
rect 114100 3680 114152 3732
rect 117412 3680 117464 3732
rect 125876 3723 125928 3732
rect 125876 3689 125885 3723
rect 125885 3689 125919 3723
rect 125919 3689 125928 3723
rect 125876 3680 125928 3689
rect 126428 3723 126480 3732
rect 126428 3689 126437 3723
rect 126437 3689 126471 3723
rect 126471 3689 126480 3723
rect 126428 3680 126480 3689
rect 126520 3680 126572 3732
rect 216588 3680 216640 3732
rect 220452 3723 220504 3732
rect 220452 3689 220461 3723
rect 220461 3689 220495 3723
rect 220495 3689 220504 3723
rect 220452 3680 220504 3689
rect 220544 3680 220596 3732
rect 310704 3680 310756 3732
rect 312728 3680 312780 3732
rect 350540 3680 350592 3732
rect 353944 3680 353996 3732
rect 410248 3680 410300 3732
rect 116032 3612 116084 3664
rect 200948 3612 201000 3664
rect 108304 3544 108356 3596
rect 114928 3544 114980 3596
rect 117320 3544 117372 3596
rect 116676 3519 116728 3528
rect 116676 3485 116685 3519
rect 116685 3485 116719 3519
rect 116719 3485 116728 3519
rect 116676 3476 116728 3485
rect 118424 3544 118476 3596
rect 211712 3612 211764 3664
rect 219716 3612 219768 3664
rect 118792 3519 118844 3528
rect 118792 3485 118801 3519
rect 118801 3485 118835 3519
rect 118835 3485 118844 3519
rect 118792 3476 118844 3485
rect 119344 3519 119396 3528
rect 119344 3485 119353 3519
rect 119353 3485 119387 3519
rect 119387 3485 119396 3519
rect 119344 3476 119396 3485
rect 120080 3519 120132 3528
rect 120080 3485 120089 3519
rect 120089 3485 120123 3519
rect 120123 3485 120132 3519
rect 120080 3476 120132 3485
rect 120540 3519 120592 3528
rect 120540 3485 120549 3519
rect 120549 3485 120583 3519
rect 120583 3485 120592 3519
rect 120540 3476 120592 3485
rect 120724 3476 120776 3528
rect 22192 3408 22244 3460
rect 116124 3451 116176 3460
rect 116124 3417 116133 3451
rect 116133 3417 116167 3451
rect 116167 3417 116176 3451
rect 116124 3408 116176 3417
rect 117596 3451 117648 3460
rect 117596 3417 117605 3451
rect 117605 3417 117639 3451
rect 117639 3417 117648 3451
rect 117596 3408 117648 3417
rect 119160 3408 119212 3460
rect 119988 3408 120040 3460
rect 120632 3408 120684 3460
rect 125140 3476 125192 3528
rect 125876 3476 125928 3528
rect 121828 3451 121880 3460
rect 121828 3417 121837 3451
rect 121837 3417 121871 3451
rect 121871 3417 121880 3451
rect 121828 3408 121880 3417
rect 122380 3408 122432 3460
rect 122564 3383 122616 3392
rect 122564 3349 122573 3383
rect 122573 3349 122607 3383
rect 122607 3349 122616 3383
rect 122564 3340 122616 3349
rect 123208 3383 123260 3392
rect 123208 3349 123217 3383
rect 123217 3349 123251 3383
rect 123251 3349 123260 3383
rect 123208 3340 123260 3349
rect 123760 3451 123812 3460
rect 123760 3417 123769 3451
rect 123769 3417 123803 3451
rect 123803 3417 123812 3451
rect 123760 3408 123812 3417
rect 125048 3451 125100 3460
rect 125048 3417 125057 3451
rect 125057 3417 125091 3451
rect 125091 3417 125100 3451
rect 125048 3408 125100 3417
rect 125232 3408 125284 3460
rect 126888 3408 126940 3460
rect 208492 3476 208544 3528
rect 208860 3519 208912 3528
rect 208860 3485 208869 3519
rect 208869 3485 208903 3519
rect 208903 3485 208912 3519
rect 208860 3476 208912 3485
rect 209044 3476 209096 3528
rect 220636 3612 220688 3664
rect 308496 3612 308548 3664
rect 308680 3612 308732 3664
rect 164332 3340 164384 3392
rect 208952 3408 209004 3460
rect 212172 3519 212224 3528
rect 212172 3485 212181 3519
rect 212181 3485 212215 3519
rect 212215 3485 212224 3519
rect 212172 3476 212224 3485
rect 212908 3476 212960 3528
rect 211712 3408 211764 3460
rect 212632 3408 212684 3460
rect 214012 3451 214064 3460
rect 214012 3417 214021 3451
rect 214021 3417 214055 3451
rect 214055 3417 214064 3451
rect 214012 3408 214064 3417
rect 215208 3476 215260 3528
rect 309692 3612 309744 3664
rect 319996 3612 320048 3664
rect 351920 3612 351972 3664
rect 354036 3612 354088 3664
rect 355876 3612 355928 3664
rect 401232 3612 401284 3664
rect 214840 3408 214892 3460
rect 215852 3451 215904 3460
rect 215852 3417 215861 3451
rect 215861 3417 215895 3451
rect 215895 3417 215904 3451
rect 215852 3408 215904 3417
rect 217140 3476 217192 3528
rect 218520 3476 218572 3528
rect 218888 3519 218940 3528
rect 218888 3485 218897 3519
rect 218897 3485 218931 3519
rect 218931 3485 218940 3519
rect 218888 3476 218940 3485
rect 219624 3476 219676 3528
rect 219716 3476 219768 3528
rect 217232 3408 217284 3460
rect 219992 3408 220044 3460
rect 220176 3340 220228 3392
rect 220636 3340 220688 3392
rect 300860 3451 300912 3460
rect 300860 3417 300869 3451
rect 300869 3417 300903 3451
rect 300903 3417 300912 3451
rect 300860 3408 300912 3417
rect 259092 3340 259144 3392
rect 300308 3340 300360 3392
rect 302792 3383 302844 3392
rect 302792 3349 302801 3383
rect 302801 3349 302835 3383
rect 302835 3349 302844 3383
rect 302792 3340 302844 3349
rect 303436 3519 303488 3528
rect 303436 3485 303445 3519
rect 303445 3485 303479 3519
rect 303479 3485 303488 3519
rect 303436 3476 303488 3485
rect 303988 3519 304040 3528
rect 303988 3485 303997 3519
rect 303997 3485 304031 3519
rect 304031 3485 304040 3519
rect 303988 3476 304040 3485
rect 304816 3476 304868 3528
rect 305276 3519 305328 3528
rect 305276 3485 305285 3519
rect 305285 3485 305319 3519
rect 305319 3485 305328 3519
rect 305276 3476 305328 3485
rect 305552 3519 305604 3528
rect 305552 3485 305561 3519
rect 305561 3485 305595 3519
rect 305595 3485 305604 3519
rect 305552 3476 305604 3485
rect 306104 3476 306156 3528
rect 306472 3519 306524 3528
rect 306472 3485 306481 3519
rect 306481 3485 306515 3519
rect 306515 3485 306524 3519
rect 306472 3476 306524 3485
rect 307116 3451 307168 3460
rect 307116 3417 307125 3451
rect 307125 3417 307159 3451
rect 307159 3417 307168 3451
rect 307116 3408 307168 3417
rect 308128 3519 308180 3528
rect 308128 3485 308137 3519
rect 308137 3485 308171 3519
rect 308171 3485 308180 3519
rect 308128 3476 308180 3485
rect 309232 3476 309284 3528
rect 309600 3476 309652 3528
rect 324504 3544 324556 3596
rect 307576 3408 307628 3460
rect 309784 3408 309836 3460
rect 310888 3519 310940 3528
rect 310888 3485 310897 3519
rect 310897 3485 310931 3519
rect 310931 3485 310940 3519
rect 310888 3476 310940 3485
rect 311164 3519 311216 3528
rect 311164 3485 311173 3519
rect 311173 3485 311207 3519
rect 311207 3485 311216 3519
rect 311164 3476 311216 3485
rect 331312 3544 331364 3596
rect 336372 3544 336424 3596
rect 406476 3544 406528 3596
rect 348240 3476 348292 3528
rect 399392 3476 399444 3528
rect 307392 3340 307444 3392
rect 309416 3340 309468 3392
rect 312268 3383 312320 3392
rect 312268 3349 312277 3383
rect 312277 3349 312311 3383
rect 312311 3349 312320 3383
rect 312268 3340 312320 3349
rect 316776 3408 316828 3460
rect 344284 3408 344336 3460
rect 356980 3408 357032 3460
rect 350448 3340 350500 3392
rect 409420 3408 409472 3460
rect 357164 3383 357216 3392
rect 357164 3349 357173 3383
rect 357173 3349 357207 3383
rect 357207 3349 357216 3383
rect 357164 3340 357216 3349
rect 393596 3383 393648 3392
rect 393596 3349 393605 3383
rect 393605 3349 393639 3383
rect 393639 3349 393648 3383
rect 393596 3340 393648 3349
rect 394240 3383 394292 3392
rect 394240 3349 394249 3383
rect 394249 3349 394283 3383
rect 394283 3349 394292 3383
rect 394240 3340 394292 3349
rect 394700 3383 394752 3392
rect 394700 3349 394709 3383
rect 394709 3349 394743 3383
rect 394743 3349 394752 3383
rect 394700 3340 394752 3349
rect 396908 3340 396960 3392
rect 397368 3340 397420 3392
rect 491300 3340 491352 3392
rect 67574 3238 67626 3290
rect 67638 3238 67690 3290
rect 67702 3238 67754 3290
rect 67766 3238 67818 3290
rect 67830 3238 67882 3290
rect 199502 3238 199554 3290
rect 199566 3238 199618 3290
rect 199630 3238 199682 3290
rect 199694 3238 199746 3290
rect 199758 3238 199810 3290
rect 331430 3238 331482 3290
rect 331494 3238 331546 3290
rect 331558 3238 331610 3290
rect 331622 3238 331674 3290
rect 331686 3238 331738 3290
rect 463358 3238 463410 3290
rect 463422 3238 463474 3290
rect 463486 3238 463538 3290
rect 463550 3238 463602 3290
rect 463614 3238 463666 3290
rect 27620 3136 27672 3188
rect 116124 3136 116176 3188
rect 22100 3068 22152 3120
rect 24860 2932 24912 2984
rect 37372 2932 37424 2984
rect 31760 2864 31812 2916
rect 108304 3000 108356 3052
rect 113364 3000 113416 3052
rect 37556 2932 37608 2984
rect 116308 3111 116360 3120
rect 116308 3077 116317 3111
rect 116317 3077 116351 3111
rect 116351 3077 116360 3111
rect 116308 3068 116360 3077
rect 114100 3043 114152 3052
rect 114100 3009 114109 3043
rect 114109 3009 114143 3043
rect 114143 3009 114152 3043
rect 114100 3000 114152 3009
rect 115664 3043 115716 3052
rect 115664 3009 115673 3043
rect 115673 3009 115707 3043
rect 115707 3009 115716 3043
rect 115664 3000 115716 3009
rect 117504 3136 117556 3188
rect 210240 3136 210292 3188
rect 118700 3111 118752 3120
rect 118700 3077 118709 3111
rect 118709 3077 118743 3111
rect 118743 3077 118752 3111
rect 118700 3068 118752 3077
rect 120264 3111 120316 3120
rect 120264 3077 120273 3111
rect 120273 3077 120307 3111
rect 120307 3077 120316 3111
rect 120264 3068 120316 3077
rect 117872 3000 117924 3052
rect 117320 2932 117372 2984
rect 119528 3000 119580 3052
rect 121368 3000 121420 3052
rect 121552 2975 121604 2984
rect 121552 2941 121561 2975
rect 121561 2941 121595 2975
rect 121595 2941 121604 2975
rect 121552 2932 121604 2941
rect 29000 2796 29052 2848
rect 121736 2864 121788 2916
rect 122564 3000 122616 3052
rect 122932 2975 122984 2984
rect 122932 2941 122941 2975
rect 122941 2941 122975 2975
rect 122975 2941 122984 2975
rect 122932 2932 122984 2941
rect 123852 3111 123904 3120
rect 123852 3077 123861 3111
rect 123861 3077 123895 3111
rect 123895 3077 123904 3111
rect 123852 3068 123904 3077
rect 123208 3043 123260 3052
rect 123208 3009 123217 3043
rect 123217 3009 123251 3043
rect 123251 3009 123260 3043
rect 123208 3000 123260 3009
rect 127348 3068 127400 3120
rect 127440 3068 127492 3120
rect 124588 3000 124640 3052
rect 125232 2932 125284 2984
rect 125416 3043 125468 3052
rect 125416 3009 125425 3043
rect 125425 3009 125459 3043
rect 125459 3009 125468 3043
rect 125416 3000 125468 3009
rect 126244 3043 126296 3052
rect 126244 3009 126253 3043
rect 126253 3009 126287 3043
rect 126287 3009 126296 3043
rect 126244 3000 126296 3009
rect 145840 3043 145892 3052
rect 145840 3009 145849 3043
rect 145849 3009 145883 3043
rect 145883 3009 145892 3043
rect 145840 3000 145892 3009
rect 164332 3043 164384 3052
rect 164332 3009 164341 3043
rect 164341 3009 164375 3043
rect 164375 3009 164384 3043
rect 164332 3000 164384 3009
rect 168012 3000 168064 3052
rect 169208 2975 169260 2984
rect 169208 2941 169217 2975
rect 169217 2941 169251 2975
rect 169251 2941 169260 2975
rect 169208 2932 169260 2941
rect 201684 3000 201736 3052
rect 202788 3043 202840 3052
rect 202788 3009 202797 3043
rect 202797 3009 202831 3043
rect 202831 3009 202840 3043
rect 202788 3000 202840 3009
rect 204904 2975 204956 2984
rect 204904 2941 204913 2975
rect 204913 2941 204947 2975
rect 204947 2941 204956 2975
rect 204904 2932 204956 2941
rect 206192 3000 206244 3052
rect 206836 3000 206888 3052
rect 208124 2975 208176 2984
rect 208124 2941 208133 2975
rect 208133 2941 208167 2975
rect 208167 2941 208176 2975
rect 208124 2932 208176 2941
rect 208584 2932 208636 2984
rect 209596 3043 209648 3052
rect 209596 3009 209605 3043
rect 209605 3009 209639 3043
rect 209639 3009 209648 3043
rect 209596 3000 209648 3009
rect 210792 3043 210844 3052
rect 210792 3009 210801 3043
rect 210801 3009 210835 3043
rect 210835 3009 210844 3043
rect 210792 3000 210844 3009
rect 213184 3000 213236 3052
rect 213552 3043 213604 3052
rect 213552 3009 213561 3043
rect 213561 3009 213595 3043
rect 213595 3009 213604 3043
rect 213552 3000 213604 3009
rect 215392 3136 215444 3188
rect 220544 3136 220596 3188
rect 221096 3179 221148 3188
rect 221096 3145 221105 3179
rect 221105 3145 221139 3179
rect 221139 3145 221148 3179
rect 221096 3136 221148 3145
rect 221188 3136 221240 3188
rect 311164 3136 311216 3188
rect 314660 3136 314712 3188
rect 314752 3179 314804 3188
rect 314752 3145 314761 3179
rect 314761 3145 314795 3179
rect 314795 3145 314804 3179
rect 314752 3136 314804 3145
rect 317880 3179 317932 3188
rect 317880 3145 317889 3179
rect 317889 3145 317923 3179
rect 317923 3145 317932 3179
rect 317880 3136 317932 3145
rect 331312 3179 331364 3188
rect 331312 3145 331321 3179
rect 331321 3145 331355 3179
rect 331355 3145 331364 3179
rect 331312 3136 331364 3145
rect 340052 3179 340104 3188
rect 340052 3145 340061 3179
rect 340061 3145 340095 3179
rect 340095 3145 340104 3179
rect 340052 3136 340104 3145
rect 344284 3179 344336 3188
rect 344284 3145 344293 3179
rect 344293 3145 344327 3179
rect 344327 3145 344336 3179
rect 344284 3136 344336 3145
rect 216588 3111 216640 3120
rect 216588 3077 216597 3111
rect 216597 3077 216631 3111
rect 216631 3077 216640 3111
rect 216588 3068 216640 3077
rect 216220 3000 216272 3052
rect 217968 3000 218020 3052
rect 210240 2975 210292 2984
rect 210240 2941 210249 2975
rect 210249 2941 210283 2975
rect 210283 2941 210292 2975
rect 210240 2932 210292 2941
rect 211436 2975 211488 2984
rect 211436 2941 211445 2975
rect 211445 2941 211479 2975
rect 211479 2941 211488 2975
rect 211436 2932 211488 2941
rect 212540 2932 212592 2984
rect 37648 2839 37700 2848
rect 37648 2805 37657 2839
rect 37657 2805 37691 2839
rect 37691 2805 37700 2839
rect 37648 2796 37700 2805
rect 74724 2796 74776 2848
rect 75000 2839 75052 2848
rect 75000 2805 75009 2839
rect 75009 2805 75043 2839
rect 75043 2805 75052 2839
rect 75000 2796 75052 2805
rect 108396 2796 108448 2848
rect 112352 2796 112404 2848
rect 114192 2796 114244 2848
rect 118056 2796 118108 2848
rect 124588 2796 124640 2848
rect 126060 2864 126112 2916
rect 126888 2864 126940 2916
rect 214012 2864 214064 2916
rect 218704 3043 218756 3052
rect 218704 3009 218713 3043
rect 218713 3009 218747 3043
rect 218747 3009 218756 3043
rect 218704 3000 218756 3009
rect 219900 3111 219952 3120
rect 219900 3077 219909 3111
rect 219909 3077 219943 3111
rect 219943 3077 219952 3111
rect 219900 3068 219952 3077
rect 219532 3000 219584 3052
rect 221372 3000 221424 3052
rect 221188 2864 221240 2916
rect 254032 3043 254084 3052
rect 254032 3009 254041 3043
rect 254041 3009 254075 3043
rect 254075 3009 254084 3043
rect 254032 3000 254084 3009
rect 259092 3043 259144 3052
rect 259092 3009 259101 3043
rect 259101 3009 259135 3043
rect 259135 3009 259144 3043
rect 259092 3000 259144 3009
rect 260288 3000 260340 3052
rect 296536 3043 296588 3052
rect 296536 3009 296545 3043
rect 296545 3009 296579 3043
rect 296579 3009 296588 3043
rect 296536 3000 296588 3009
rect 297364 3043 297416 3052
rect 297364 3009 297373 3043
rect 297373 3009 297407 3043
rect 297407 3009 297416 3043
rect 297364 3000 297416 3009
rect 298652 3043 298704 3052
rect 298652 3009 298661 3043
rect 298661 3009 298695 3043
rect 298695 3009 298704 3043
rect 298652 3000 298704 3009
rect 300216 3043 300268 3052
rect 300216 3009 300225 3043
rect 300225 3009 300259 3043
rect 300259 3009 300268 3043
rect 300216 3000 300268 3009
rect 300860 3000 300912 3052
rect 301136 3043 301188 3052
rect 301136 3009 301145 3043
rect 301145 3009 301179 3043
rect 301179 3009 301188 3043
rect 301136 3000 301188 3009
rect 301228 3000 301280 3052
rect 303436 3000 303488 3052
rect 303804 2975 303856 2984
rect 303804 2941 303813 2975
rect 303813 2941 303847 2975
rect 303847 2941 303856 2975
rect 303804 2932 303856 2941
rect 304356 3043 304408 3052
rect 304356 3009 304365 3043
rect 304365 3009 304399 3043
rect 304399 3009 304408 3043
rect 304356 3000 304408 3009
rect 305368 2932 305420 2984
rect 306196 3000 306248 3052
rect 306564 3000 306616 3052
rect 306840 3000 306892 3052
rect 301228 2864 301280 2916
rect 127440 2796 127492 2848
rect 143172 2839 143224 2848
rect 143172 2805 143181 2839
rect 143181 2805 143215 2839
rect 143215 2805 143224 2839
rect 143172 2796 143224 2805
rect 152188 2796 152240 2848
rect 164792 2839 164844 2848
rect 164792 2805 164801 2839
rect 164801 2805 164835 2839
rect 164835 2805 164844 2839
rect 164792 2796 164844 2805
rect 168012 2839 168064 2848
rect 168012 2805 168021 2839
rect 168021 2805 168055 2839
rect 168055 2805 168064 2839
rect 168012 2796 168064 2805
rect 201684 2839 201736 2848
rect 201684 2805 201693 2839
rect 201693 2805 201727 2839
rect 201727 2805 201736 2839
rect 201684 2796 201736 2805
rect 206192 2796 206244 2848
rect 206836 2839 206888 2848
rect 206836 2805 206845 2839
rect 206845 2805 206879 2839
rect 206879 2805 206888 2839
rect 206836 2796 206888 2805
rect 218428 2796 218480 2848
rect 221648 2839 221700 2848
rect 221648 2805 221657 2839
rect 221657 2805 221691 2839
rect 221691 2805 221700 2839
rect 221648 2796 221700 2805
rect 247132 2796 247184 2848
rect 251732 2796 251784 2848
rect 260288 2839 260340 2848
rect 260288 2805 260297 2839
rect 260297 2805 260331 2839
rect 260331 2805 260340 2839
rect 260288 2796 260340 2805
rect 295800 2796 295852 2848
rect 299572 2839 299624 2848
rect 299572 2805 299581 2839
rect 299581 2805 299615 2839
rect 299615 2805 299624 2839
rect 299572 2796 299624 2805
rect 301136 2796 301188 2848
rect 304356 2796 304408 2848
rect 305460 2796 305512 2848
rect 306656 2864 306708 2916
rect 307392 3111 307444 3120
rect 307392 3077 307401 3111
rect 307401 3077 307435 3111
rect 307435 3077 307444 3111
rect 307392 3068 307444 3077
rect 309416 3111 309468 3120
rect 309416 3077 309425 3111
rect 309425 3077 309459 3111
rect 309459 3077 309468 3111
rect 309416 3068 309468 3077
rect 310704 3111 310756 3120
rect 310704 3077 310713 3111
rect 310713 3077 310747 3111
rect 310747 3077 310756 3111
rect 310704 3068 310756 3077
rect 307852 3000 307904 3052
rect 308588 3043 308640 3052
rect 308588 3009 308597 3043
rect 308597 3009 308631 3043
rect 308631 3009 308640 3043
rect 308588 3000 308640 3009
rect 307392 2932 307444 2984
rect 308496 2932 308548 2984
rect 312728 3043 312780 3052
rect 312728 3009 312737 3043
rect 312737 3009 312771 3043
rect 312771 3009 312780 3043
rect 312728 3000 312780 3009
rect 314016 3043 314068 3052
rect 314016 3009 314025 3043
rect 314025 3009 314059 3043
rect 314059 3009 314068 3043
rect 314016 3000 314068 3009
rect 317880 3000 317932 3052
rect 315764 2975 315816 2984
rect 315764 2941 315773 2975
rect 315773 2941 315807 2975
rect 315807 2941 315816 2975
rect 315764 2932 315816 2941
rect 323400 2932 323452 2984
rect 307760 2796 307812 2848
rect 309048 2796 309100 2848
rect 313372 2839 313424 2848
rect 313372 2805 313381 2839
rect 313381 2805 313415 2839
rect 313415 2805 313424 2839
rect 313372 2796 313424 2805
rect 342168 3068 342220 3120
rect 348240 3136 348292 3188
rect 350724 3136 350776 3188
rect 353300 3000 353352 3052
rect 353944 3179 353996 3188
rect 353944 3145 353953 3179
rect 353953 3145 353987 3179
rect 353987 3145 353996 3179
rect 353944 3136 353996 3145
rect 362224 3111 362276 3120
rect 362224 3077 362233 3111
rect 362233 3077 362267 3111
rect 362267 3077 362276 3111
rect 362224 3068 362276 3077
rect 382740 3136 382792 3188
rect 478880 3136 478932 3188
rect 411076 3068 411128 3120
rect 416320 3111 416372 3120
rect 416320 3077 416329 3111
rect 416329 3077 416363 3111
rect 416363 3077 416372 3111
rect 416320 3068 416372 3077
rect 422576 3068 422628 3120
rect 499764 3068 499816 3120
rect 340880 2932 340932 2984
rect 349804 2864 349856 2916
rect 357164 3000 357216 3052
rect 390192 3043 390244 3052
rect 390192 3009 390201 3043
rect 390201 3009 390235 3043
rect 390235 3009 390244 3043
rect 390192 3000 390244 3009
rect 390560 3043 390612 3052
rect 390560 3009 390569 3043
rect 390569 3009 390603 3043
rect 390603 3009 390612 3043
rect 390560 3000 390612 3009
rect 354036 2932 354088 2984
rect 391112 2932 391164 2984
rect 394240 3000 394292 3052
rect 394424 3043 394476 3052
rect 394424 3009 394433 3043
rect 394433 3009 394467 3043
rect 394467 3009 394476 3043
rect 394424 3000 394476 3009
rect 393596 2932 393648 2984
rect 396080 3000 396132 3052
rect 396724 3043 396776 3052
rect 396724 3009 396733 3043
rect 396733 3009 396767 3043
rect 396767 3009 396776 3043
rect 396724 3000 396776 3009
rect 401784 3000 401836 3052
rect 359556 2864 359608 2916
rect 484584 3000 484636 3052
rect 488632 2932 488684 2984
rect 470416 2907 470468 2916
rect 470416 2873 470425 2907
rect 470425 2873 470459 2907
rect 470459 2873 470468 2907
rect 470416 2864 470468 2873
rect 318984 2796 319036 2848
rect 319444 2796 319496 2848
rect 323768 2839 323820 2848
rect 323768 2805 323777 2839
rect 323777 2805 323811 2839
rect 323811 2805 323820 2839
rect 323768 2796 323820 2805
rect 324688 2796 324740 2848
rect 325148 2796 325200 2848
rect 332784 2796 332836 2848
rect 337292 2796 337344 2848
rect 337844 2796 337896 2848
rect 341524 2839 341576 2848
rect 341524 2805 341533 2839
rect 341533 2805 341567 2839
rect 341567 2805 341576 2839
rect 341524 2796 341576 2805
rect 342076 2839 342128 2848
rect 342076 2805 342085 2839
rect 342085 2805 342119 2839
rect 342119 2805 342128 2839
rect 342076 2796 342128 2805
rect 345572 2839 345624 2848
rect 345572 2805 345581 2839
rect 345581 2805 345615 2839
rect 345615 2805 345624 2839
rect 345572 2796 345624 2805
rect 346676 2839 346728 2848
rect 346676 2805 346685 2839
rect 346685 2805 346719 2839
rect 346719 2805 346728 2839
rect 346676 2796 346728 2805
rect 348424 2796 348476 2848
rect 349712 2796 349764 2848
rect 350632 2796 350684 2848
rect 352380 2796 352432 2848
rect 353668 2796 353720 2848
rect 354496 2839 354548 2848
rect 354496 2805 354505 2839
rect 354505 2805 354539 2839
rect 354539 2805 354548 2839
rect 354496 2796 354548 2805
rect 356060 2796 356112 2848
rect 358176 2839 358228 2848
rect 358176 2805 358185 2839
rect 358185 2805 358219 2839
rect 358219 2805 358228 2839
rect 358176 2796 358228 2805
rect 380900 2839 380952 2848
rect 380900 2805 380909 2839
rect 380909 2805 380943 2839
rect 380943 2805 380952 2839
rect 380900 2796 380952 2805
rect 390560 2796 390612 2848
rect 395988 2796 396040 2848
rect 396172 2839 396224 2848
rect 396172 2805 396181 2839
rect 396181 2805 396215 2839
rect 396215 2805 396224 2839
rect 396172 2796 396224 2805
rect 398932 2839 398984 2848
rect 398932 2805 398941 2839
rect 398941 2805 398975 2839
rect 398975 2805 398984 2839
rect 398932 2796 398984 2805
rect 399852 2796 399904 2848
rect 401140 2796 401192 2848
rect 408500 2839 408552 2848
rect 408500 2805 408509 2839
rect 408509 2805 408543 2839
rect 408543 2805 408552 2839
rect 408500 2796 408552 2805
rect 434996 2839 435048 2848
rect 434996 2805 435005 2839
rect 435005 2805 435039 2839
rect 435039 2805 435048 2839
rect 434996 2796 435048 2805
rect 435732 2796 435784 2848
rect 66914 2694 66966 2746
rect 66978 2694 67030 2746
rect 67042 2694 67094 2746
rect 67106 2694 67158 2746
rect 67170 2694 67222 2746
rect 198842 2694 198894 2746
rect 198906 2694 198958 2746
rect 198970 2694 199022 2746
rect 199034 2694 199086 2746
rect 199098 2694 199150 2746
rect 330770 2694 330822 2746
rect 330834 2694 330886 2746
rect 330898 2694 330950 2746
rect 330962 2694 331014 2746
rect 331026 2694 331078 2746
rect 462698 2694 462750 2746
rect 462762 2694 462814 2746
rect 462826 2694 462878 2746
rect 462890 2694 462942 2746
rect 462954 2694 463006 2746
rect 1860 2635 1912 2644
rect 1860 2601 1869 2635
rect 1869 2601 1903 2635
rect 1903 2601 1912 2635
rect 1860 2592 1912 2601
rect 19892 2635 19944 2644
rect 19892 2601 19901 2635
rect 19901 2601 19935 2635
rect 19935 2601 19944 2635
rect 19892 2592 19944 2601
rect 29184 2592 29236 2644
rect 53840 2592 53892 2644
rect 58164 2635 58216 2644
rect 58164 2601 58173 2635
rect 58173 2601 58207 2635
rect 58207 2601 58216 2635
rect 58164 2592 58216 2601
rect 56508 2524 56560 2576
rect 63592 2592 63644 2644
rect 70400 2635 70452 2644
rect 70400 2601 70409 2635
rect 70409 2601 70443 2635
rect 70443 2601 70452 2635
rect 70400 2592 70452 2601
rect 71044 2592 71096 2644
rect 73988 2635 74040 2644
rect 73988 2601 73997 2635
rect 73997 2601 74031 2635
rect 74031 2601 74040 2635
rect 73988 2592 74040 2601
rect 74540 2592 74592 2644
rect 164792 2592 164844 2644
rect 179420 2592 179472 2644
rect 211804 2592 211856 2644
rect 21916 2456 21968 2508
rect 55864 2456 55916 2508
rect 31760 2388 31812 2440
rect 35900 2388 35952 2440
rect 37648 2388 37700 2440
rect 41972 2388 42024 2440
rect 48320 2388 48372 2440
rect 24308 2320 24360 2372
rect 2596 2295 2648 2304
rect 2596 2261 2605 2295
rect 2605 2261 2639 2295
rect 2639 2261 2648 2295
rect 2596 2252 2648 2261
rect 26700 2252 26752 2304
rect 35900 2295 35952 2304
rect 35900 2261 35909 2295
rect 35909 2261 35943 2295
rect 35943 2261 35952 2295
rect 35900 2252 35952 2261
rect 36728 2363 36780 2372
rect 36728 2329 36737 2363
rect 36737 2329 36771 2363
rect 36771 2329 36780 2363
rect 36728 2320 36780 2329
rect 37924 2295 37976 2304
rect 37924 2261 37933 2295
rect 37933 2261 37967 2295
rect 37967 2261 37976 2295
rect 37924 2252 37976 2261
rect 41972 2295 42024 2304
rect 41972 2261 41981 2295
rect 41981 2261 42015 2295
rect 42015 2261 42024 2295
rect 41972 2252 42024 2261
rect 42892 2363 42944 2372
rect 42892 2329 42901 2363
rect 42901 2329 42935 2363
rect 42935 2329 42944 2363
rect 42892 2320 42944 2329
rect 54668 2431 54720 2440
rect 54668 2397 54677 2431
rect 54677 2397 54711 2431
rect 54711 2397 54720 2431
rect 54668 2388 54720 2397
rect 58164 2388 58216 2440
rect 143172 2524 143224 2576
rect 148232 2567 148284 2576
rect 148232 2533 148241 2567
rect 148241 2533 148275 2567
rect 148275 2533 148284 2567
rect 148232 2524 148284 2533
rect 58992 2363 59044 2372
rect 58992 2329 59001 2363
rect 59001 2329 59035 2363
rect 59035 2329 59044 2363
rect 58992 2320 59044 2329
rect 48320 2295 48372 2304
rect 48320 2261 48329 2295
rect 48329 2261 48363 2295
rect 48363 2261 48372 2295
rect 48320 2252 48372 2261
rect 55864 2252 55916 2304
rect 63500 2431 63552 2440
rect 63500 2397 63509 2431
rect 63509 2397 63543 2431
rect 63543 2397 63552 2431
rect 63500 2388 63552 2397
rect 70768 2320 70820 2372
rect 74540 2456 74592 2508
rect 75000 2456 75052 2508
rect 110788 2499 110840 2508
rect 71044 2431 71096 2440
rect 71044 2397 71053 2431
rect 71053 2397 71087 2431
rect 71087 2397 71096 2431
rect 71044 2388 71096 2397
rect 74632 2388 74684 2440
rect 74724 2431 74776 2440
rect 74724 2397 74733 2431
rect 74733 2397 74767 2431
rect 74767 2397 74776 2431
rect 74724 2388 74776 2397
rect 92020 2431 92072 2440
rect 92020 2397 92029 2431
rect 92029 2397 92063 2431
rect 92063 2397 92072 2431
rect 92020 2388 92072 2397
rect 75276 2363 75328 2372
rect 75276 2329 75285 2363
rect 75285 2329 75319 2363
rect 75319 2329 75328 2363
rect 75276 2320 75328 2329
rect 62580 2295 62632 2304
rect 62580 2261 62589 2295
rect 62589 2261 62623 2295
rect 62623 2261 62632 2295
rect 62580 2252 62632 2261
rect 66260 2295 66312 2304
rect 66260 2261 66269 2295
rect 66269 2261 66303 2295
rect 66303 2261 66312 2295
rect 66260 2252 66312 2261
rect 92296 2388 92348 2440
rect 98644 2431 98696 2440
rect 98644 2397 98653 2431
rect 98653 2397 98687 2431
rect 98687 2397 98696 2431
rect 98644 2388 98696 2397
rect 103888 2431 103940 2440
rect 103888 2397 103897 2431
rect 103897 2397 103931 2431
rect 103931 2397 103940 2431
rect 103888 2388 103940 2397
rect 107660 2431 107712 2440
rect 107660 2397 107669 2431
rect 107669 2397 107703 2431
rect 107703 2397 107712 2431
rect 107660 2388 107712 2397
rect 108396 2431 108448 2440
rect 108396 2397 108405 2431
rect 108405 2397 108439 2431
rect 108439 2397 108448 2431
rect 108396 2388 108448 2397
rect 110788 2465 110797 2499
rect 110797 2465 110831 2499
rect 110831 2465 110840 2499
rect 110788 2456 110840 2465
rect 113364 2456 113416 2508
rect 114928 2499 114980 2508
rect 114928 2465 114937 2499
rect 114937 2465 114971 2499
rect 114971 2465 114980 2499
rect 114928 2456 114980 2465
rect 301412 2592 301464 2644
rect 302884 2635 302936 2644
rect 302884 2601 302893 2635
rect 302893 2601 302927 2635
rect 302927 2601 302936 2635
rect 302884 2592 302936 2601
rect 304724 2635 304776 2644
rect 304724 2601 304733 2635
rect 304733 2601 304767 2635
rect 304767 2601 304776 2635
rect 304724 2592 304776 2601
rect 308404 2635 308456 2644
rect 308404 2601 308413 2635
rect 308413 2601 308447 2635
rect 308447 2601 308456 2635
rect 308404 2592 308456 2601
rect 308588 2592 308640 2644
rect 112352 2431 112404 2440
rect 112352 2397 112361 2431
rect 112361 2397 112395 2431
rect 112395 2397 112404 2431
rect 112352 2388 112404 2397
rect 114192 2388 114244 2440
rect 116216 2388 116268 2440
rect 117872 2388 117924 2440
rect 118056 2431 118108 2440
rect 118056 2397 118065 2431
rect 118065 2397 118099 2431
rect 118099 2397 118108 2431
rect 118056 2388 118108 2397
rect 120632 2431 120684 2440
rect 120632 2397 120641 2431
rect 120641 2397 120675 2431
rect 120675 2397 120684 2431
rect 120632 2388 120684 2397
rect 122380 2388 122432 2440
rect 123484 2388 123536 2440
rect 124496 2388 124548 2440
rect 96896 2363 96948 2372
rect 96896 2329 96905 2363
rect 96905 2329 96939 2363
rect 96939 2329 96948 2363
rect 96896 2320 96948 2329
rect 105084 2363 105136 2372
rect 105084 2329 105093 2363
rect 105093 2329 105127 2363
rect 105127 2329 105136 2363
rect 105084 2320 105136 2329
rect 108948 2363 109000 2372
rect 108948 2329 108957 2363
rect 108957 2329 108991 2363
rect 108991 2329 109000 2363
rect 108948 2320 109000 2329
rect 112904 2363 112956 2372
rect 112904 2329 112913 2363
rect 112913 2329 112947 2363
rect 112947 2329 112956 2363
rect 112904 2320 112956 2329
rect 117504 2363 117556 2372
rect 117504 2329 117513 2363
rect 117513 2329 117547 2363
rect 117547 2329 117556 2363
rect 117504 2320 117556 2329
rect 118700 2363 118752 2372
rect 118700 2329 118709 2363
rect 118709 2329 118743 2363
rect 118743 2329 118752 2363
rect 118700 2320 118752 2329
rect 120172 2363 120224 2372
rect 120172 2329 120181 2363
rect 120181 2329 120215 2363
rect 120215 2329 120224 2363
rect 120172 2320 120224 2329
rect 121460 2363 121512 2372
rect 121460 2329 121469 2363
rect 121469 2329 121503 2363
rect 121503 2329 121512 2363
rect 121460 2320 121512 2329
rect 122840 2363 122892 2372
rect 122840 2329 122849 2363
rect 122849 2329 122883 2363
rect 122883 2329 122892 2363
rect 122840 2320 122892 2329
rect 123852 2363 123904 2372
rect 123852 2329 123861 2363
rect 123861 2329 123895 2363
rect 123895 2329 123904 2363
rect 123852 2320 123904 2329
rect 125232 2363 125284 2372
rect 125232 2329 125241 2363
rect 125241 2329 125275 2363
rect 125275 2329 125284 2363
rect 125232 2320 125284 2329
rect 126060 2431 126112 2440
rect 126060 2397 126069 2431
rect 126069 2397 126103 2431
rect 126103 2397 126112 2431
rect 126060 2388 126112 2397
rect 126612 2431 126664 2440
rect 126612 2397 126621 2431
rect 126621 2397 126655 2431
rect 126655 2397 126664 2431
rect 126612 2388 126664 2397
rect 126428 2320 126480 2372
rect 131396 2431 131448 2440
rect 131396 2397 131405 2431
rect 131405 2397 131439 2431
rect 131439 2397 131448 2431
rect 131396 2388 131448 2397
rect 137284 2431 137336 2440
rect 137284 2397 137293 2431
rect 137293 2397 137327 2431
rect 137327 2397 137336 2431
rect 137284 2388 137336 2397
rect 143172 2388 143224 2440
rect 143908 2431 143960 2440
rect 143908 2397 143917 2431
rect 143917 2397 143951 2431
rect 143951 2397 143960 2431
rect 143908 2388 143960 2397
rect 145840 2388 145892 2440
rect 148232 2388 148284 2440
rect 152188 2431 152240 2440
rect 152188 2397 152197 2431
rect 152197 2397 152231 2431
rect 152231 2397 152240 2431
rect 152188 2388 152240 2397
rect 150992 2363 151044 2372
rect 150992 2329 151001 2363
rect 151001 2329 151035 2363
rect 151035 2329 151044 2363
rect 150992 2320 151044 2329
rect 156696 2431 156748 2440
rect 156696 2397 156705 2431
rect 156705 2397 156739 2431
rect 156739 2397 156748 2431
rect 156696 2388 156748 2397
rect 154028 2363 154080 2372
rect 154028 2329 154037 2363
rect 154037 2329 154071 2363
rect 154071 2329 154080 2363
rect 154028 2320 154080 2329
rect 157892 2363 157944 2372
rect 157892 2329 157901 2363
rect 157901 2329 157935 2363
rect 157935 2329 157944 2363
rect 157892 2320 157944 2329
rect 164332 2431 164384 2440
rect 164332 2397 164341 2431
rect 164341 2397 164375 2431
rect 164375 2397 164384 2431
rect 164332 2388 164384 2397
rect 164792 2388 164844 2440
rect 161848 2363 161900 2372
rect 161848 2329 161857 2363
rect 161857 2329 161891 2363
rect 161891 2329 161900 2363
rect 161848 2320 161900 2329
rect 165528 2363 165580 2372
rect 165528 2329 165537 2363
rect 165537 2329 165571 2363
rect 165571 2329 165580 2363
rect 165528 2320 165580 2329
rect 169024 2363 169076 2372
rect 169024 2329 169033 2363
rect 169033 2329 169067 2363
rect 169067 2329 169076 2363
rect 169024 2320 169076 2329
rect 110052 2295 110104 2304
rect 110052 2261 110061 2295
rect 110061 2261 110095 2295
rect 110095 2261 110104 2295
rect 110052 2252 110104 2261
rect 126888 2252 126940 2304
rect 128820 2295 128872 2304
rect 128820 2261 128829 2295
rect 128829 2261 128863 2295
rect 128863 2261 128872 2295
rect 128820 2252 128872 2261
rect 130200 2295 130252 2304
rect 130200 2261 130209 2295
rect 130209 2261 130243 2295
rect 130243 2261 130252 2295
rect 130200 2252 130252 2261
rect 136088 2295 136140 2304
rect 136088 2261 136097 2295
rect 136097 2261 136131 2295
rect 136131 2261 136140 2295
rect 136088 2252 136140 2261
rect 146116 2295 146168 2304
rect 146116 2261 146125 2295
rect 146125 2261 146159 2295
rect 146159 2261 146168 2295
rect 146116 2252 146168 2261
rect 152740 2295 152792 2304
rect 152740 2261 152749 2295
rect 152749 2261 152783 2295
rect 152783 2261 152792 2295
rect 152740 2252 152792 2261
rect 160468 2295 160520 2304
rect 160468 2261 160477 2295
rect 160477 2261 160511 2295
rect 160511 2261 160520 2295
rect 160468 2252 160520 2261
rect 164148 2295 164200 2304
rect 164148 2261 164157 2295
rect 164157 2261 164191 2295
rect 164191 2261 164200 2295
rect 164148 2252 164200 2261
rect 192208 2431 192260 2440
rect 192208 2397 192217 2431
rect 192217 2397 192251 2431
rect 192251 2397 192260 2431
rect 192208 2388 192260 2397
rect 170772 2295 170824 2304
rect 170772 2261 170781 2295
rect 170781 2261 170815 2295
rect 170815 2261 170824 2295
rect 170772 2252 170824 2261
rect 182916 2295 182968 2304
rect 182916 2261 182925 2295
rect 182925 2261 182959 2295
rect 182959 2261 182968 2295
rect 182916 2252 182968 2261
rect 200212 2431 200264 2440
rect 200212 2397 200221 2431
rect 200221 2397 200255 2431
rect 200255 2397 200264 2431
rect 200212 2388 200264 2397
rect 199384 2320 199436 2372
rect 203892 2431 203944 2440
rect 203892 2397 203901 2431
rect 203901 2397 203935 2431
rect 203935 2397 203944 2431
rect 203892 2388 203944 2397
rect 207664 2431 207716 2440
rect 207664 2397 207673 2431
rect 207673 2397 207707 2431
rect 207707 2397 207716 2431
rect 207664 2388 207716 2397
rect 208400 2388 208452 2440
rect 209412 2431 209464 2440
rect 206100 2363 206152 2372
rect 206100 2329 206109 2363
rect 206109 2329 206143 2363
rect 206143 2329 206152 2363
rect 206100 2320 206152 2329
rect 209412 2397 209421 2431
rect 209421 2397 209455 2431
rect 209455 2397 209464 2431
rect 209412 2388 209464 2397
rect 208860 2363 208912 2372
rect 208860 2329 208869 2363
rect 208869 2329 208903 2363
rect 208903 2329 208912 2363
rect 208860 2320 208912 2329
rect 210240 2363 210292 2372
rect 210240 2329 210249 2363
rect 210249 2329 210283 2363
rect 210283 2329 210292 2363
rect 210240 2320 210292 2329
rect 211528 2431 211580 2440
rect 211528 2397 211537 2431
rect 211537 2397 211571 2431
rect 211571 2397 211580 2431
rect 211528 2388 211580 2397
rect 211804 2499 211856 2508
rect 211804 2465 211813 2499
rect 211813 2465 211847 2499
rect 211847 2465 211856 2499
rect 211804 2456 211856 2465
rect 214932 2456 214984 2508
rect 216864 2456 216916 2508
rect 219164 2499 219216 2508
rect 219164 2465 219173 2499
rect 219173 2465 219207 2499
rect 219207 2465 219216 2499
rect 219164 2456 219216 2465
rect 213644 2388 213696 2440
rect 214288 2388 214340 2440
rect 216680 2388 216732 2440
rect 216772 2388 216824 2440
rect 211620 2320 211672 2372
rect 212448 2320 212500 2372
rect 212816 2363 212868 2372
rect 212816 2329 212825 2363
rect 212825 2329 212859 2363
rect 212859 2329 212868 2363
rect 212816 2320 212868 2329
rect 214012 2363 214064 2372
rect 214012 2329 214021 2363
rect 214021 2329 214055 2363
rect 214055 2329 214064 2363
rect 214012 2320 214064 2329
rect 215392 2363 215444 2372
rect 215392 2329 215401 2363
rect 215401 2329 215435 2363
rect 215435 2329 215444 2363
rect 215392 2320 215444 2329
rect 216588 2363 216640 2372
rect 216588 2329 216597 2363
rect 216597 2329 216631 2363
rect 216631 2329 216640 2363
rect 216588 2320 216640 2329
rect 193588 2295 193640 2304
rect 193588 2261 193597 2295
rect 193597 2261 193631 2295
rect 193631 2261 193640 2295
rect 193588 2252 193640 2261
rect 197912 2295 197964 2304
rect 197912 2261 197921 2295
rect 197921 2261 197955 2295
rect 197955 2261 197964 2295
rect 197912 2252 197964 2261
rect 200396 2295 200448 2304
rect 200396 2261 200405 2295
rect 200405 2261 200439 2295
rect 200439 2261 200448 2295
rect 200396 2252 200448 2261
rect 202696 2295 202748 2304
rect 202696 2261 202705 2295
rect 202705 2261 202739 2295
rect 202739 2261 202748 2295
rect 202696 2252 202748 2261
rect 204904 2295 204956 2304
rect 204904 2261 204913 2295
rect 204913 2261 204947 2295
rect 204947 2261 204956 2295
rect 204904 2252 204956 2261
rect 217968 2252 218020 2304
rect 218428 2431 218480 2440
rect 218428 2397 218437 2431
rect 218437 2397 218471 2431
rect 218471 2397 218480 2431
rect 218428 2388 218480 2397
rect 221648 2456 221700 2508
rect 220360 2388 220412 2440
rect 221004 2431 221056 2440
rect 221004 2397 221013 2431
rect 221013 2397 221047 2431
rect 221047 2397 221056 2431
rect 221004 2388 221056 2397
rect 223028 2363 223080 2372
rect 223028 2329 223037 2363
rect 223037 2329 223071 2363
rect 223071 2329 223080 2363
rect 223028 2320 223080 2329
rect 224960 2431 225012 2440
rect 224960 2397 224969 2431
rect 224969 2397 225003 2431
rect 225003 2397 225012 2431
rect 224960 2388 225012 2397
rect 230756 2431 230808 2440
rect 230756 2397 230765 2431
rect 230765 2397 230799 2431
rect 230799 2397 230808 2431
rect 230756 2388 230808 2397
rect 226156 2363 226208 2372
rect 226156 2329 226165 2363
rect 226165 2329 226199 2363
rect 226199 2329 226208 2363
rect 226156 2320 226208 2329
rect 231952 2363 232004 2372
rect 231952 2329 231961 2363
rect 231961 2329 231995 2363
rect 231995 2329 232004 2363
rect 231952 2320 232004 2329
rect 237748 2431 237800 2440
rect 237748 2397 237757 2431
rect 237757 2397 237791 2431
rect 237791 2397 237800 2431
rect 237748 2388 237800 2397
rect 239036 2431 239088 2440
rect 239036 2397 239045 2431
rect 239045 2397 239079 2431
rect 239079 2397 239088 2431
rect 239036 2388 239088 2397
rect 247132 2431 247184 2440
rect 247132 2397 247141 2431
rect 247141 2397 247175 2431
rect 247175 2397 247184 2431
rect 247132 2388 247184 2397
rect 244188 2363 244240 2372
rect 244188 2329 244197 2363
rect 244197 2329 244231 2363
rect 244231 2329 244240 2363
rect 244188 2320 244240 2329
rect 246304 2363 246356 2372
rect 246304 2329 246313 2363
rect 246313 2329 246347 2363
rect 246347 2329 246356 2363
rect 246304 2320 246356 2329
rect 221372 2252 221424 2304
rect 224224 2295 224276 2304
rect 224224 2261 224233 2295
rect 224233 2261 224267 2295
rect 224267 2261 224276 2295
rect 224224 2252 224276 2261
rect 236276 2295 236328 2304
rect 236276 2261 236285 2295
rect 236285 2261 236319 2295
rect 236319 2261 236328 2295
rect 236276 2252 236328 2261
rect 237012 2295 237064 2304
rect 237012 2261 237021 2295
rect 237021 2261 237055 2295
rect 237055 2261 237064 2295
rect 237012 2252 237064 2261
rect 248052 2295 248104 2304
rect 248052 2261 248061 2295
rect 248061 2261 248095 2295
rect 248095 2261 248104 2295
rect 291108 2499 291160 2508
rect 251732 2431 251784 2440
rect 251732 2397 251741 2431
rect 251741 2397 251775 2431
rect 251775 2397 251784 2431
rect 251732 2388 251784 2397
rect 254032 2388 254084 2440
rect 255780 2388 255832 2440
rect 248052 2252 248104 2261
rect 254308 2295 254360 2304
rect 254308 2261 254317 2295
rect 254317 2261 254351 2295
rect 254351 2261 254360 2295
rect 254308 2252 254360 2261
rect 255780 2295 255832 2304
rect 255780 2261 255789 2295
rect 255789 2261 255823 2295
rect 255823 2261 255832 2295
rect 255780 2252 255832 2261
rect 257068 2363 257120 2372
rect 257068 2329 257077 2363
rect 257077 2329 257111 2363
rect 257111 2329 257120 2363
rect 257068 2320 257120 2329
rect 260012 2431 260064 2440
rect 260012 2397 260021 2431
rect 260021 2397 260055 2431
rect 260055 2397 260064 2431
rect 260012 2388 260064 2397
rect 262312 2431 262364 2440
rect 262312 2397 262321 2431
rect 262321 2397 262355 2431
rect 262355 2397 262364 2431
rect 262312 2388 262364 2397
rect 263508 2431 263560 2440
rect 263508 2397 263517 2431
rect 263517 2397 263551 2431
rect 263551 2397 263560 2431
rect 263508 2388 263560 2397
rect 273076 2431 273128 2440
rect 264336 2363 264388 2372
rect 264336 2329 264345 2363
rect 264345 2329 264379 2363
rect 264379 2329 264388 2363
rect 264336 2320 264388 2329
rect 258264 2252 258316 2304
rect 258356 2295 258408 2304
rect 258356 2261 258365 2295
rect 258365 2261 258399 2295
rect 258399 2261 258408 2295
rect 258356 2252 258408 2261
rect 273076 2397 273085 2431
rect 273085 2397 273119 2431
rect 273119 2397 273128 2431
rect 273076 2388 273128 2397
rect 277124 2363 277176 2372
rect 277124 2329 277133 2363
rect 277133 2329 277167 2363
rect 277167 2329 277176 2363
rect 277124 2320 277176 2329
rect 287428 2431 287480 2440
rect 287428 2397 287437 2431
rect 287437 2397 287471 2431
rect 287471 2397 287480 2431
rect 287428 2388 287480 2397
rect 285956 2363 286008 2372
rect 285956 2329 285965 2363
rect 285965 2329 285999 2363
rect 285999 2329 286008 2363
rect 285956 2320 286008 2329
rect 291108 2465 291117 2499
rect 291117 2465 291151 2499
rect 291151 2465 291160 2499
rect 291108 2456 291160 2465
rect 293776 2499 293828 2508
rect 293776 2465 293785 2499
rect 293785 2465 293819 2499
rect 293819 2465 293828 2499
rect 293776 2456 293828 2465
rect 292580 2388 292632 2440
rect 295432 2431 295484 2440
rect 295432 2397 295441 2431
rect 295441 2397 295475 2431
rect 295475 2397 295484 2431
rect 295432 2388 295484 2397
rect 296536 2388 296588 2440
rect 296996 2431 297048 2440
rect 296996 2397 297005 2431
rect 297005 2397 297039 2431
rect 297039 2397 297048 2431
rect 296996 2388 297048 2397
rect 298652 2388 298704 2440
rect 299572 2431 299624 2440
rect 299572 2397 299581 2431
rect 299581 2397 299615 2431
rect 299615 2397 299624 2431
rect 299572 2388 299624 2397
rect 300308 2431 300360 2440
rect 300308 2397 300317 2431
rect 300317 2397 300351 2431
rect 300351 2397 300360 2431
rect 300308 2388 300360 2397
rect 295800 2363 295852 2372
rect 295800 2329 295809 2363
rect 295809 2329 295843 2363
rect 295843 2329 295852 2363
rect 295800 2320 295852 2329
rect 299020 2363 299072 2372
rect 299020 2329 299029 2363
rect 299029 2329 299063 2363
rect 299063 2329 299072 2363
rect 299020 2320 299072 2329
rect 300768 2363 300820 2372
rect 300768 2329 300777 2363
rect 300777 2329 300811 2363
rect 300811 2329 300820 2363
rect 300768 2320 300820 2329
rect 302792 2524 302844 2576
rect 302792 2388 302844 2440
rect 309048 2524 309100 2576
rect 305460 2456 305512 2508
rect 310888 2456 310940 2508
rect 304172 2388 304224 2440
rect 306012 2431 306064 2440
rect 306012 2397 306021 2431
rect 306021 2397 306055 2431
rect 306055 2397 306064 2431
rect 306012 2388 306064 2397
rect 306748 2431 306800 2440
rect 306748 2397 306757 2431
rect 306757 2397 306791 2431
rect 306791 2397 306800 2431
rect 306748 2388 306800 2397
rect 310612 2388 310664 2440
rect 310704 2431 310756 2440
rect 310704 2397 310713 2431
rect 310713 2397 310747 2431
rect 310747 2397 310756 2431
rect 310704 2388 310756 2397
rect 312268 2524 312320 2576
rect 313188 2524 313240 2576
rect 314292 2592 314344 2644
rect 318340 2635 318392 2644
rect 318340 2601 318349 2635
rect 318349 2601 318383 2635
rect 318383 2601 318392 2635
rect 318340 2592 318392 2601
rect 319628 2635 319680 2644
rect 319628 2601 319637 2635
rect 319637 2601 319671 2635
rect 319671 2601 319680 2635
rect 319628 2592 319680 2601
rect 319720 2592 319772 2644
rect 350448 2635 350500 2644
rect 350448 2601 350457 2635
rect 350457 2601 350491 2635
rect 350491 2601 350500 2635
rect 350448 2592 350500 2601
rect 355140 2635 355192 2644
rect 355140 2601 355149 2635
rect 355149 2601 355183 2635
rect 355183 2601 355192 2635
rect 355140 2592 355192 2601
rect 355784 2592 355836 2644
rect 359556 2635 359608 2644
rect 359556 2601 359565 2635
rect 359565 2601 359599 2635
rect 359599 2601 359608 2635
rect 359556 2592 359608 2601
rect 362500 2635 362552 2644
rect 362500 2601 362509 2635
rect 362509 2601 362543 2635
rect 362543 2601 362552 2635
rect 362500 2592 362552 2601
rect 380532 2635 380584 2644
rect 380532 2601 380541 2635
rect 380541 2601 380575 2635
rect 380575 2601 380584 2635
rect 380532 2592 380584 2601
rect 382740 2635 382792 2644
rect 382740 2601 382749 2635
rect 382749 2601 382783 2635
rect 382783 2601 382792 2635
rect 382740 2592 382792 2601
rect 387156 2635 387208 2644
rect 387156 2601 387165 2635
rect 387165 2601 387199 2635
rect 387199 2601 387208 2635
rect 387156 2592 387208 2601
rect 395620 2635 395672 2644
rect 395620 2601 395629 2635
rect 395629 2601 395663 2635
rect 395663 2601 395672 2635
rect 395620 2592 395672 2601
rect 398564 2635 398616 2644
rect 398564 2601 398573 2635
rect 398573 2601 398607 2635
rect 398607 2601 398616 2635
rect 398564 2592 398616 2601
rect 325240 2524 325292 2576
rect 325332 2567 325384 2576
rect 325332 2533 325341 2567
rect 325341 2533 325375 2567
rect 325375 2533 325384 2567
rect 325332 2524 325384 2533
rect 325424 2524 325476 2576
rect 342076 2524 342128 2576
rect 407856 2592 407908 2644
rect 408500 2592 408552 2644
rect 492680 2592 492732 2644
rect 311164 2456 311216 2508
rect 303988 2363 304040 2372
rect 303988 2329 303997 2363
rect 303997 2329 304031 2363
rect 304031 2329 304040 2363
rect 303988 2320 304040 2329
rect 305460 2363 305512 2372
rect 305460 2329 305469 2363
rect 305469 2329 305503 2363
rect 305503 2329 305512 2363
rect 305460 2320 305512 2329
rect 307300 2363 307352 2372
rect 307300 2329 307309 2363
rect 307309 2329 307343 2363
rect 307343 2329 307352 2363
rect 307300 2320 307352 2329
rect 265716 2295 265768 2304
rect 265716 2261 265725 2295
rect 265725 2261 265759 2295
rect 265759 2261 265768 2295
rect 265716 2252 265768 2261
rect 271788 2252 271840 2304
rect 278320 2295 278372 2304
rect 278320 2261 278329 2295
rect 278329 2261 278363 2295
rect 278363 2261 278372 2295
rect 278320 2252 278372 2261
rect 288348 2252 288400 2304
rect 292580 2295 292632 2304
rect 292580 2261 292589 2295
rect 292589 2261 292623 2295
rect 292623 2261 292632 2295
rect 292580 2252 292632 2261
rect 305000 2252 305052 2304
rect 309232 2363 309284 2372
rect 309232 2329 309241 2363
rect 309241 2329 309275 2363
rect 309275 2329 309284 2363
rect 309232 2320 309284 2329
rect 315948 2388 316000 2440
rect 316592 2388 316644 2440
rect 310612 2252 310664 2304
rect 311348 2252 311400 2304
rect 311532 2295 311584 2304
rect 311532 2261 311541 2295
rect 311541 2261 311575 2295
rect 311575 2261 311584 2295
rect 311532 2252 311584 2261
rect 313280 2363 313332 2372
rect 313280 2329 313289 2363
rect 313289 2329 313323 2363
rect 313323 2329 313332 2363
rect 313280 2320 313332 2329
rect 315764 2320 315816 2372
rect 317052 2363 317104 2372
rect 317052 2329 317061 2363
rect 317061 2329 317095 2363
rect 317095 2329 317104 2363
rect 317052 2320 317104 2329
rect 318340 2388 318392 2440
rect 318984 2431 319036 2440
rect 318984 2397 318993 2431
rect 318993 2397 319027 2431
rect 319027 2397 319036 2431
rect 318984 2388 319036 2397
rect 319444 2431 319496 2440
rect 319444 2397 319453 2431
rect 319453 2397 319487 2431
rect 319487 2397 319496 2431
rect 319444 2388 319496 2397
rect 319720 2320 319772 2372
rect 313372 2252 313424 2304
rect 314752 2252 314804 2304
rect 323400 2295 323452 2304
rect 323400 2261 323409 2295
rect 323409 2261 323443 2295
rect 323443 2261 323452 2295
rect 323400 2252 323452 2261
rect 324688 2431 324740 2440
rect 324688 2397 324697 2431
rect 324697 2397 324731 2431
rect 324731 2397 324740 2431
rect 324688 2388 324740 2397
rect 325148 2431 325200 2440
rect 325148 2397 325157 2431
rect 325157 2397 325191 2431
rect 325191 2397 325200 2431
rect 325148 2388 325200 2397
rect 327172 2431 327224 2440
rect 327172 2397 327181 2431
rect 327181 2397 327215 2431
rect 327215 2397 327224 2431
rect 327172 2388 327224 2397
rect 330024 2431 330076 2440
rect 330024 2397 330033 2431
rect 330033 2397 330067 2431
rect 330067 2397 330076 2431
rect 330024 2388 330076 2397
rect 331220 2363 331272 2372
rect 331220 2329 331229 2363
rect 331229 2329 331263 2363
rect 331263 2329 331272 2363
rect 331220 2320 331272 2329
rect 332324 2431 332376 2440
rect 332324 2397 332333 2431
rect 332333 2397 332367 2431
rect 332367 2397 332376 2431
rect 332324 2388 332376 2397
rect 336372 2431 336424 2440
rect 336372 2397 336381 2431
rect 336381 2397 336415 2431
rect 336415 2397 336424 2431
rect 336372 2388 336424 2397
rect 337844 2431 337896 2440
rect 337844 2397 337853 2431
rect 337853 2397 337887 2431
rect 337887 2397 337896 2431
rect 337844 2388 337896 2397
rect 341524 2388 341576 2440
rect 342076 2388 342128 2440
rect 342168 2431 342220 2440
rect 342168 2397 342177 2431
rect 342177 2397 342211 2431
rect 342211 2397 342220 2431
rect 342168 2388 342220 2397
rect 345572 2388 345624 2440
rect 346216 2388 346268 2440
rect 346584 2431 346636 2440
rect 346584 2397 346593 2431
rect 346593 2397 346627 2431
rect 346627 2397 346636 2431
rect 346584 2388 346636 2397
rect 350632 2388 350684 2440
rect 353668 2431 353720 2440
rect 353668 2397 353677 2431
rect 353677 2397 353711 2431
rect 353711 2397 353720 2431
rect 353668 2388 353720 2397
rect 356060 2431 356112 2440
rect 356060 2397 356069 2431
rect 356069 2397 356103 2431
rect 356103 2397 356112 2431
rect 356060 2388 356112 2397
rect 332784 2320 332836 2372
rect 335268 2363 335320 2372
rect 335268 2329 335277 2363
rect 335277 2329 335311 2363
rect 335311 2329 335320 2363
rect 335268 2320 335320 2329
rect 337292 2363 337344 2372
rect 337292 2329 337301 2363
rect 337301 2329 337335 2363
rect 337335 2329 337344 2363
rect 337292 2320 337344 2329
rect 339960 2363 340012 2372
rect 339960 2329 339969 2363
rect 339969 2329 340003 2363
rect 340003 2329 340012 2363
rect 339960 2320 340012 2329
rect 341984 2320 342036 2372
rect 323768 2252 323820 2304
rect 324504 2295 324556 2304
rect 324504 2261 324513 2295
rect 324513 2261 324547 2295
rect 324547 2261 324556 2295
rect 324504 2252 324556 2261
rect 326436 2295 326488 2304
rect 326436 2261 326445 2295
rect 326445 2261 326479 2295
rect 326479 2261 326488 2295
rect 326436 2252 326488 2261
rect 329288 2295 329340 2304
rect 329288 2261 329297 2295
rect 329297 2261 329331 2295
rect 329331 2261 329340 2295
rect 329288 2252 329340 2261
rect 332508 2295 332560 2304
rect 332508 2261 332517 2295
rect 332517 2261 332551 2295
rect 332551 2261 332560 2295
rect 332508 2252 332560 2261
rect 337200 2295 337252 2304
rect 337200 2261 337209 2295
rect 337209 2261 337243 2295
rect 337243 2261 337252 2295
rect 337200 2252 337252 2261
rect 338028 2295 338080 2304
rect 338028 2261 338037 2295
rect 338037 2261 338071 2295
rect 338071 2261 338080 2295
rect 338028 2252 338080 2261
rect 342352 2295 342404 2304
rect 342352 2261 342361 2295
rect 342361 2261 342395 2295
rect 342395 2261 342404 2295
rect 342352 2252 342404 2261
rect 346676 2320 346728 2372
rect 348424 2363 348476 2372
rect 348424 2329 348433 2363
rect 348433 2329 348467 2363
rect 348467 2329 348476 2363
rect 348424 2320 348476 2329
rect 349712 2363 349764 2372
rect 349712 2329 349721 2363
rect 349721 2329 349755 2363
rect 349755 2329 349764 2363
rect 349712 2320 349764 2329
rect 352380 2363 352432 2372
rect 352380 2329 352389 2363
rect 352389 2329 352423 2363
rect 352423 2329 352432 2363
rect 352380 2320 352432 2329
rect 353300 2363 353352 2372
rect 353300 2329 353309 2363
rect 353309 2329 353343 2363
rect 353343 2329 353352 2363
rect 353300 2320 353352 2329
rect 355140 2320 355192 2372
rect 345664 2295 345716 2304
rect 345664 2261 345673 2295
rect 345673 2261 345707 2295
rect 345707 2261 345716 2295
rect 345664 2252 345716 2261
rect 346768 2295 346820 2304
rect 346768 2261 346777 2295
rect 346777 2261 346811 2295
rect 346811 2261 346820 2295
rect 346768 2252 346820 2261
rect 349620 2295 349672 2304
rect 349620 2261 349629 2295
rect 349629 2261 349663 2295
rect 349663 2261 349672 2295
rect 349620 2252 349672 2261
rect 352288 2295 352340 2304
rect 352288 2261 352297 2295
rect 352297 2261 352331 2295
rect 352331 2261 352340 2295
rect 352288 2252 352340 2261
rect 354404 2295 354456 2304
rect 354404 2261 354413 2295
rect 354413 2261 354447 2295
rect 354447 2261 354456 2295
rect 354404 2252 354456 2261
rect 367284 2499 367336 2508
rect 367284 2465 367293 2499
rect 367293 2465 367327 2499
rect 367327 2465 367336 2499
rect 367284 2456 367336 2465
rect 358176 2388 358228 2440
rect 359556 2388 359608 2440
rect 362224 2388 362276 2440
rect 357900 2363 357952 2372
rect 357900 2329 357909 2363
rect 357909 2329 357943 2363
rect 357943 2329 357952 2363
rect 357900 2320 357952 2329
rect 371148 2363 371200 2372
rect 371148 2329 371157 2363
rect 371157 2329 371191 2363
rect 371191 2329 371200 2363
rect 371148 2320 371200 2329
rect 380900 2388 380952 2440
rect 381268 2431 381320 2440
rect 381268 2397 381277 2431
rect 381277 2397 381311 2431
rect 381311 2397 381320 2431
rect 381268 2388 381320 2397
rect 382740 2388 382792 2440
rect 385316 2499 385368 2508
rect 385316 2465 385325 2499
rect 385325 2465 385359 2499
rect 385359 2465 385368 2499
rect 385316 2456 385368 2465
rect 403992 2499 404044 2508
rect 403992 2465 404001 2499
rect 404001 2465 404035 2499
rect 404035 2465 404044 2499
rect 403992 2456 404044 2465
rect 372436 2363 372488 2372
rect 372436 2329 372445 2363
rect 372445 2329 372479 2363
rect 372479 2329 372488 2363
rect 372436 2320 372488 2329
rect 387156 2388 387208 2440
rect 388444 2431 388496 2440
rect 388444 2397 388453 2431
rect 388453 2397 388487 2431
rect 388487 2397 388496 2431
rect 388444 2388 388496 2397
rect 389272 2363 389324 2372
rect 389272 2329 389281 2363
rect 389281 2329 389315 2363
rect 389315 2329 389324 2363
rect 389272 2320 389324 2329
rect 391112 2431 391164 2440
rect 391112 2397 391121 2431
rect 391121 2397 391155 2431
rect 391155 2397 391164 2431
rect 391112 2388 391164 2397
rect 394700 2388 394752 2440
rect 396908 2431 396960 2440
rect 396908 2397 396917 2431
rect 396917 2397 396951 2431
rect 396951 2397 396960 2431
rect 396908 2388 396960 2397
rect 397368 2431 397420 2440
rect 397368 2397 397377 2431
rect 397377 2397 397411 2431
rect 397411 2397 397420 2431
rect 397368 2388 397420 2397
rect 398932 2388 398984 2440
rect 391664 2363 391716 2372
rect 391664 2329 391673 2363
rect 391673 2329 391707 2363
rect 391707 2329 391716 2363
rect 391664 2320 391716 2329
rect 393872 2363 393924 2372
rect 393872 2329 393881 2363
rect 393881 2329 393915 2363
rect 393915 2329 393924 2363
rect 393872 2320 393924 2329
rect 396172 2320 396224 2372
rect 386512 2295 386564 2304
rect 386512 2261 386521 2295
rect 386521 2261 386555 2295
rect 386555 2261 386564 2295
rect 386512 2252 386564 2261
rect 390468 2295 390520 2304
rect 390468 2261 390477 2295
rect 390477 2261 390511 2295
rect 390511 2261 390520 2295
rect 390468 2252 390520 2261
rect 399300 2363 399352 2372
rect 399300 2329 399309 2363
rect 399309 2329 399343 2363
rect 399343 2329 399352 2363
rect 399300 2320 399352 2329
rect 399852 2431 399904 2440
rect 399852 2397 399861 2431
rect 399861 2397 399895 2431
rect 399895 2397 399904 2431
rect 399852 2388 399904 2397
rect 401140 2431 401192 2440
rect 401140 2397 401149 2431
rect 401149 2397 401183 2431
rect 401183 2397 401192 2431
rect 401140 2388 401192 2397
rect 407212 2499 407264 2508
rect 407212 2465 407221 2499
rect 407221 2465 407255 2499
rect 407255 2465 407264 2499
rect 407212 2456 407264 2465
rect 408500 2456 408552 2508
rect 411812 2499 411864 2508
rect 411812 2465 411821 2499
rect 411821 2465 411855 2499
rect 411855 2465 411864 2499
rect 411812 2456 411864 2465
rect 422576 2567 422628 2576
rect 422576 2533 422585 2567
rect 422585 2533 422619 2567
rect 422619 2533 422628 2567
rect 422576 2524 422628 2533
rect 434628 2567 434680 2576
rect 434628 2533 434637 2567
rect 434637 2533 434671 2567
rect 434671 2533 434680 2567
rect 434628 2524 434680 2533
rect 434996 2524 435048 2576
rect 505376 2524 505428 2576
rect 408316 2388 408368 2440
rect 400864 2252 400916 2304
rect 401508 2363 401560 2372
rect 401508 2329 401517 2363
rect 401517 2329 401551 2363
rect 401551 2329 401560 2363
rect 401508 2320 401560 2329
rect 405188 2363 405240 2372
rect 405188 2329 405197 2363
rect 405197 2329 405231 2363
rect 405231 2329 405240 2363
rect 405188 2320 405240 2329
rect 409696 2320 409748 2372
rect 407672 2252 407724 2304
rect 416320 2388 416372 2440
rect 421380 2431 421432 2440
rect 421380 2397 421389 2431
rect 421389 2397 421423 2431
rect 421423 2397 421432 2431
rect 421380 2388 421432 2397
rect 422576 2388 422628 2440
rect 425152 2363 425204 2372
rect 425152 2329 425161 2363
rect 425161 2329 425195 2363
rect 425195 2329 425204 2363
rect 425152 2320 425204 2329
rect 434996 2388 435048 2440
rect 435732 2431 435784 2440
rect 435732 2397 435741 2431
rect 435741 2397 435775 2431
rect 435775 2397 435784 2431
rect 435732 2388 435784 2397
rect 435456 2363 435508 2372
rect 435456 2329 435465 2363
rect 435465 2329 435499 2363
rect 435499 2329 435508 2363
rect 435456 2320 435508 2329
rect 439412 2363 439464 2372
rect 439412 2329 439421 2363
rect 439421 2329 439455 2363
rect 439455 2329 439464 2363
rect 439412 2320 439464 2329
rect 447784 2363 447836 2372
rect 447784 2329 447793 2363
rect 447793 2329 447827 2363
rect 447827 2329 447836 2363
rect 447784 2320 447836 2329
rect 465724 2431 465776 2440
rect 465724 2397 465733 2431
rect 465733 2397 465767 2431
rect 465767 2397 465776 2431
rect 465724 2388 465776 2397
rect 470416 2388 470468 2440
rect 474372 2363 474424 2372
rect 474372 2329 474381 2363
rect 474381 2329 474415 2363
rect 474415 2329 474424 2363
rect 474372 2320 474424 2329
rect 478972 2363 479024 2372
rect 478972 2329 478981 2363
rect 478981 2329 479015 2363
rect 479015 2329 479024 2363
rect 478972 2320 479024 2329
rect 413008 2295 413060 2304
rect 413008 2261 413017 2295
rect 413017 2261 413051 2295
rect 413051 2261 413060 2295
rect 413008 2252 413060 2261
rect 416596 2295 416648 2304
rect 416596 2261 416605 2295
rect 416605 2261 416639 2295
rect 416639 2261 416648 2295
rect 416596 2252 416648 2261
rect 426532 2295 426584 2304
rect 426532 2261 426541 2295
rect 426541 2261 426575 2295
rect 426575 2261 426584 2295
rect 426532 2252 426584 2261
rect 440608 2295 440660 2304
rect 440608 2261 440617 2295
rect 440617 2261 440651 2295
rect 440651 2261 440660 2295
rect 440608 2252 440660 2261
rect 448612 2295 448664 2304
rect 448612 2261 448621 2295
rect 448621 2261 448655 2295
rect 448655 2261 448664 2295
rect 448612 2252 448664 2261
rect 452660 2295 452712 2304
rect 452660 2261 452669 2295
rect 452669 2261 452703 2295
rect 452703 2261 452712 2295
rect 452660 2252 452712 2261
rect 453396 2295 453448 2304
rect 453396 2261 453405 2295
rect 453405 2261 453439 2295
rect 453439 2261 453448 2295
rect 453396 2252 453448 2261
rect 461860 2295 461912 2304
rect 461860 2261 461869 2295
rect 461869 2261 461903 2295
rect 461903 2261 461912 2295
rect 461860 2252 461912 2261
rect 466552 2295 466604 2304
rect 466552 2261 466561 2295
rect 466561 2261 466595 2295
rect 466595 2261 466604 2295
rect 466552 2252 466604 2261
rect 470692 2295 470744 2304
rect 470692 2261 470701 2295
rect 470701 2261 470735 2295
rect 470735 2261 470744 2295
rect 470692 2252 470744 2261
rect 475476 2295 475528 2304
rect 475476 2261 475485 2295
rect 475485 2261 475519 2295
rect 475519 2261 475528 2295
rect 475476 2252 475528 2261
rect 479800 2295 479852 2304
rect 479800 2261 479809 2295
rect 479809 2261 479843 2295
rect 479843 2261 479852 2295
rect 479800 2252 479852 2261
rect 492128 2295 492180 2304
rect 492128 2261 492137 2295
rect 492137 2261 492171 2295
rect 492171 2261 492180 2295
rect 492128 2252 492180 2261
rect 500868 2252 500920 2304
rect 67574 2150 67626 2202
rect 67638 2150 67690 2202
rect 67702 2150 67754 2202
rect 67766 2150 67818 2202
rect 67830 2150 67882 2202
rect 199502 2150 199554 2202
rect 199566 2150 199618 2202
rect 199630 2150 199682 2202
rect 199694 2150 199746 2202
rect 199758 2150 199810 2202
rect 331430 2150 331482 2202
rect 331494 2150 331546 2202
rect 331558 2150 331610 2202
rect 331622 2150 331674 2202
rect 331686 2150 331738 2202
rect 463358 2150 463410 2202
rect 463422 2150 463474 2202
rect 463486 2150 463538 2202
rect 463550 2150 463602 2202
rect 463614 2150 463666 2202
rect 26240 2048 26292 2100
rect 31668 2048 31720 2100
rect 37924 2048 37976 2100
rect 103888 2048 103940 2100
rect 108948 2048 109000 2100
rect 202696 2048 202748 2100
rect 226156 2048 226208 2100
rect 306196 2048 306248 2100
rect 307852 2048 307904 2100
rect 316592 2048 316644 2100
rect 22652 1980 22704 2032
rect 62580 1980 62632 2032
rect 70768 1980 70820 2032
rect 120080 1980 120132 2032
rect 128820 1980 128872 2032
rect 223028 1980 223080 2032
rect 231952 1980 232004 2032
rect 306288 1980 306340 2032
rect 306472 1980 306524 2032
rect 349620 2048 349672 2100
rect 386512 2048 386564 2100
rect 478972 2048 479024 2100
rect 25964 1912 26016 1964
rect 41972 1912 42024 1964
rect 42892 1912 42944 1964
rect 136088 1912 136140 1964
rect 154028 1912 154080 1964
rect 248052 1912 248104 1964
rect 337200 1980 337252 2032
rect 350540 1980 350592 2032
rect 425152 1980 425204 2032
rect 426532 1980 426584 2032
rect 494060 1980 494112 2032
rect 21824 1844 21876 1896
rect 66260 1844 66312 1896
rect 75276 1844 75328 1896
rect 168012 1844 168064 1896
rect 200396 1844 200448 1896
rect 211528 1844 211580 1896
rect 244188 1844 244240 1896
rect 307760 1844 307812 1896
rect 24032 1776 24084 1828
rect 31208 1776 31260 1828
rect 27528 1708 27580 1760
rect 31668 1776 31720 1828
rect 48320 1776 48372 1828
rect 74632 1776 74684 1828
rect 111800 1776 111852 1828
rect 212172 1776 212224 1828
rect 307116 1776 307168 1828
rect 311348 1776 311400 1828
rect 313188 1844 313240 1896
rect 335268 1912 335320 1964
rect 349804 1912 349856 1964
rect 371148 1912 371200 1964
rect 390468 1912 390520 1964
rect 397828 1912 397880 1964
rect 440608 1912 440660 1964
rect 488540 1912 488592 1964
rect 346308 1844 346360 1896
rect 350632 1844 350684 1896
rect 389180 1844 389232 1896
rect 399300 1844 399352 1896
rect 399484 1844 399536 1896
rect 408040 1844 408092 1896
rect 448612 1844 448664 1896
rect 485872 1844 485924 1896
rect 346676 1776 346728 1828
rect 408316 1776 408368 1828
rect 453396 1776 453448 1828
rect 484768 1776 484820 1828
rect 126060 1708 126112 1760
rect 127348 1708 127400 1760
rect 216588 1708 216640 1760
rect 307024 1708 307076 1760
rect 2596 1640 2648 1692
rect 31392 1640 31444 1692
rect 31668 1640 31720 1692
rect 96896 1640 96948 1692
rect 112904 1640 112956 1692
rect 206836 1640 206888 1692
rect 208400 1640 208452 1692
rect 246304 1640 246356 1692
rect 305552 1640 305604 1692
rect 319996 1708 320048 1760
rect 329288 1708 329340 1760
rect 338028 1708 338080 1760
rect 389272 1708 389324 1760
rect 399852 1708 399904 1760
rect 408408 1708 408460 1760
rect 475476 1708 475528 1760
rect 502340 1708 502392 1760
rect 21640 1572 21692 1624
rect 24860 1572 24912 1624
rect 28264 1504 28316 1556
rect 31484 1572 31536 1624
rect 115664 1572 115716 1624
rect 208860 1572 208912 1624
rect 213184 1572 213236 1624
rect 307392 1572 307444 1624
rect 345664 1640 345716 1692
rect 354496 1640 354548 1692
rect 447784 1640 447836 1692
rect 466552 1640 466604 1692
rect 489828 1640 489880 1692
rect 352288 1572 352340 1624
rect 380900 1572 380952 1624
rect 474372 1572 474424 1624
rect 479800 1572 479852 1624
rect 496636 1572 496688 1624
rect 28080 1436 28132 1488
rect 33692 1504 33744 1556
rect 58992 1504 59044 1556
rect 152740 1504 152792 1556
rect 206100 1504 206152 1556
rect 300308 1504 300360 1556
rect 306104 1504 306156 1556
rect 354404 1504 354456 1556
rect 399576 1504 399628 1556
rect 105084 1436 105136 1488
rect 116124 1436 116176 1488
rect 120540 1436 120592 1488
rect 212816 1436 212868 1488
rect 213920 1436 213972 1488
rect 309232 1436 309284 1488
rect 332600 1436 332652 1488
rect 401140 1436 401192 1488
rect 401508 1504 401560 1556
rect 407580 1504 407632 1556
rect 407672 1504 407724 1556
rect 405096 1436 405148 1488
rect 406936 1436 406988 1488
rect 410524 1436 410576 1488
rect 28632 1368 28684 1420
rect 23204 1300 23256 1352
rect 26056 1300 26108 1352
rect 26148 1300 26200 1352
rect 31024 1300 31076 1352
rect 216680 1368 216732 1420
rect 311532 1368 311584 1420
rect 400956 1368 401008 1420
rect 402704 1368 402756 1420
rect 405188 1368 405240 1420
rect 407212 1368 407264 1420
rect 461860 1504 461912 1556
rect 495624 1504 495676 1556
rect 478420 1368 478472 1420
rect 32588 1300 32640 1352
rect 33784 1300 33836 1352
rect 117320 1300 117372 1352
rect 117872 1300 117924 1352
rect 210240 1300 210292 1352
rect 306288 1300 306340 1352
rect 325148 1300 325200 1352
rect 346216 1300 346268 1352
rect 355968 1300 356020 1352
rect 358176 1300 358228 1352
rect 407488 1300 407540 1352
rect 408408 1300 408460 1352
rect 21916 1232 21968 1284
rect 29000 1232 29052 1284
rect 30012 1232 30064 1284
rect 31208 1232 31260 1284
rect 31576 1232 31628 1284
rect 117504 1232 117556 1284
rect 121828 1232 121880 1284
rect 215208 1232 215260 1284
rect 306012 1232 306064 1284
rect 389180 1232 389232 1284
rect 394700 1232 394752 1284
rect 398012 1232 398064 1284
rect 398104 1232 398156 1284
rect 20628 1096 20680 1148
rect 20996 756 21048 808
rect 21732 892 21784 944
rect 22100 892 22152 944
rect 23756 1164 23808 1216
rect 28264 1164 28316 1216
rect 24860 1096 24912 1148
rect 28540 1096 28592 1148
rect 27620 1028 27672 1080
rect 23388 960 23440 1012
rect 21824 756 21876 808
rect 21824 484 21876 536
rect 22652 756 22704 808
rect 22928 688 22980 740
rect 23204 688 23256 740
rect 23756 756 23808 808
rect 24032 688 24084 740
rect 24308 756 24360 808
rect 24584 756 24636 808
rect 24860 756 24912 808
rect 26240 892 26292 944
rect 25412 756 25464 808
rect 26424 824 26476 876
rect 27620 892 27672 944
rect 31116 1164 31168 1216
rect 36636 1164 36688 1216
rect 108396 1164 108448 1216
rect 120080 1164 120132 1216
rect 160468 1164 160520 1216
rect 161848 1164 161900 1216
rect 255780 1164 255832 1216
rect 306196 1164 306248 1216
rect 319444 1164 319496 1216
rect 323768 1164 323820 1216
rect 398840 1164 398892 1216
rect 399024 1232 399076 1284
rect 435732 1300 435784 1352
rect 480996 1436 481048 1488
rect 478788 1368 478840 1420
rect 492128 1368 492180 1420
rect 479616 1300 479668 1352
rect 484676 1300 484728 1352
rect 484768 1300 484820 1352
rect 401048 1164 401100 1216
rect 401140 1164 401192 1216
rect 480352 1232 480404 1284
rect 480904 1232 480956 1284
rect 485780 1232 485832 1284
rect 485872 1232 485924 1284
rect 488816 1232 488868 1284
rect 494704 1300 494756 1352
rect 25964 756 26016 808
rect 26148 756 26200 808
rect 26700 756 26752 808
rect 26976 756 27028 808
rect 27528 756 27580 808
rect 28632 824 28684 876
rect 28080 756 28132 808
rect 28356 756 28408 808
rect 29092 892 29144 944
rect 31208 1096 31260 1148
rect 31484 1096 31536 1148
rect 118148 1096 118200 1148
rect 182916 1096 182968 1148
rect 277124 1096 277176 1148
rect 318984 1096 319036 1148
rect 399668 1096 399720 1148
rect 402704 1096 402756 1148
rect 406752 1096 406804 1148
rect 30012 1028 30064 1080
rect 36820 1028 36872 1080
rect 119988 1028 120040 1080
rect 211068 1028 211120 1080
rect 237012 1028 237064 1080
rect 331220 1028 331272 1080
rect 341524 1028 341576 1080
rect 390560 1028 390612 1080
rect 397920 1028 397972 1080
rect 399576 1028 399628 1080
rect 399760 1028 399812 1080
rect 400956 1028 401008 1080
rect 31760 960 31812 1012
rect 112352 960 112404 1012
rect 116124 960 116176 1012
rect 197912 960 197964 1012
rect 199384 960 199436 1012
rect 292580 960 292632 1012
rect 299572 960 299624 1012
rect 393872 960 393924 1012
rect 28632 416 28684 468
rect 29184 756 29236 808
rect 29736 756 29788 808
rect 31300 824 31352 876
rect 36452 892 36504 944
rect 36544 892 36596 944
rect 122840 892 122892 944
rect 210792 892 210844 944
rect 305184 892 305236 944
rect 307760 892 307812 944
rect 337844 892 337896 944
rect 391664 892 391716 944
rect 401140 960 401192 1012
rect 398012 892 398064 944
rect 406936 1028 406988 1080
rect 401324 892 401376 944
rect 31668 824 31720 876
rect 31760 824 31812 876
rect 31852 824 31904 876
rect 121644 824 121696 876
rect 157892 824 157944 876
rect 251732 824 251784 876
rect 254308 824 254360 876
rect 306748 824 306800 876
rect 313372 824 313424 876
rect 36820 756 36872 808
rect 123852 756 123904 808
rect 165528 756 165580 808
rect 258356 756 258408 808
rect 265716 756 265768 808
rect 357900 756 357952 808
rect 111800 688 111852 740
rect 169024 688 169076 740
rect 257068 688 257120 740
rect 346308 688 346360 740
rect 398196 824 398248 876
rect 406384 892 406436 944
rect 401600 824 401652 876
rect 407488 1096 407540 1148
rect 408868 1096 408920 1148
rect 407212 960 407264 1012
rect 411444 1028 411496 1080
rect 413008 1164 413060 1216
rect 486884 1164 486936 1216
rect 488540 1164 488592 1216
rect 500132 1164 500184 1216
rect 416596 1096 416648 1148
rect 480904 1028 480956 1080
rect 480996 1028 481048 1080
rect 482560 1028 482612 1080
rect 482652 1028 482704 1080
rect 494704 1028 494756 1080
rect 407580 960 407632 1012
rect 494520 960 494572 1012
rect 479616 892 479668 944
rect 479708 892 479760 944
rect 397828 756 397880 808
rect 399300 688 399352 740
rect 32864 620 32916 672
rect 117596 620 117648 672
rect 120356 620 120408 672
rect 211436 620 211488 672
rect 212448 620 212500 672
rect 305460 620 305512 672
rect 307300 620 307352 672
rect 332600 620 332652 672
rect 332784 620 332836 672
rect 350540 620 350592 672
rect 395988 620 396040 672
rect 399944 620 399996 672
rect 36452 552 36504 604
rect 125048 552 125100 604
rect 146116 552 146168 604
rect 204904 552 204956 604
rect 206192 552 206244 604
rect 299020 552 299072 604
rect 324688 552 324740 604
rect 397920 552 397972 604
rect 36636 484 36688 536
rect 193588 484 193640 536
rect 285956 484 286008 536
rect 295800 484 295852 536
rect 338028 484 338080 536
rect 33692 416 33744 468
rect 121460 416 121512 468
rect 152188 416 152240 468
rect 208400 416 208452 468
rect 258264 416 258316 468
rect 346584 416 346636 468
rect 356060 416 356112 468
rect 398012 416 398064 468
rect 170772 348 170824 400
rect 264336 348 264388 400
rect 278320 348 278372 400
rect 349804 348 349856 400
rect 352380 348 352432 400
rect 398196 348 398248 400
rect 32588 280 32640 332
rect 121552 280 121604 332
rect 121736 280 121788 332
rect 212632 280 212684 332
rect 247132 280 247184 332
rect 339960 280 340012 332
rect 349712 280 349764 332
rect 398104 280 398156 332
rect 31392 212 31444 264
rect 118700 212 118752 264
rect 218428 212 218480 264
rect 313280 212 313332 264
rect 348424 212 348476 264
rect 399852 212 399904 264
rect 31576 144 31628 196
rect 120172 144 120224 196
rect 215852 144 215904 196
rect 310428 144 310480 196
rect 346768 144 346820 196
rect 399484 144 399536 196
rect 125232 76 125284 128
rect 337292 76 337344 128
rect 399760 76 399812 128
rect 31760 8 31812 60
rect 123760 8 123812 60
rect 315764 8 315816 60
rect 399944 8 399996 60
rect 400220 620 400272 672
rect 400496 416 400548 468
rect 400772 756 400824 808
rect 400956 756 401008 808
rect 401324 756 401376 808
rect 401784 756 401836 808
rect 402060 756 402112 808
rect 402336 756 402388 808
rect 402612 756 402664 808
rect 403164 756 403216 808
rect 403440 620 403492 672
rect 403440 484 403492 536
rect 403716 756 403768 808
rect 403992 756 404044 808
rect 404268 756 404320 808
rect 404544 756 404596 808
rect 404820 756 404872 808
rect 405096 756 405148 808
rect 405372 756 405424 808
rect 405924 756 405976 808
rect 406200 756 406252 808
rect 406200 484 406252 536
rect 406476 756 406528 808
rect 406752 756 406804 808
rect 407212 756 407264 808
rect 407304 756 407356 808
rect 407764 756 407816 808
rect 407764 620 407816 672
rect 408040 756 408092 808
rect 408316 756 408368 808
rect 408592 756 408644 808
rect 408868 756 408920 808
rect 409696 824 409748 876
rect 409420 756 409472 808
rect 409696 484 409748 536
rect 409972 756 410024 808
rect 410248 756 410300 808
rect 410524 756 410576 808
rect 410800 756 410852 808
rect 411076 756 411128 808
rect 411444 824 411496 876
rect 478880 756 478932 808
rect 479708 552 479760 604
rect 470692 8 470744 60
rect 479708 8 479760 60
rect 480352 756 480404 808
rect 481640 756 481692 808
rect 482560 756 482612 808
rect 484584 756 484636 808
rect 484676 756 484728 808
rect 485780 756 485832 808
rect 486884 756 486936 808
rect 488632 756 488684 808
rect 488816 756 488868 808
rect 489920 756 489972 808
rect 491300 756 491352 808
rect 492680 756 492732 808
rect 494060 756 494112 808
rect 494520 688 494572 740
rect 495624 756 495676 808
rect 496636 756 496688 808
rect 499764 756 499816 808
rect 500132 756 500184 808
rect 500868 824 500920 876
rect 502340 756 502392 808
rect 505376 756 505428 808
<< metal2 >>
rect -1076 9784 -756 9796
rect -1076 9728 -1064 9784
rect -1008 9728 -984 9784
rect -928 9728 -904 9784
rect -848 9728 -824 9784
rect -768 9728 -756 9784
rect -1076 9704 -756 9728
rect -1076 9648 -1064 9704
rect -1008 9648 -984 9704
rect -928 9648 -904 9704
rect -848 9648 -824 9704
rect -768 9648 -756 9704
rect -1076 9624 -756 9648
rect -1076 9568 -1064 9624
rect -1008 9568 -984 9624
rect -928 9568 -904 9624
rect -848 9568 -824 9624
rect -768 9568 -756 9624
rect -1076 9544 -756 9568
rect -1076 9488 -1064 9544
rect -1008 9488 -984 9544
rect -928 9488 -904 9544
rect -848 9488 -824 9544
rect -768 9488 -756 9544
rect -1076 7740 -756 9488
rect 1860 9240 1912 9246
rect 1860 9182 1912 9188
rect 34428 9240 34480 9246
rect 34428 9182 34480 9188
rect 52368 9240 52420 9246
rect 52368 9182 52420 9188
rect -1076 7684 -1064 7740
rect -1008 7684 -984 7740
rect -928 7684 -904 7740
rect -848 7684 -824 7740
rect -768 7684 -756 7740
rect -1076 7660 -756 7684
rect -1076 7604 -1064 7660
rect -1008 7604 -984 7660
rect -928 7604 -904 7660
rect -848 7604 -824 7660
rect -768 7604 -756 7660
rect -1076 7580 -756 7604
rect -1076 7524 -1064 7580
rect -1008 7524 -984 7580
rect -928 7524 -904 7580
rect -848 7524 -824 7580
rect -768 7524 -756 7580
rect -1076 7500 -756 7524
rect -1076 7444 -1064 7500
rect -1008 7444 -984 7500
rect -928 7444 -904 7500
rect -848 7444 -824 7500
rect -768 7444 -756 7500
rect -1076 6381 -756 7444
rect -1076 6325 -1064 6381
rect -1008 6325 -984 6381
rect -928 6325 -904 6381
rect -848 6325 -824 6381
rect -768 6325 -756 6381
rect -1076 6301 -756 6325
rect -1076 6245 -1064 6301
rect -1008 6245 -984 6301
rect -928 6245 -904 6301
rect -848 6245 -824 6301
rect -768 6245 -756 6301
rect -1076 6221 -756 6245
rect -1076 6165 -1064 6221
rect -1008 6165 -984 6221
rect -928 6165 -904 6221
rect -848 6165 -824 6221
rect -768 6165 -756 6221
rect -1076 6141 -756 6165
rect -1076 6085 -1064 6141
rect -1008 6085 -984 6141
rect -928 6085 -904 6141
rect -848 6085 -824 6141
rect -768 6085 -756 6141
rect -1076 5022 -756 6085
rect -1076 4966 -1064 5022
rect -1008 4966 -984 5022
rect -928 4966 -904 5022
rect -848 4966 -824 5022
rect -768 4966 -756 5022
rect -1076 4942 -756 4966
rect -1076 4886 -1064 4942
rect -1008 4886 -984 4942
rect -928 4886 -904 4942
rect -848 4886 -824 4942
rect -768 4886 -756 4942
rect -1076 4862 -756 4886
rect -1076 4806 -1064 4862
rect -1008 4806 -984 4862
rect -928 4806 -904 4862
rect -848 4806 -824 4862
rect -768 4806 -756 4862
rect -1076 4782 -756 4806
rect -1076 4726 -1064 4782
rect -1008 4726 -984 4782
rect -928 4726 -904 4782
rect -848 4726 -824 4782
rect -768 4726 -756 4782
rect -1076 3663 -756 4726
rect -1076 3607 -1064 3663
rect -1008 3607 -984 3663
rect -928 3607 -904 3663
rect -848 3607 -824 3663
rect -768 3607 -756 3663
rect -1076 3583 -756 3607
rect -1076 3527 -1064 3583
rect -1008 3527 -984 3583
rect -928 3527 -904 3583
rect -848 3527 -824 3583
rect -768 3527 -756 3583
rect -1076 3503 -756 3527
rect -1076 3447 -1064 3503
rect -1008 3447 -984 3503
rect -928 3447 -904 3503
rect -848 3447 -824 3503
rect -768 3447 -756 3503
rect -1076 3423 -756 3447
rect -1076 3367 -1064 3423
rect -1008 3367 -984 3423
rect -928 3367 -904 3423
rect -848 3367 -824 3423
rect -768 3367 -756 3423
rect -1076 304 -756 3367
rect -416 9124 -96 9136
rect -416 9068 -404 9124
rect -348 9068 -324 9124
rect -268 9068 -244 9124
rect -188 9068 -164 9124
rect -108 9068 -96 9124
rect -416 9044 -96 9068
rect -416 8988 -404 9044
rect -348 8988 -324 9044
rect -268 8988 -244 9044
rect -188 8988 -164 9044
rect -108 8988 -96 9044
rect -416 8964 -96 8988
rect -416 8908 -404 8964
rect -348 8908 -324 8964
rect -268 8908 -244 8964
rect -188 8908 -164 8964
rect -108 8908 -96 8964
rect -416 8884 -96 8908
rect -416 8828 -404 8884
rect -348 8828 -324 8884
rect -268 8828 -244 8884
rect -188 8828 -164 8884
rect -108 8828 -96 8884
rect -416 7080 -96 8828
rect -416 7024 -404 7080
rect -348 7024 -324 7080
rect -268 7024 -244 7080
rect -188 7024 -164 7080
rect -108 7024 -96 7080
rect -416 7000 -96 7024
rect -416 6944 -404 7000
rect -348 6944 -324 7000
rect -268 6944 -244 7000
rect -188 6944 -164 7000
rect -108 6944 -96 7000
rect -416 6920 -96 6944
rect -416 6864 -404 6920
rect -348 6864 -324 6920
rect -268 6864 -244 6920
rect -188 6864 -164 6920
rect -108 6864 -96 6920
rect -416 6840 -96 6864
rect -416 6784 -404 6840
rect -348 6784 -324 6840
rect -268 6784 -244 6840
rect -188 6784 -164 6840
rect -108 6784 -96 6840
rect -416 5721 -96 6784
rect -416 5665 -404 5721
rect -348 5665 -324 5721
rect -268 5665 -244 5721
rect -188 5665 -164 5721
rect -108 5665 -96 5721
rect -416 5641 -96 5665
rect -416 5585 -404 5641
rect -348 5585 -324 5641
rect -268 5585 -244 5641
rect -188 5585 -164 5641
rect -108 5585 -96 5641
rect -416 5561 -96 5585
rect -416 5505 -404 5561
rect -348 5505 -324 5561
rect -268 5505 -244 5561
rect -188 5505 -164 5561
rect -108 5505 -96 5561
rect -416 5481 -96 5505
rect -416 5425 -404 5481
rect -348 5425 -324 5481
rect -268 5425 -244 5481
rect -188 5425 -164 5481
rect -108 5425 -96 5481
rect -416 4362 -96 5425
rect -416 4306 -404 4362
rect -348 4306 -324 4362
rect -268 4306 -244 4362
rect -188 4306 -164 4362
rect -108 4306 -96 4362
rect -416 4282 -96 4306
rect -416 4226 -404 4282
rect -348 4226 -324 4282
rect -268 4226 -244 4282
rect -188 4226 -164 4282
rect -108 4226 -96 4282
rect -416 4202 -96 4226
rect -416 4146 -404 4202
rect -348 4146 -324 4202
rect -268 4146 -244 4202
rect -188 4146 -164 4202
rect -108 4146 -96 4202
rect -416 4122 -96 4146
rect -416 4066 -404 4122
rect -348 4066 -324 4122
rect -268 4066 -244 4122
rect -188 4066 -164 4122
rect -108 4066 -96 4122
rect -416 3003 -96 4066
rect -416 2947 -404 3003
rect -348 2947 -324 3003
rect -268 2947 -244 3003
rect -188 2947 -164 3003
rect -108 2947 -96 3003
rect -416 2923 -96 2947
rect -416 2867 -404 2923
rect -348 2867 -324 2923
rect -268 2867 -244 2923
rect -188 2867 -164 2923
rect -108 2867 -96 2923
rect -416 2843 -96 2867
rect -416 2787 -404 2843
rect -348 2787 -324 2843
rect -268 2787 -244 2843
rect -188 2787 -164 2843
rect -108 2787 -96 2843
rect -416 2763 -96 2787
rect -416 2707 -404 2763
rect -348 2707 -324 2763
rect -268 2707 -244 2763
rect -188 2707 -164 2763
rect -108 2707 -96 2763
rect -416 964 -96 2707
rect 1872 2650 1900 9182
rect 17868 8900 17920 8906
rect 17868 8842 17920 8848
rect 17880 6866 17908 8842
rect 31300 7200 31352 7206
rect 31300 7142 31352 7148
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 19892 6860 19944 6866
rect 19892 6802 19944 6808
rect 19904 2650 19932 6802
rect 27712 6112 27764 6118
rect 27712 6054 27764 6060
rect 26424 5772 26476 5778
rect 26424 5714 26476 5720
rect 24584 5636 24636 5642
rect 24584 5578 24636 5584
rect 23388 4548 23440 4554
rect 23388 4490 23440 4496
rect 22928 4276 22980 4282
rect 22928 4218 22980 4224
rect 20996 4208 21048 4214
rect 20996 4150 21048 4156
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 1860 2644 1912 2650
rect 1860 2586 1912 2592
rect 19892 2644 19944 2650
rect 19892 2586 19944 2592
rect 2596 2304 2648 2310
rect 2596 2246 2648 2252
rect 2608 1698 2636 2246
rect 2596 1692 2648 1698
rect 2596 1634 2648 1640
rect 20732 1442 20760 4014
rect 20640 1414 20760 1442
rect 20640 1154 20668 1414
rect 20628 1148 20680 1154
rect 20628 1090 20680 1096
rect -416 908 -404 964
rect -348 908 -324 964
rect -268 908 -244 964
rect -188 908 -164 964
rect -108 908 -96 964
rect -416 884 -96 908
rect -416 828 -404 884
rect -348 828 -324 884
rect -268 828 -244 884
rect -188 828 -164 884
rect -108 828 -96 884
rect -416 804 -96 828
rect 21008 814 21036 4150
rect 22192 3460 22244 3466
rect 22192 3402 22244 3408
rect 22100 3120 22152 3126
rect 22100 3062 22152 3068
rect 21916 2508 21968 2514
rect 21916 2450 21968 2456
rect 21824 1896 21876 1902
rect 21824 1838 21876 1844
rect 21640 1624 21692 1630
rect 21640 1566 21692 1572
rect -416 748 -404 804
rect -348 748 -324 804
rect -268 748 -244 804
rect -188 748 -164 804
rect -108 748 -96 804
rect 20996 808 21048 814
rect 20996 750 21048 756
rect -416 724 -96 748
rect -416 668 -404 724
rect -348 668 -324 724
rect -268 668 -244 724
rect -188 668 -164 724
rect -108 668 -96 724
rect -416 656 -96 668
rect 21652 490 21680 1566
rect 21732 944 21784 950
rect 21732 886 21784 892
rect 21744 626 21772 886
rect 21836 814 21864 1838
rect 21928 1290 21956 2450
rect 21916 1284 21968 1290
rect 21916 1226 21968 1232
rect 22112 950 22140 3062
rect 22100 944 22152 950
rect 22100 886 22152 892
rect 21824 808 21876 814
rect 21824 750 21876 756
rect 22204 626 22232 3402
rect 22652 2032 22704 2038
rect 22652 1974 22704 1980
rect 22664 814 22692 1974
rect 22652 808 22704 814
rect 22652 750 22704 756
rect 22940 746 22968 4218
rect 23204 1352 23256 1358
rect 23204 1294 23256 1300
rect 23216 746 23244 1294
rect 23400 1018 23428 4490
rect 24308 2372 24360 2378
rect 24308 2314 24360 2320
rect 24032 1828 24084 1834
rect 24032 1770 24084 1776
rect 23756 1216 23808 1222
rect 23756 1158 23808 1164
rect 23388 1012 23440 1018
rect 23388 954 23440 960
rect 23768 814 23796 1158
rect 23756 808 23808 814
rect 23756 750 23808 756
rect 24044 746 24072 1770
rect 24320 814 24348 2314
rect 24596 814 24624 5578
rect 25412 5568 25464 5574
rect 25412 5510 25464 5516
rect 24860 2984 24912 2990
rect 24860 2926 24912 2932
rect 24872 1630 24900 2926
rect 24860 1624 24912 1630
rect 24860 1566 24912 1572
rect 24860 1148 24912 1154
rect 24860 1090 24912 1096
rect 24872 814 24900 1090
rect 25424 814 25452 5510
rect 26240 2100 26292 2106
rect 26240 2042 26292 2048
rect 25964 1964 26016 1970
rect 25964 1906 26016 1912
rect 25976 814 26004 1906
rect 26054 1592 26110 1601
rect 26054 1527 26110 1536
rect 26068 1358 26096 1527
rect 26056 1352 26108 1358
rect 26056 1294 26108 1300
rect 26148 1352 26200 1358
rect 26148 1294 26200 1300
rect 26160 814 26188 1294
rect 26252 950 26280 2042
rect 26240 944 26292 950
rect 26240 886 26292 892
rect 26436 882 26464 5714
rect 27620 3188 27672 3194
rect 27620 3130 27672 3136
rect 26700 2304 26752 2310
rect 26700 2246 26752 2252
rect 26424 876 26476 882
rect 26424 818 26476 824
rect 26712 814 26740 2246
rect 27528 1760 27580 1766
rect 27528 1702 27580 1708
rect 26974 1456 27030 1465
rect 26974 1391 27030 1400
rect 26988 814 27016 1391
rect 27540 814 27568 1702
rect 27632 1086 27660 3130
rect 27620 1080 27672 1086
rect 27620 1022 27672 1028
rect 27620 944 27672 950
rect 27724 932 27752 6054
rect 29736 5908 29788 5914
rect 29736 5850 29788 5856
rect 28356 4616 28408 4622
rect 28356 4558 28408 4564
rect 28264 1556 28316 1562
rect 28264 1498 28316 1504
rect 28080 1488 28132 1494
rect 28080 1430 28132 1436
rect 27672 904 27752 932
rect 27620 886 27672 892
rect 28092 814 28120 1430
rect 28276 1222 28304 1498
rect 28264 1216 28316 1222
rect 28264 1158 28316 1164
rect 28368 814 28396 4558
rect 29000 2848 29052 2854
rect 29000 2790 29052 2796
rect 28632 1420 28684 1426
rect 28632 1362 28684 1368
rect 28538 1184 28594 1193
rect 28538 1119 28540 1128
rect 28592 1119 28594 1128
rect 28540 1090 28592 1096
rect 28644 882 28672 1362
rect 29012 1290 29040 2790
rect 29184 2644 29236 2650
rect 29184 2586 29236 2592
rect 29090 1864 29146 1873
rect 29090 1799 29146 1808
rect 29000 1284 29052 1290
rect 29000 1226 29052 1232
rect 29104 950 29132 1799
rect 29092 944 29144 950
rect 29092 886 29144 892
rect 28632 876 28684 882
rect 28632 818 28684 824
rect 29196 814 29224 2586
rect 29748 814 29776 5850
rect 31208 1828 31260 1834
rect 31208 1770 31260 1776
rect 31220 1737 31248 1770
rect 31206 1728 31262 1737
rect 31206 1663 31262 1672
rect 31024 1352 31076 1358
rect 31024 1294 31076 1300
rect 31206 1320 31262 1329
rect 30012 1284 30064 1290
rect 30012 1226 30064 1232
rect 30024 1086 30052 1226
rect 30012 1080 30064 1086
rect 30012 1022 30064 1028
rect 24308 808 24360 814
rect 24308 750 24360 756
rect 24584 808 24636 814
rect 24584 750 24636 756
rect 24860 808 24912 814
rect 24860 750 24912 756
rect 25412 808 25464 814
rect 25412 750 25464 756
rect 25964 808 26016 814
rect 25964 750 26016 756
rect 26148 808 26200 814
rect 26148 750 26200 756
rect 26700 808 26752 814
rect 26700 750 26752 756
rect 26976 808 27028 814
rect 26976 750 27028 756
rect 27528 808 27580 814
rect 27528 750 27580 756
rect 28080 808 28132 814
rect 28080 750 28132 756
rect 28356 808 28408 814
rect 28356 750 28408 756
rect 29184 808 29236 814
rect 29184 750 29236 756
rect 29736 808 29788 814
rect 29736 750 29788 756
rect 22928 740 22980 746
rect 22928 682 22980 688
rect 23204 740 23256 746
rect 23204 682 23256 688
rect 24032 740 24084 746
rect 24032 682 24084 688
rect 21744 598 22232 626
rect 21824 536 21876 542
rect 21652 484 21824 490
rect 21652 478 21876 484
rect 28630 504 28686 513
rect 21652 462 21864 478
rect 28630 439 28632 448
rect 28684 439 28686 448
rect 28632 410 28684 416
rect -1076 248 -1064 304
rect -1008 248 -984 304
rect -928 248 -904 304
rect -848 248 -824 304
rect -768 248 -756 304
rect -1076 224 -756 248
rect -1076 168 -1064 224
rect -1008 168 -984 224
rect -928 168 -904 224
rect -848 168 -824 224
rect -768 168 -756 224
rect 31036 218 31064 1294
rect 31206 1255 31208 1264
rect 31260 1255 31262 1264
rect 31208 1226 31260 1232
rect 31116 1216 31168 1222
rect 31116 1158 31168 1164
rect 31128 354 31156 1158
rect 31208 1148 31260 1154
rect 31208 1090 31260 1096
rect 31220 762 31248 1090
rect 31312 882 31340 7142
rect 34440 6866 34468 9182
rect 52380 6866 52408 9182
rect 66908 9124 67228 9796
rect 66908 9068 66920 9124
rect 66976 9068 67000 9124
rect 67056 9068 67080 9124
rect 67136 9068 67160 9124
rect 67216 9068 67228 9124
rect 66908 9044 67228 9068
rect 66908 8988 66920 9044
rect 66976 8988 67000 9044
rect 67056 8988 67080 9044
rect 67136 8988 67160 9044
rect 67216 8988 67228 9044
rect 66908 8964 67228 8988
rect 66908 8908 66920 8964
rect 66976 8908 67000 8964
rect 67056 8908 67080 8964
rect 67136 8908 67160 8964
rect 67216 8908 67228 8964
rect 66908 8884 67228 8908
rect 66908 8828 66920 8884
rect 66976 8828 67000 8884
rect 67056 8828 67080 8884
rect 67136 8828 67160 8884
rect 67216 8828 67228 8884
rect 66908 7098 67228 8828
rect 66908 7046 66914 7098
rect 66966 7080 66978 7098
rect 67030 7080 67042 7098
rect 67094 7080 67106 7098
rect 67158 7080 67170 7098
rect 66976 7046 66978 7080
rect 67158 7046 67160 7080
rect 67222 7046 67228 7098
rect 66908 7024 66920 7046
rect 66976 7024 67000 7046
rect 67056 7024 67080 7046
rect 67136 7024 67160 7046
rect 67216 7024 67228 7046
rect 66908 7000 67228 7024
rect 66908 6944 66920 7000
rect 66976 6944 67000 7000
rect 67056 6944 67080 7000
rect 67136 6944 67160 7000
rect 67216 6944 67228 7000
rect 66908 6920 67228 6944
rect 34428 6860 34480 6866
rect 34428 6802 34480 6808
rect 37648 6860 37700 6866
rect 37648 6802 37700 6808
rect 52368 6860 52420 6866
rect 52368 6802 52420 6808
rect 53840 6860 53892 6866
rect 53840 6802 53892 6808
rect 66908 6864 66920 6920
rect 66976 6864 67000 6920
rect 67056 6864 67080 6920
rect 67136 6864 67160 6920
rect 67216 6864 67228 6920
rect 66908 6840 67228 6864
rect 37372 2984 37424 2990
rect 37556 2984 37608 2990
rect 37424 2932 37556 2938
rect 37372 2926 37608 2932
rect 31760 2916 31812 2922
rect 37384 2910 37596 2926
rect 31760 2858 31812 2864
rect 31772 2446 31800 2858
rect 37660 2854 37688 6802
rect 37648 2848 37700 2854
rect 37648 2790 37700 2796
rect 37660 2446 37688 2790
rect 53852 2650 53880 6802
rect 66908 6784 66920 6840
rect 66976 6784 67000 6840
rect 67056 6784 67080 6840
rect 67136 6784 67160 6840
rect 67216 6784 67228 6840
rect 66908 6010 67228 6784
rect 66908 5958 66914 6010
rect 66966 5958 66978 6010
rect 67030 5958 67042 6010
rect 67094 5958 67106 6010
rect 67158 5958 67170 6010
rect 67222 5958 67228 6010
rect 66908 5721 67228 5958
rect 66908 5665 66920 5721
rect 66976 5665 67000 5721
rect 67056 5665 67080 5721
rect 67136 5665 67160 5721
rect 67216 5665 67228 5721
rect 66908 5641 67228 5665
rect 66908 5585 66920 5641
rect 66976 5585 67000 5641
rect 67056 5585 67080 5641
rect 67136 5585 67160 5641
rect 67216 5585 67228 5641
rect 66908 5561 67228 5585
rect 66908 5505 66920 5561
rect 66976 5505 67000 5561
rect 67056 5505 67080 5561
rect 67136 5505 67160 5561
rect 67216 5505 67228 5561
rect 66908 5481 67228 5505
rect 66908 5425 66920 5481
rect 66976 5425 67000 5481
rect 67056 5425 67080 5481
rect 67136 5425 67160 5481
rect 67216 5425 67228 5481
rect 63592 5160 63644 5166
rect 63592 5102 63644 5108
rect 63500 4820 63552 4826
rect 63500 4762 63552 4768
rect 58164 4548 58216 4554
rect 58164 4490 58216 4496
rect 56508 3936 56560 3942
rect 56508 3878 56560 3884
rect 53840 2644 53892 2650
rect 53840 2586 53892 2592
rect 56520 2582 56548 3878
rect 58176 2650 58204 4490
rect 58164 2644 58216 2650
rect 58164 2586 58216 2592
rect 56508 2576 56560 2582
rect 54666 2544 54722 2553
rect 56508 2518 56560 2524
rect 54666 2479 54722 2488
rect 55864 2508 55916 2514
rect 54680 2446 54708 2479
rect 55864 2450 55916 2456
rect 31760 2440 31812 2446
rect 31760 2382 31812 2388
rect 35900 2440 35952 2446
rect 35900 2382 35952 2388
rect 37648 2440 37700 2446
rect 37648 2382 37700 2388
rect 41972 2440 42024 2446
rect 41972 2382 42024 2388
rect 48320 2440 48372 2446
rect 48320 2382 48372 2388
rect 54668 2440 54720 2446
rect 54668 2382 54720 2388
rect 35912 2310 35940 2382
rect 36728 2372 36780 2378
rect 36728 2314 36780 2320
rect 35900 2304 35952 2310
rect 35900 2246 35952 2252
rect 31668 2100 31720 2106
rect 31668 2042 31720 2048
rect 31680 1834 31708 2042
rect 36740 2009 36768 2314
rect 41984 2310 42012 2382
rect 42892 2372 42944 2378
rect 42892 2314 42944 2320
rect 37924 2304 37976 2310
rect 37924 2246 37976 2252
rect 41972 2304 42024 2310
rect 41972 2246 42024 2252
rect 37936 2106 37964 2246
rect 37924 2100 37976 2106
rect 37924 2042 37976 2048
rect 36726 2000 36782 2009
rect 41984 1970 42012 2246
rect 42904 1970 42932 2314
rect 48332 2310 48360 2382
rect 55876 2310 55904 2450
rect 58176 2446 58204 2586
rect 63512 2446 63540 4762
rect 63604 2650 63632 5102
rect 66908 4922 67228 5425
rect 66908 4870 66914 4922
rect 66966 4870 66978 4922
rect 67030 4870 67042 4922
rect 67094 4870 67106 4922
rect 67158 4870 67170 4922
rect 67222 4870 67228 4922
rect 66908 4362 67228 4870
rect 66908 4306 66920 4362
rect 66976 4306 67000 4362
rect 67056 4306 67080 4362
rect 67136 4306 67160 4362
rect 67216 4306 67228 4362
rect 66908 4282 67228 4306
rect 66908 4226 66920 4282
rect 66976 4226 67000 4282
rect 67056 4226 67080 4282
rect 67136 4226 67160 4282
rect 67216 4226 67228 4282
rect 66908 4202 67228 4226
rect 66908 4146 66920 4202
rect 66976 4146 67000 4202
rect 67056 4146 67080 4202
rect 67136 4146 67160 4202
rect 67216 4146 67228 4202
rect 66908 4122 67228 4146
rect 66908 4066 66920 4122
rect 66976 4066 67000 4122
rect 67056 4066 67080 4122
rect 67136 4066 67160 4122
rect 67216 4066 67228 4122
rect 66908 3834 67228 4066
rect 66908 3782 66914 3834
rect 66966 3782 66978 3834
rect 67030 3782 67042 3834
rect 67094 3782 67106 3834
rect 67158 3782 67170 3834
rect 67222 3782 67228 3834
rect 66908 3003 67228 3782
rect 66908 2947 66920 3003
rect 66976 2947 67000 3003
rect 67056 2947 67080 3003
rect 67136 2947 67160 3003
rect 67216 2947 67228 3003
rect 66908 2923 67228 2947
rect 66908 2867 66920 2923
rect 66976 2867 67000 2923
rect 67056 2867 67080 2923
rect 67136 2867 67160 2923
rect 67216 2867 67228 2923
rect 66908 2843 67228 2867
rect 66908 2787 66920 2843
rect 66976 2787 67000 2843
rect 67056 2787 67080 2843
rect 67136 2787 67160 2843
rect 67216 2787 67228 2843
rect 66908 2763 67228 2787
rect 66908 2746 66920 2763
rect 66976 2746 67000 2763
rect 67056 2746 67080 2763
rect 67136 2746 67160 2763
rect 67216 2746 67228 2763
rect 66908 2694 66914 2746
rect 66976 2707 66978 2746
rect 67158 2707 67160 2746
rect 66966 2694 66978 2707
rect 67030 2694 67042 2707
rect 67094 2694 67106 2707
rect 67158 2694 67170 2707
rect 67222 2694 67228 2746
rect 63592 2644 63644 2650
rect 63592 2586 63644 2592
rect 58164 2440 58216 2446
rect 58164 2382 58216 2388
rect 63500 2440 63552 2446
rect 63500 2382 63552 2388
rect 58992 2372 59044 2378
rect 58992 2314 59044 2320
rect 48320 2304 48372 2310
rect 48320 2246 48372 2252
rect 55864 2304 55916 2310
rect 55864 2246 55916 2252
rect 36726 1935 36782 1944
rect 41972 1964 42024 1970
rect 41972 1906 42024 1912
rect 42892 1964 42944 1970
rect 42892 1906 42944 1912
rect 36542 1864 36598 1873
rect 31668 1828 31720 1834
rect 48332 1834 48360 2246
rect 36542 1799 36598 1808
rect 48320 1828 48372 1834
rect 31668 1770 31720 1776
rect 33782 1728 33838 1737
rect 31404 1698 31708 1714
rect 31392 1692 31720 1698
rect 31444 1686 31668 1692
rect 31392 1634 31444 1640
rect 33782 1663 33838 1672
rect 31668 1634 31720 1640
rect 31484 1624 31536 1630
rect 31484 1566 31536 1572
rect 32862 1592 32918 1601
rect 31496 1154 31524 1566
rect 32862 1527 32918 1536
rect 33692 1556 33744 1562
rect 31850 1456 31906 1465
rect 31850 1391 31906 1400
rect 31758 1320 31814 1329
rect 31576 1284 31628 1290
rect 31758 1255 31814 1264
rect 31576 1226 31628 1232
rect 31588 1193 31616 1226
rect 31574 1184 31630 1193
rect 31484 1148 31536 1154
rect 31574 1119 31630 1128
rect 31484 1090 31536 1096
rect 31772 1018 31800 1255
rect 31760 1012 31812 1018
rect 31760 954 31812 960
rect 31864 882 31892 1391
rect 32588 1352 32640 1358
rect 32588 1294 32640 1300
rect 31300 876 31352 882
rect 31668 876 31720 882
rect 31300 818 31352 824
rect 31588 836 31668 864
rect 31588 762 31616 836
rect 31668 818 31720 824
rect 31760 876 31812 882
rect 31760 818 31812 824
rect 31852 876 31904 882
rect 31852 818 31904 824
rect 31220 734 31616 762
rect 31128 326 31616 354
rect 31392 264 31444 270
rect 31036 212 31392 218
rect 31036 206 31444 212
rect 31036 190 31432 206
rect 31588 202 31616 326
rect 31576 196 31628 202
rect -1076 144 -756 168
rect -1076 88 -1064 144
rect -1008 88 -984 144
rect -928 88 -904 144
rect -848 88 -824 144
rect -768 88 -756 144
rect 31576 138 31628 144
rect -1076 64 -756 88
rect 31772 66 31800 818
rect 32600 338 32628 1294
rect 32876 678 32904 1527
rect 33692 1498 33744 1504
rect 32864 672 32916 678
rect 32864 614 32916 620
rect 33704 474 33732 1498
rect 33796 1358 33824 1663
rect 33784 1352 33836 1358
rect 33784 1294 33836 1300
rect 36556 950 36584 1799
rect 48320 1770 48372 1776
rect 59004 1562 59032 2314
rect 62580 2304 62632 2310
rect 62580 2246 62632 2252
rect 66260 2304 66312 2310
rect 66260 2246 66312 2252
rect 62592 2038 62620 2246
rect 62580 2032 62632 2038
rect 62580 1974 62632 1980
rect 66272 1902 66300 2246
rect 66260 1896 66312 1902
rect 66260 1838 66312 1844
rect 58992 1556 59044 1562
rect 58992 1498 59044 1504
rect 36636 1216 36688 1222
rect 36636 1158 36688 1164
rect 36452 944 36504 950
rect 36452 886 36504 892
rect 36544 944 36596 950
rect 36544 886 36596 892
rect 36464 610 36492 886
rect 36452 604 36504 610
rect 36452 546 36504 552
rect 36648 542 36676 1158
rect 36820 1080 36872 1086
rect 36820 1022 36872 1028
rect 36832 814 36860 1022
rect 66908 964 67228 2694
rect 66908 908 66920 964
rect 66976 908 67000 964
rect 67056 908 67080 964
rect 67136 908 67160 964
rect 67216 908 67228 964
rect 66908 884 67228 908
rect 66908 828 66920 884
rect 66976 828 67000 884
rect 67056 828 67080 884
rect 67136 828 67160 884
rect 67216 828 67228 884
rect 36820 808 36872 814
rect 36820 750 36872 756
rect 66908 804 67228 828
rect 66908 748 66920 804
rect 66976 748 67000 804
rect 67056 748 67080 804
rect 67136 748 67160 804
rect 67216 748 67228 804
rect 66908 724 67228 748
rect 66908 668 66920 724
rect 66976 668 67000 724
rect 67056 668 67080 724
rect 67136 668 67160 724
rect 67216 668 67228 724
rect 36636 536 36688 542
rect 36636 478 36688 484
rect 33692 468 33744 474
rect 33692 410 33744 416
rect 32588 332 32640 338
rect 32588 274 32640 280
rect -1076 8 -1064 64
rect -1008 8 -984 64
rect -928 8 -904 64
rect -848 8 -824 64
rect -768 8 -756 64
rect -1076 -4 -756 8
rect 31760 60 31812 66
rect 31760 2 31812 8
rect 66908 -4 67228 668
rect 67568 9784 67888 9796
rect 67568 9728 67580 9784
rect 67636 9728 67660 9784
rect 67716 9728 67740 9784
rect 67796 9728 67820 9784
rect 67876 9728 67888 9784
rect 67568 9704 67888 9728
rect 67568 9648 67580 9704
rect 67636 9648 67660 9704
rect 67716 9648 67740 9704
rect 67796 9648 67820 9704
rect 67876 9648 67888 9704
rect 67568 9624 67888 9648
rect 67568 9568 67580 9624
rect 67636 9568 67660 9624
rect 67716 9568 67740 9624
rect 67796 9568 67820 9624
rect 67876 9568 67888 9624
rect 67568 9544 67888 9568
rect 67568 9488 67580 9544
rect 67636 9488 67660 9544
rect 67716 9488 67740 9544
rect 67796 9488 67820 9544
rect 67876 9488 67888 9544
rect 67568 7740 67888 9488
rect 68928 9240 68980 9246
rect 68928 9182 68980 9188
rect 102232 9240 102284 9246
rect 102232 9182 102284 9188
rect 119988 9240 120040 9246
rect 119988 9182 120040 9188
rect 136548 9240 136600 9246
rect 136548 9182 136600 9188
rect 187608 9240 187660 9246
rect 187608 9182 187660 9188
rect 67568 7684 67580 7740
rect 67636 7684 67660 7740
rect 67716 7684 67740 7740
rect 67796 7684 67820 7740
rect 67876 7684 67888 7740
rect 67568 7660 67888 7684
rect 67568 7642 67580 7660
rect 67636 7642 67660 7660
rect 67716 7642 67740 7660
rect 67796 7642 67820 7660
rect 67876 7642 67888 7660
rect 67568 7590 67574 7642
rect 67636 7604 67638 7642
rect 67818 7604 67820 7642
rect 67626 7590 67638 7604
rect 67690 7590 67702 7604
rect 67754 7590 67766 7604
rect 67818 7590 67830 7604
rect 67882 7590 67888 7642
rect 67568 7580 67888 7590
rect 67568 7524 67580 7580
rect 67636 7524 67660 7580
rect 67716 7524 67740 7580
rect 67796 7524 67820 7580
rect 67876 7524 67888 7580
rect 67568 7500 67888 7524
rect 67568 7444 67580 7500
rect 67636 7444 67660 7500
rect 67716 7444 67740 7500
rect 67796 7444 67820 7500
rect 67876 7444 67888 7500
rect 67568 6554 67888 7444
rect 68940 6866 68968 9182
rect 85488 8900 85540 8906
rect 85488 8842 85540 8848
rect 85500 6866 85528 8842
rect 68928 6860 68980 6866
rect 68928 6802 68980 6808
rect 73988 6860 74040 6866
rect 73988 6802 74040 6808
rect 85488 6860 85540 6866
rect 85488 6802 85540 6808
rect 92020 6860 92072 6866
rect 92020 6802 92072 6808
rect 67568 6502 67574 6554
rect 67626 6502 67638 6554
rect 67690 6502 67702 6554
rect 67754 6502 67766 6554
rect 67818 6502 67830 6554
rect 67882 6502 67888 6554
rect 67568 6381 67888 6502
rect 67568 6325 67580 6381
rect 67636 6325 67660 6381
rect 67716 6325 67740 6381
rect 67796 6325 67820 6381
rect 67876 6325 67888 6381
rect 67568 6301 67888 6325
rect 67568 6245 67580 6301
rect 67636 6245 67660 6301
rect 67716 6245 67740 6301
rect 67796 6245 67820 6301
rect 67876 6245 67888 6301
rect 67568 6221 67888 6245
rect 67568 6165 67580 6221
rect 67636 6165 67660 6221
rect 67716 6165 67740 6221
rect 67796 6165 67820 6221
rect 67876 6165 67888 6221
rect 67568 6141 67888 6165
rect 67568 6085 67580 6141
rect 67636 6085 67660 6141
rect 67716 6085 67740 6141
rect 67796 6085 67820 6141
rect 67876 6085 67888 6141
rect 67568 5466 67888 6085
rect 67568 5414 67574 5466
rect 67626 5414 67638 5466
rect 67690 5414 67702 5466
rect 67754 5414 67766 5466
rect 67818 5414 67830 5466
rect 67882 5414 67888 5466
rect 67568 5022 67888 5414
rect 67568 4966 67580 5022
rect 67636 4966 67660 5022
rect 67716 4966 67740 5022
rect 67796 4966 67820 5022
rect 67876 4966 67888 5022
rect 67568 4942 67888 4966
rect 67568 4886 67580 4942
rect 67636 4886 67660 4942
rect 67716 4886 67740 4942
rect 67796 4886 67820 4942
rect 67876 4886 67888 4942
rect 67568 4862 67888 4886
rect 67568 4806 67580 4862
rect 67636 4806 67660 4862
rect 67716 4806 67740 4862
rect 67796 4806 67820 4862
rect 67876 4806 67888 4862
rect 67568 4782 67888 4806
rect 67568 4726 67580 4782
rect 67636 4726 67660 4782
rect 67716 4726 67740 4782
rect 67796 4726 67820 4782
rect 67876 4726 67888 4782
rect 67568 4378 67888 4726
rect 67568 4326 67574 4378
rect 67626 4326 67638 4378
rect 67690 4326 67702 4378
rect 67754 4326 67766 4378
rect 67818 4326 67830 4378
rect 67882 4326 67888 4378
rect 67568 3663 67888 4326
rect 70400 4208 70452 4214
rect 70400 4150 70452 4156
rect 67568 3607 67580 3663
rect 67636 3607 67660 3663
rect 67716 3607 67740 3663
rect 67796 3607 67820 3663
rect 67876 3607 67888 3663
rect 67568 3583 67888 3607
rect 67568 3527 67580 3583
rect 67636 3527 67660 3583
rect 67716 3527 67740 3583
rect 67796 3527 67820 3583
rect 67876 3527 67888 3583
rect 67568 3503 67888 3527
rect 67568 3447 67580 3503
rect 67636 3447 67660 3503
rect 67716 3447 67740 3503
rect 67796 3447 67820 3503
rect 67876 3447 67888 3503
rect 67568 3423 67888 3447
rect 67568 3367 67580 3423
rect 67636 3367 67660 3423
rect 67716 3367 67740 3423
rect 67796 3367 67820 3423
rect 67876 3367 67888 3423
rect 67568 3290 67888 3367
rect 67568 3238 67574 3290
rect 67626 3238 67638 3290
rect 67690 3238 67702 3290
rect 67754 3238 67766 3290
rect 67818 3238 67830 3290
rect 67882 3238 67888 3290
rect 67568 2202 67888 3238
rect 70412 2650 70440 4150
rect 74000 2650 74028 6802
rect 74724 2848 74776 2854
rect 74724 2790 74776 2796
rect 75000 2848 75052 2854
rect 75000 2790 75052 2796
rect 70400 2644 70452 2650
rect 70400 2586 70452 2592
rect 71044 2644 71096 2650
rect 71044 2586 71096 2592
rect 73988 2644 74040 2650
rect 73988 2586 74040 2592
rect 74540 2644 74592 2650
rect 74540 2586 74592 2592
rect 71056 2446 71084 2586
rect 74552 2514 74580 2586
rect 74540 2508 74592 2514
rect 74540 2450 74592 2456
rect 74736 2446 74764 2790
rect 75012 2514 75040 2790
rect 75000 2508 75052 2514
rect 75000 2450 75052 2456
rect 92032 2446 92060 6802
rect 102244 6186 102272 9182
rect 120000 6866 120028 9182
rect 125416 7200 125468 7206
rect 125416 7142 125468 7148
rect 125876 7200 125928 7206
rect 125876 7142 125928 7148
rect 125140 6996 125192 7002
rect 125140 6938 125192 6944
rect 124496 6928 124548 6934
rect 124496 6870 124548 6876
rect 119988 6860 120040 6866
rect 119988 6802 120040 6808
rect 114192 6248 114244 6254
rect 114192 6190 114244 6196
rect 102232 6180 102284 6186
rect 102232 6122 102284 6128
rect 110052 6180 110104 6186
rect 110052 6122 110104 6128
rect 98644 4208 98696 4214
rect 98644 4150 98696 4156
rect 98656 2446 98684 4150
rect 108304 3596 108356 3602
rect 108304 3538 108356 3544
rect 108316 3058 108344 3538
rect 108304 3052 108356 3058
rect 108304 2994 108356 3000
rect 108396 2848 108448 2854
rect 108396 2790 108448 2796
rect 108408 2446 108436 2790
rect 71044 2440 71096 2446
rect 71044 2382 71096 2388
rect 74632 2440 74684 2446
rect 74632 2382 74684 2388
rect 74724 2440 74776 2446
rect 74724 2382 74776 2388
rect 92020 2440 92072 2446
rect 92296 2440 92348 2446
rect 92072 2388 92296 2394
rect 92020 2382 92348 2388
rect 98644 2440 98696 2446
rect 98644 2382 98696 2388
rect 103888 2440 103940 2446
rect 107660 2440 107712 2446
rect 103888 2382 103940 2388
rect 107658 2408 107660 2417
rect 108396 2440 108448 2446
rect 107712 2408 107714 2417
rect 70768 2372 70820 2378
rect 70768 2314 70820 2320
rect 67568 2150 67574 2202
rect 67626 2150 67638 2202
rect 67690 2150 67702 2202
rect 67754 2150 67766 2202
rect 67818 2150 67830 2202
rect 67882 2150 67888 2202
rect 67568 304 67888 2150
rect 70780 2038 70808 2314
rect 70768 2032 70820 2038
rect 70768 1974 70820 1980
rect 74644 1834 74672 2382
rect 75276 2372 75328 2378
rect 92032 2366 92336 2382
rect 96896 2372 96948 2378
rect 75276 2314 75328 2320
rect 96896 2314 96948 2320
rect 75288 1902 75316 2314
rect 75276 1896 75328 1902
rect 75276 1838 75328 1844
rect 74632 1828 74684 1834
rect 74632 1770 74684 1776
rect 96908 1698 96936 2314
rect 103900 2106 103928 2382
rect 105084 2372 105136 2378
rect 108396 2382 108448 2388
rect 107658 2343 107714 2352
rect 105084 2314 105136 2320
rect 103888 2100 103940 2106
rect 103888 2042 103940 2048
rect 96896 1692 96948 1698
rect 96896 1634 96948 1640
rect 105096 1494 105124 2314
rect 105084 1488 105136 1494
rect 105084 1430 105136 1436
rect 108408 1222 108436 2382
rect 108948 2372 109000 2378
rect 108948 2314 109000 2320
rect 108960 2106 108988 2314
rect 110064 2310 110092 6122
rect 110788 5228 110840 5234
rect 110788 5170 110840 5176
rect 110800 2514 110828 5170
rect 114100 3732 114152 3738
rect 114100 3674 114152 3680
rect 114112 3058 114140 3674
rect 113364 3052 113416 3058
rect 113364 2994 113416 3000
rect 114100 3052 114152 3058
rect 114100 2994 114152 3000
rect 112352 2848 112404 2854
rect 112352 2790 112404 2796
rect 110788 2508 110840 2514
rect 110788 2450 110840 2456
rect 112364 2446 112392 2790
rect 113376 2514 113404 2994
rect 114204 2854 114232 6190
rect 120264 6112 120316 6118
rect 120264 6054 120316 6060
rect 117320 5840 117372 5846
rect 117320 5782 117372 5788
rect 116216 5024 116268 5030
rect 116216 4966 116268 4972
rect 116676 5024 116728 5030
rect 116676 4966 116728 4972
rect 115664 4480 115716 4486
rect 115664 4422 115716 4428
rect 116032 4480 116084 4486
rect 116032 4422 116084 4428
rect 114928 3596 114980 3602
rect 114928 3538 114980 3544
rect 114192 2848 114244 2854
rect 114192 2790 114244 2796
rect 113364 2508 113416 2514
rect 113364 2450 113416 2456
rect 114204 2446 114232 2790
rect 114940 2514 114968 3538
rect 115676 3058 115704 4422
rect 116044 4162 116072 4422
rect 115768 4146 116072 4162
rect 115756 4140 116072 4146
rect 115808 4134 116072 4140
rect 115756 4082 115808 4088
rect 116044 3670 116072 4134
rect 116032 3664 116084 3670
rect 116032 3606 116084 3612
rect 116124 3460 116176 3466
rect 116124 3402 116176 3408
rect 116136 3194 116164 3402
rect 116124 3188 116176 3194
rect 116124 3130 116176 3136
rect 115664 3052 115716 3058
rect 115664 2994 115716 3000
rect 114928 2508 114980 2514
rect 114928 2450 114980 2456
rect 112352 2440 112404 2446
rect 112352 2382 112404 2388
rect 114192 2440 114244 2446
rect 114192 2382 114244 2388
rect 110052 2304 110104 2310
rect 110052 2246 110104 2252
rect 108948 2100 109000 2106
rect 108948 2042 109000 2048
rect 111800 1828 111852 1834
rect 111800 1770 111852 1776
rect 108396 1216 108448 1222
rect 108396 1158 108448 1164
rect 111812 746 111840 1770
rect 112364 1018 112392 2382
rect 112904 2372 112956 2378
rect 112904 2314 112956 2320
rect 112916 1698 112944 2314
rect 112904 1692 112956 1698
rect 112904 1634 112956 1640
rect 115676 1630 115704 2994
rect 116228 2446 116256 4966
rect 116584 4480 116636 4486
rect 116584 4422 116636 4428
rect 116308 4276 116360 4282
rect 116308 4218 116360 4224
rect 116320 3126 116348 4218
rect 116596 4146 116624 4422
rect 116584 4140 116636 4146
rect 116584 4082 116636 4088
rect 116688 3942 116716 4966
rect 116676 3936 116728 3942
rect 116676 3878 116728 3884
rect 116688 3534 116716 3878
rect 117332 3602 117360 5782
rect 120080 5772 120132 5778
rect 120080 5714 120132 5720
rect 117412 5704 117464 5710
rect 117412 5646 117464 5652
rect 117424 3738 117452 5646
rect 118792 5636 118844 5642
rect 118792 5578 118844 5584
rect 119344 5636 119396 5642
rect 119344 5578 119396 5584
rect 118700 5568 118752 5574
rect 118700 5510 118752 5516
rect 117504 5024 117556 5030
rect 117504 4966 117556 4972
rect 118056 5024 118108 5030
rect 118056 4966 118108 4972
rect 117412 3732 117464 3738
rect 117412 3674 117464 3680
rect 117320 3596 117372 3602
rect 117320 3538 117372 3544
rect 116676 3528 116728 3534
rect 116676 3470 116728 3476
rect 117516 3194 117544 4966
rect 117872 4480 117924 4486
rect 117872 4422 117924 4428
rect 117596 3460 117648 3466
rect 117596 3402 117648 3408
rect 117504 3188 117556 3194
rect 117504 3130 117556 3136
rect 116308 3120 116360 3126
rect 116308 3062 116360 3068
rect 117320 2984 117372 2990
rect 117320 2926 117372 2932
rect 116216 2440 116268 2446
rect 116216 2382 116268 2388
rect 115664 1624 115716 1630
rect 115664 1566 115716 1572
rect 116124 1488 116176 1494
rect 116124 1430 116176 1436
rect 116136 1018 116164 1430
rect 117332 1358 117360 2926
rect 117504 2372 117556 2378
rect 117504 2314 117556 2320
rect 117320 1352 117372 1358
rect 117320 1294 117372 1300
rect 117516 1290 117544 2314
rect 117504 1284 117556 1290
rect 117504 1226 117556 1232
rect 112352 1012 112404 1018
rect 112352 954 112404 960
rect 116124 1012 116176 1018
rect 116124 954 116176 960
rect 111800 740 111852 746
rect 111800 682 111852 688
rect 117608 678 117636 3402
rect 117884 3058 117912 4422
rect 117872 3052 117924 3058
rect 117872 2994 117924 3000
rect 118068 2854 118096 4966
rect 118424 4480 118476 4486
rect 118424 4422 118476 4428
rect 118148 4072 118200 4078
rect 118148 4014 118200 4020
rect 118056 2848 118108 2854
rect 118056 2790 118108 2796
rect 118068 2446 118096 2790
rect 117872 2440 117924 2446
rect 117872 2382 117924 2388
rect 118056 2440 118108 2446
rect 118056 2382 118108 2388
rect 117884 1358 117912 2382
rect 117872 1352 117924 1358
rect 117872 1294 117924 1300
rect 118160 1154 118188 4014
rect 118436 3602 118464 4422
rect 118424 3596 118476 3602
rect 118424 3538 118476 3544
rect 118712 3126 118740 5510
rect 118804 3534 118832 5578
rect 118976 4480 119028 4486
rect 118976 4422 119028 4428
rect 118988 4146 119016 4422
rect 118976 4140 119028 4146
rect 118976 4082 119028 4088
rect 119160 4004 119212 4010
rect 119160 3946 119212 3952
rect 118792 3528 118844 3534
rect 118792 3470 118844 3476
rect 119172 3466 119200 3946
rect 119356 3942 119384 5578
rect 119528 4480 119580 4486
rect 119528 4422 119580 4428
rect 119344 3936 119396 3942
rect 119344 3878 119396 3884
rect 119356 3534 119384 3878
rect 119344 3528 119396 3534
rect 119344 3470 119396 3476
rect 119160 3460 119212 3466
rect 119160 3402 119212 3408
rect 118700 3120 118752 3126
rect 118700 3062 118752 3068
rect 119540 3058 119568 4422
rect 120092 3534 120120 5714
rect 120080 3528 120132 3534
rect 120080 3470 120132 3476
rect 119988 3460 120040 3466
rect 119988 3402 120040 3408
rect 119528 3052 119580 3058
rect 119528 2994 119580 3000
rect 118700 2372 118752 2378
rect 118700 2314 118752 2320
rect 118148 1148 118200 1154
rect 118148 1090 118200 1096
rect 117596 672 117648 678
rect 117596 614 117648 620
rect 67568 248 67580 304
rect 67636 248 67660 304
rect 67716 248 67740 304
rect 67796 248 67820 304
rect 67876 248 67888 304
rect 118712 270 118740 2314
rect 120000 1086 120028 3402
rect 120276 3126 120304 6054
rect 123852 5908 123904 5914
rect 123852 5850 123904 5856
rect 120632 4616 120684 4622
rect 120632 4558 120684 4564
rect 120644 4146 120672 4558
rect 120724 4480 120776 4486
rect 120724 4422 120776 4428
rect 121368 4480 121420 4486
rect 121368 4422 121420 4428
rect 122380 4480 122432 4486
rect 122380 4422 122432 4428
rect 120356 4140 120408 4146
rect 120356 4082 120408 4088
rect 120632 4140 120684 4146
rect 120632 4082 120684 4088
rect 120264 3120 120316 3126
rect 120264 3062 120316 3068
rect 120172 2372 120224 2378
rect 120172 2314 120224 2320
rect 120080 2032 120132 2038
rect 120080 1974 120132 1980
rect 120092 1222 120120 1974
rect 120080 1216 120132 1222
rect 120080 1158 120132 1164
rect 119988 1080 120040 1086
rect 119988 1022 120040 1028
rect 67568 224 67888 248
rect 67568 168 67580 224
rect 67636 168 67660 224
rect 67716 168 67740 224
rect 67796 168 67820 224
rect 67876 168 67888 224
rect 118700 264 118752 270
rect 118700 206 118752 212
rect 120184 202 120212 2314
rect 120368 678 120396 4082
rect 120540 3528 120592 3534
rect 120540 3470 120592 3476
rect 120552 1494 120580 3470
rect 120644 3466 120672 4082
rect 120736 3534 120764 4422
rect 120816 3936 120868 3942
rect 120816 3878 120868 3884
rect 120724 3528 120776 3534
rect 120724 3470 120776 3476
rect 120632 3460 120684 3466
rect 120632 3402 120684 3408
rect 120828 2774 120856 3878
rect 121380 3058 121408 4422
rect 121644 4072 121696 4078
rect 121644 4014 121696 4020
rect 121368 3052 121420 3058
rect 121368 2994 121420 3000
rect 121552 2984 121604 2990
rect 121552 2926 121604 2932
rect 120644 2746 120856 2774
rect 120644 2446 120672 2746
rect 120632 2440 120684 2446
rect 120632 2382 120684 2388
rect 121460 2372 121512 2378
rect 121460 2314 121512 2320
rect 120540 1488 120592 1494
rect 120540 1430 120592 1436
rect 120356 672 120408 678
rect 120356 614 120408 620
rect 121472 474 121500 2314
rect 121460 468 121512 474
rect 121460 410 121512 416
rect 121564 338 121592 2926
rect 121656 882 121684 4014
rect 122392 3466 122420 4422
rect 122656 4072 122708 4078
rect 122656 4014 122708 4020
rect 123484 4072 123536 4078
rect 123484 4014 123536 4020
rect 121828 3460 121880 3466
rect 121828 3402 121880 3408
rect 122380 3460 122432 3466
rect 122380 3402 122432 3408
rect 121736 2916 121788 2922
rect 121736 2858 121788 2864
rect 121644 876 121696 882
rect 121644 818 121696 824
rect 121748 338 121776 2858
rect 121840 1290 121868 3402
rect 122392 2446 122420 3402
rect 122564 3392 122616 3398
rect 122564 3334 122616 3340
rect 122576 3233 122604 3334
rect 122562 3224 122618 3233
rect 122562 3159 122618 3168
rect 122576 3058 122604 3159
rect 122564 3052 122616 3058
rect 122564 2994 122616 3000
rect 122380 2440 122432 2446
rect 122380 2382 122432 2388
rect 122668 2281 122696 4014
rect 123208 3392 123260 3398
rect 123208 3334 123260 3340
rect 123220 3058 123248 3334
rect 123208 3052 123260 3058
rect 123208 2994 123260 3000
rect 122932 2984 122984 2990
rect 122932 2926 122984 2932
rect 122840 2372 122892 2378
rect 122840 2314 122892 2320
rect 122654 2272 122710 2281
rect 122654 2207 122710 2216
rect 121828 1284 121880 1290
rect 121828 1226 121880 1232
rect 122852 950 122880 2314
rect 122840 944 122892 950
rect 122840 886 122892 892
rect 122944 513 122972 2926
rect 123220 2145 123248 2994
rect 123496 2446 123524 4014
rect 123760 3460 123812 3466
rect 123760 3402 123812 3408
rect 123484 2440 123536 2446
rect 123484 2382 123536 2388
rect 123206 2136 123262 2145
rect 123206 2071 123262 2080
rect 122930 504 122986 513
rect 122930 439 122986 448
rect 121552 332 121604 338
rect 121552 274 121604 280
rect 121736 332 121788 338
rect 121736 274 121788 280
rect 67568 144 67888 168
rect 67568 88 67580 144
rect 67636 88 67660 144
rect 67716 88 67740 144
rect 67796 88 67820 144
rect 67876 88 67888 144
rect 120172 196 120224 202
rect 120172 138 120224 144
rect 67568 64 67888 88
rect 123772 66 123800 3402
rect 123864 3126 123892 5850
rect 124508 4146 124536 6870
rect 125152 4146 125180 6938
rect 124496 4140 124548 4146
rect 124496 4082 124548 4088
rect 125140 4140 125192 4146
rect 125140 4082 125192 4088
rect 123852 3120 123904 3126
rect 123852 3062 123904 3068
rect 124508 2446 124536 4082
rect 125152 3534 125180 4082
rect 125140 3528 125192 3534
rect 125140 3470 125192 3476
rect 125048 3460 125100 3466
rect 125048 3402 125100 3408
rect 125232 3460 125284 3466
rect 125232 3402 125284 3408
rect 124588 3052 124640 3058
rect 124588 2994 124640 3000
rect 124600 2854 124628 2994
rect 124588 2848 124640 2854
rect 124588 2790 124640 2796
rect 124496 2440 124548 2446
rect 124496 2382 124548 2388
rect 123852 2372 123904 2378
rect 123852 2314 123904 2320
rect 123864 814 123892 2314
rect 123852 808 123904 814
rect 123852 750 123904 756
rect 125060 610 125088 3402
rect 125244 2990 125272 3402
rect 125428 3058 125456 7142
rect 125888 3738 125916 7142
rect 126796 6860 126848 6866
rect 126796 6802 126848 6808
rect 126244 6112 126296 6118
rect 126244 6054 126296 6060
rect 125876 3732 125928 3738
rect 125876 3674 125928 3680
rect 125888 3534 125916 3674
rect 125876 3528 125928 3534
rect 125876 3470 125928 3476
rect 126256 3058 126284 6054
rect 126428 4684 126480 4690
rect 126428 4626 126480 4632
rect 126440 3738 126468 4626
rect 126612 4548 126664 4554
rect 126612 4490 126664 4496
rect 126520 4072 126572 4078
rect 126520 4014 126572 4020
rect 126532 3738 126560 4014
rect 126428 3732 126480 3738
rect 126428 3674 126480 3680
rect 126520 3732 126572 3738
rect 126520 3674 126572 3680
rect 125416 3052 125468 3058
rect 125416 2994 125468 3000
rect 126244 3052 126296 3058
rect 126244 2994 126296 3000
rect 125232 2984 125284 2990
rect 125232 2926 125284 2932
rect 126060 2916 126112 2922
rect 126060 2858 126112 2864
rect 126072 2446 126100 2858
rect 126060 2440 126112 2446
rect 126060 2382 126112 2388
rect 125232 2372 125284 2378
rect 125232 2314 125284 2320
rect 125048 604 125100 610
rect 125048 546 125100 552
rect 125244 134 125272 2314
rect 126072 1766 126100 2382
rect 126440 2378 126468 3674
rect 126624 2446 126652 4490
rect 126808 2774 126836 6802
rect 136560 6186 136588 9182
rect 153108 8968 153160 8974
rect 153108 8910 153160 8916
rect 171048 8968 171100 8974
rect 171048 8910 171100 8916
rect 153120 6186 153148 8910
rect 171060 6186 171088 8910
rect 187620 6186 187648 9182
rect 198836 9124 199156 9796
rect 198836 9068 198848 9124
rect 198904 9068 198928 9124
rect 198984 9068 199008 9124
rect 199064 9068 199088 9124
rect 199144 9068 199156 9124
rect 198836 9044 199156 9068
rect 198836 8988 198848 9044
rect 198904 8988 198928 9044
rect 198984 8988 199008 9044
rect 199064 8988 199088 9044
rect 199144 8988 199156 9044
rect 198836 8964 199156 8988
rect 198836 8908 198848 8964
rect 198904 8908 198928 8964
rect 198984 8908 199008 8964
rect 199064 8908 199088 8964
rect 199144 8908 199156 8964
rect 198836 8884 199156 8908
rect 198836 8828 198848 8884
rect 198904 8828 198928 8884
rect 198984 8828 199008 8884
rect 199064 8828 199088 8884
rect 199144 8828 199156 8884
rect 198836 7098 199156 8828
rect 198836 7046 198842 7098
rect 198894 7080 198906 7098
rect 198958 7080 198970 7098
rect 199022 7080 199034 7098
rect 199086 7080 199098 7098
rect 198904 7046 198906 7080
rect 199086 7046 199088 7080
rect 199150 7046 199156 7098
rect 198836 7024 198848 7046
rect 198904 7024 198928 7046
rect 198984 7024 199008 7046
rect 199064 7024 199088 7046
rect 199144 7024 199156 7046
rect 198836 7000 199156 7024
rect 198836 6944 198848 7000
rect 198904 6944 198928 7000
rect 198984 6944 199008 7000
rect 199064 6944 199088 7000
rect 199144 6944 199156 7000
rect 198836 6920 199156 6944
rect 198836 6864 198848 6920
rect 198904 6864 198928 6920
rect 198984 6864 199008 6920
rect 199064 6864 199088 6920
rect 199144 6864 199156 6920
rect 198836 6840 199156 6864
rect 198836 6784 198848 6840
rect 198904 6784 198928 6840
rect 198984 6784 199008 6840
rect 199064 6784 199088 6840
rect 199144 6784 199156 6840
rect 136548 6180 136600 6186
rect 136548 6122 136600 6128
rect 145840 6180 145892 6186
rect 145840 6122 145892 6128
rect 153108 6180 153160 6186
rect 153108 6122 153160 6128
rect 164148 6180 164200 6186
rect 164148 6122 164200 6128
rect 171048 6180 171100 6186
rect 171048 6122 171100 6128
rect 179420 6180 179472 6186
rect 179420 6122 179472 6128
rect 187608 6180 187660 6186
rect 187608 6122 187660 6128
rect 137284 5092 137336 5098
rect 137284 5034 137336 5040
rect 131396 4752 131448 4758
rect 131396 4694 131448 4700
rect 126888 3460 126940 3466
rect 126888 3402 126940 3408
rect 126900 2922 126928 3402
rect 127348 3120 127400 3126
rect 127348 3062 127400 3068
rect 127440 3120 127492 3126
rect 127440 3062 127492 3068
rect 126888 2916 126940 2922
rect 126888 2858 126940 2864
rect 126808 2746 126928 2774
rect 126612 2440 126664 2446
rect 126612 2382 126664 2388
rect 126428 2372 126480 2378
rect 126428 2314 126480 2320
rect 126900 2310 126928 2746
rect 126888 2304 126940 2310
rect 126888 2246 126940 2252
rect 127360 1766 127388 3062
rect 127452 2854 127480 3062
rect 127440 2848 127492 2854
rect 127440 2790 127492 2796
rect 131408 2446 131436 4694
rect 137296 2446 137324 5034
rect 143908 4616 143960 4622
rect 143908 4558 143960 4564
rect 143172 2848 143224 2854
rect 143172 2790 143224 2796
rect 143184 2582 143212 2790
rect 143172 2576 143224 2582
rect 143172 2518 143224 2524
rect 143184 2446 143212 2518
rect 143920 2446 143948 4558
rect 145852 3058 145880 6122
rect 150992 5160 151044 5166
rect 150992 5102 151044 5108
rect 145840 3052 145892 3058
rect 145840 2994 145892 3000
rect 145852 2446 145880 2994
rect 148232 2576 148284 2582
rect 148230 2544 148232 2553
rect 148284 2544 148286 2553
rect 148230 2479 148286 2488
rect 148244 2446 148272 2479
rect 131396 2440 131448 2446
rect 131396 2382 131448 2388
rect 137284 2440 137336 2446
rect 137284 2382 137336 2388
rect 143172 2440 143224 2446
rect 143172 2382 143224 2388
rect 143908 2440 143960 2446
rect 143908 2382 143960 2388
rect 145840 2440 145892 2446
rect 145840 2382 145892 2388
rect 148232 2440 148284 2446
rect 148232 2382 148284 2388
rect 151004 2378 151032 5102
rect 156696 4820 156748 4826
rect 156696 4762 156748 4768
rect 152188 2848 152240 2854
rect 152188 2790 152240 2796
rect 152200 2446 152228 2790
rect 156708 2446 156736 4762
rect 152188 2440 152240 2446
rect 152188 2382 152240 2388
rect 156696 2440 156748 2446
rect 156696 2382 156748 2388
rect 150992 2372 151044 2378
rect 150992 2314 151044 2320
rect 128820 2304 128872 2310
rect 128820 2246 128872 2252
rect 130200 2304 130252 2310
rect 130200 2246 130252 2252
rect 136088 2304 136140 2310
rect 136088 2246 136140 2252
rect 146116 2304 146168 2310
rect 146116 2246 146168 2252
rect 128832 2038 128860 2246
rect 128820 2032 128872 2038
rect 130212 2009 130240 2246
rect 128820 1974 128872 1980
rect 130198 2000 130254 2009
rect 136100 1970 136128 2246
rect 130198 1935 130254 1944
rect 136088 1964 136140 1970
rect 136088 1906 136140 1912
rect 126060 1760 126112 1766
rect 126060 1702 126112 1708
rect 127348 1760 127400 1766
rect 127348 1702 127400 1708
rect 146128 610 146156 2246
rect 146116 604 146168 610
rect 146116 546 146168 552
rect 152200 474 152228 2382
rect 154028 2372 154080 2378
rect 154028 2314 154080 2320
rect 157892 2372 157944 2378
rect 157892 2314 157944 2320
rect 161848 2372 161900 2378
rect 161848 2314 161900 2320
rect 152740 2304 152792 2310
rect 152740 2246 152792 2252
rect 152752 1562 152780 2246
rect 154040 1970 154068 2314
rect 154028 1964 154080 1970
rect 154028 1906 154080 1912
rect 152740 1556 152792 1562
rect 152740 1498 152792 1504
rect 157904 882 157932 2314
rect 160468 2304 160520 2310
rect 160468 2246 160520 2252
rect 160480 1222 160508 2246
rect 161860 1222 161888 2314
rect 164160 2310 164188 6122
rect 169208 5908 169260 5914
rect 169208 5850 169260 5856
rect 164332 3392 164384 3398
rect 164332 3334 164384 3340
rect 164344 3058 164372 3334
rect 164332 3052 164384 3058
rect 164332 2994 164384 3000
rect 168012 3052 168064 3058
rect 168012 2994 168064 3000
rect 164344 2446 164372 2994
rect 168024 2854 168052 2994
rect 169220 2990 169248 5850
rect 169208 2984 169260 2990
rect 169208 2926 169260 2932
rect 164792 2848 164844 2854
rect 164792 2790 164844 2796
rect 168012 2848 168064 2854
rect 168012 2790 168064 2796
rect 164804 2650 164832 2790
rect 164792 2644 164844 2650
rect 164792 2586 164844 2592
rect 164804 2446 164832 2586
rect 164332 2440 164384 2446
rect 164332 2382 164384 2388
rect 164792 2440 164844 2446
rect 164792 2382 164844 2388
rect 165528 2372 165580 2378
rect 165528 2314 165580 2320
rect 164148 2304 164200 2310
rect 164148 2246 164200 2252
rect 160468 1216 160520 1222
rect 160468 1158 160520 1164
rect 161848 1216 161900 1222
rect 161848 1158 161900 1164
rect 157892 876 157944 882
rect 157892 818 157944 824
rect 165540 814 165568 2314
rect 168024 1902 168052 2790
rect 179432 2650 179460 6122
rect 198836 6010 199156 6784
rect 198836 5958 198842 6010
rect 198894 5958 198906 6010
rect 198958 5958 198970 6010
rect 199022 5958 199034 6010
rect 199086 5958 199098 6010
rect 199150 5958 199156 6010
rect 198836 5721 199156 5958
rect 198836 5665 198848 5721
rect 198904 5665 198928 5721
rect 198984 5665 199008 5721
rect 199064 5665 199088 5721
rect 199144 5665 199156 5721
rect 198836 5641 199156 5665
rect 198836 5585 198848 5641
rect 198904 5585 198928 5641
rect 198984 5585 199008 5641
rect 199064 5585 199088 5641
rect 199144 5585 199156 5641
rect 198836 5561 199156 5585
rect 198836 5505 198848 5561
rect 198904 5505 198928 5561
rect 198984 5505 199008 5561
rect 199064 5505 199088 5561
rect 199144 5505 199156 5561
rect 198836 5481 199156 5505
rect 198836 5425 198848 5481
rect 198904 5425 198928 5481
rect 198984 5425 199008 5481
rect 199064 5425 199088 5481
rect 199144 5425 199156 5481
rect 198836 4922 199156 5425
rect 198836 4870 198842 4922
rect 198894 4870 198906 4922
rect 198958 4870 198970 4922
rect 199022 4870 199034 4922
rect 199086 4870 199098 4922
rect 199150 4870 199156 4922
rect 198836 4362 199156 4870
rect 198836 4306 198848 4362
rect 198904 4306 198928 4362
rect 198984 4306 199008 4362
rect 199064 4306 199088 4362
rect 199144 4306 199156 4362
rect 198836 4282 199156 4306
rect 198836 4226 198848 4282
rect 198904 4226 198928 4282
rect 198984 4226 199008 4282
rect 199064 4226 199088 4282
rect 199144 4226 199156 4282
rect 192208 4208 192260 4214
rect 192208 4150 192260 4156
rect 198836 4202 199156 4226
rect 179420 2644 179472 2650
rect 179420 2586 179472 2592
rect 192220 2446 192248 4150
rect 198836 4146 198848 4202
rect 198904 4146 198928 4202
rect 198984 4146 199008 4202
rect 199064 4146 199088 4202
rect 199144 4146 199156 4202
rect 198836 4122 199156 4146
rect 198836 4066 198848 4122
rect 198904 4066 198928 4122
rect 198984 4066 199008 4122
rect 199064 4066 199088 4122
rect 199144 4066 199156 4122
rect 198836 3834 199156 4066
rect 198836 3782 198842 3834
rect 198894 3782 198906 3834
rect 198958 3782 198970 3834
rect 199022 3782 199034 3834
rect 199086 3782 199098 3834
rect 199150 3782 199156 3834
rect 198836 3003 199156 3782
rect 198836 2947 198848 3003
rect 198904 2947 198928 3003
rect 198984 2947 199008 3003
rect 199064 2947 199088 3003
rect 199144 2947 199156 3003
rect 198836 2923 199156 2947
rect 198836 2867 198848 2923
rect 198904 2867 198928 2923
rect 198984 2867 199008 2923
rect 199064 2867 199088 2923
rect 199144 2867 199156 2923
rect 198836 2843 199156 2867
rect 198836 2787 198848 2843
rect 198904 2787 198928 2843
rect 198984 2787 199008 2843
rect 199064 2787 199088 2843
rect 199144 2787 199156 2843
rect 198836 2763 199156 2787
rect 198836 2746 198848 2763
rect 198904 2746 198928 2763
rect 198984 2746 199008 2763
rect 199064 2746 199088 2763
rect 199144 2746 199156 2763
rect 198836 2694 198842 2746
rect 198904 2707 198906 2746
rect 199086 2707 199088 2746
rect 198894 2694 198906 2707
rect 198958 2694 198970 2707
rect 199022 2694 199034 2707
rect 199086 2694 199098 2707
rect 199150 2694 199156 2746
rect 192208 2440 192260 2446
rect 192208 2382 192260 2388
rect 169024 2372 169076 2378
rect 169024 2314 169076 2320
rect 168012 1896 168064 1902
rect 168012 1838 168064 1844
rect 165528 808 165580 814
rect 165528 750 165580 756
rect 169036 746 169064 2314
rect 170772 2304 170824 2310
rect 170772 2246 170824 2252
rect 182916 2304 182968 2310
rect 182916 2246 182968 2252
rect 193588 2304 193640 2310
rect 193588 2246 193640 2252
rect 197912 2304 197964 2310
rect 197912 2246 197964 2252
rect 169024 740 169076 746
rect 169024 682 169076 688
rect 152188 468 152240 474
rect 152188 410 152240 416
rect 170784 406 170812 2246
rect 182928 1154 182956 2246
rect 182916 1148 182968 1154
rect 182916 1090 182968 1096
rect 193600 542 193628 2246
rect 197924 1018 197952 2246
rect 197912 1012 197964 1018
rect 197912 954 197964 960
rect 198836 964 199156 2694
rect 199496 9784 199816 9796
rect 199496 9728 199508 9784
rect 199564 9728 199588 9784
rect 199644 9728 199668 9784
rect 199724 9728 199748 9784
rect 199804 9728 199816 9784
rect 199496 9704 199816 9728
rect 199496 9648 199508 9704
rect 199564 9648 199588 9704
rect 199644 9648 199668 9704
rect 199724 9648 199748 9704
rect 199804 9648 199816 9704
rect 199496 9624 199816 9648
rect 199496 9568 199508 9624
rect 199564 9568 199588 9624
rect 199644 9568 199668 9624
rect 199724 9568 199748 9624
rect 199804 9568 199816 9624
rect 199496 9544 199816 9568
rect 199496 9488 199508 9544
rect 199564 9488 199588 9544
rect 199644 9488 199668 9544
rect 199724 9488 199748 9544
rect 199804 9488 199816 9544
rect 199496 7740 199816 9488
rect 204168 9240 204220 9246
rect 204168 9182 204220 9188
rect 222108 9240 222160 9246
rect 222108 9182 222160 9188
rect 273168 9240 273220 9246
rect 273168 9182 273220 9188
rect 289452 9240 289504 9246
rect 289452 9182 289504 9188
rect 199496 7684 199508 7740
rect 199564 7684 199588 7740
rect 199644 7684 199668 7740
rect 199724 7684 199748 7740
rect 199804 7684 199816 7740
rect 199496 7660 199816 7684
rect 199496 7642 199508 7660
rect 199564 7642 199588 7660
rect 199644 7642 199668 7660
rect 199724 7642 199748 7660
rect 199804 7642 199816 7660
rect 199496 7590 199502 7642
rect 199564 7604 199566 7642
rect 199746 7604 199748 7642
rect 199554 7590 199566 7604
rect 199618 7590 199630 7604
rect 199682 7590 199694 7604
rect 199746 7590 199758 7604
rect 199810 7590 199816 7642
rect 199496 7580 199816 7590
rect 199496 7524 199508 7580
rect 199564 7524 199588 7580
rect 199644 7524 199668 7580
rect 199724 7524 199748 7580
rect 199804 7524 199816 7580
rect 199496 7500 199816 7524
rect 199496 7444 199508 7500
rect 199564 7444 199588 7500
rect 199644 7444 199668 7500
rect 199724 7444 199748 7500
rect 199804 7444 199816 7500
rect 199496 6554 199816 7444
rect 202788 7268 202840 7274
rect 202788 7210 202840 7216
rect 199496 6502 199502 6554
rect 199554 6502 199566 6554
rect 199618 6502 199630 6554
rect 199682 6502 199694 6554
rect 199746 6502 199758 6554
rect 199810 6502 199816 6554
rect 199496 6381 199816 6502
rect 199496 6325 199508 6381
rect 199564 6325 199588 6381
rect 199644 6325 199668 6381
rect 199724 6325 199748 6381
rect 199804 6325 199816 6381
rect 199496 6301 199816 6325
rect 199496 6245 199508 6301
rect 199564 6245 199588 6301
rect 199644 6245 199668 6301
rect 199724 6245 199748 6301
rect 199804 6245 199816 6301
rect 199496 6221 199816 6245
rect 199496 6165 199508 6221
rect 199564 6165 199588 6221
rect 199644 6165 199668 6221
rect 199724 6165 199748 6221
rect 199804 6165 199816 6221
rect 199496 6141 199816 6165
rect 199496 6085 199508 6141
rect 199564 6085 199588 6141
rect 199644 6085 199668 6141
rect 199724 6085 199748 6141
rect 199804 6085 199816 6141
rect 200212 6180 200264 6186
rect 200212 6122 200264 6128
rect 199496 5466 199816 6085
rect 199496 5414 199502 5466
rect 199554 5414 199566 5466
rect 199618 5414 199630 5466
rect 199682 5414 199694 5466
rect 199746 5414 199758 5466
rect 199810 5414 199816 5466
rect 199496 5022 199816 5414
rect 199496 4966 199508 5022
rect 199564 4966 199588 5022
rect 199644 4966 199668 5022
rect 199724 4966 199748 5022
rect 199804 4966 199816 5022
rect 199496 4942 199816 4966
rect 199496 4886 199508 4942
rect 199564 4886 199588 4942
rect 199644 4886 199668 4942
rect 199724 4886 199748 4942
rect 199804 4886 199816 4942
rect 199496 4862 199816 4886
rect 199496 4806 199508 4862
rect 199564 4806 199588 4862
rect 199644 4806 199668 4862
rect 199724 4806 199748 4862
rect 199804 4806 199816 4862
rect 199496 4782 199816 4806
rect 199496 4726 199508 4782
rect 199564 4726 199588 4782
rect 199644 4726 199668 4782
rect 199724 4726 199748 4782
rect 199804 4726 199816 4782
rect 199496 4378 199816 4726
rect 199496 4326 199502 4378
rect 199554 4326 199566 4378
rect 199618 4326 199630 4378
rect 199682 4326 199694 4378
rect 199746 4326 199758 4378
rect 199810 4326 199816 4378
rect 199496 3663 199816 4326
rect 199496 3607 199508 3663
rect 199564 3607 199588 3663
rect 199644 3607 199668 3663
rect 199724 3607 199748 3663
rect 199804 3607 199816 3663
rect 199496 3583 199816 3607
rect 199496 3527 199508 3583
rect 199564 3527 199588 3583
rect 199644 3527 199668 3583
rect 199724 3527 199748 3583
rect 199804 3527 199816 3583
rect 199496 3503 199816 3527
rect 199496 3447 199508 3503
rect 199564 3447 199588 3503
rect 199644 3447 199668 3503
rect 199724 3447 199748 3503
rect 199804 3447 199816 3503
rect 199496 3423 199816 3447
rect 199496 3367 199508 3423
rect 199564 3367 199588 3423
rect 199644 3367 199668 3423
rect 199724 3367 199748 3423
rect 199804 3367 199816 3423
rect 199496 3290 199816 3367
rect 199496 3238 199502 3290
rect 199554 3238 199566 3290
rect 199618 3238 199630 3290
rect 199682 3238 199694 3290
rect 199746 3238 199758 3290
rect 199810 3238 199816 3290
rect 199384 2372 199436 2378
rect 199384 2314 199436 2320
rect 199396 1018 199424 2314
rect 199496 2202 199816 3238
rect 200224 2446 200252 6122
rect 200948 4072 201000 4078
rect 200948 4014 201000 4020
rect 200960 3670 200988 4014
rect 200948 3664 201000 3670
rect 200948 3606 201000 3612
rect 202800 3058 202828 7210
rect 204180 6186 204208 9182
rect 218520 7472 218572 7478
rect 218520 7414 218572 7420
rect 217140 6996 217192 7002
rect 217140 6938 217192 6944
rect 218060 6996 218112 7002
rect 218060 6938 218112 6944
rect 208584 6248 208636 6254
rect 208584 6190 208636 6196
rect 209412 6248 209464 6254
rect 209412 6190 209464 6196
rect 204168 6180 204220 6186
rect 204168 6122 204220 6128
rect 207664 5840 207716 5846
rect 207664 5782 207716 5788
rect 204904 5228 204956 5234
rect 204904 5170 204956 5176
rect 203892 4208 203944 4214
rect 203892 4150 203944 4156
rect 201684 3052 201736 3058
rect 201684 2994 201736 3000
rect 202788 3052 202840 3058
rect 202788 2994 202840 3000
rect 201696 2854 201724 2994
rect 201684 2848 201736 2854
rect 201684 2790 201736 2796
rect 200212 2440 200264 2446
rect 201696 2417 201724 2790
rect 203904 2446 203932 4150
rect 204916 2990 204944 5170
rect 206192 3052 206244 3058
rect 206192 2994 206244 3000
rect 206836 3052 206888 3058
rect 206836 2994 206888 3000
rect 204904 2984 204956 2990
rect 204904 2926 204956 2932
rect 206204 2854 206232 2994
rect 206848 2854 206876 2994
rect 206192 2848 206244 2854
rect 206192 2790 206244 2796
rect 206836 2848 206888 2854
rect 206836 2790 206888 2796
rect 203892 2440 203944 2446
rect 200212 2382 200264 2388
rect 201682 2408 201738 2417
rect 203892 2382 203944 2388
rect 201682 2343 201738 2352
rect 206100 2372 206152 2378
rect 206100 2314 206152 2320
rect 200396 2304 200448 2310
rect 200396 2246 200448 2252
rect 202696 2304 202748 2310
rect 202696 2246 202748 2252
rect 204904 2304 204956 2310
rect 204904 2246 204956 2252
rect 199496 2150 199502 2202
rect 199554 2150 199566 2202
rect 199618 2150 199630 2202
rect 199682 2150 199694 2202
rect 199746 2150 199758 2202
rect 199810 2150 199816 2202
rect 198836 908 198848 964
rect 198904 908 198928 964
rect 198984 908 199008 964
rect 199064 908 199088 964
rect 199144 908 199156 964
rect 199384 1012 199436 1018
rect 199384 954 199436 960
rect 198836 884 199156 908
rect 198836 828 198848 884
rect 198904 828 198928 884
rect 198984 828 199008 884
rect 199064 828 199088 884
rect 199144 828 199156 884
rect 198836 804 199156 828
rect 198836 748 198848 804
rect 198904 748 198928 804
rect 198984 748 199008 804
rect 199064 748 199088 804
rect 199144 748 199156 804
rect 198836 724 199156 748
rect 198836 668 198848 724
rect 198904 668 198928 724
rect 198984 668 199008 724
rect 199064 668 199088 724
rect 199144 668 199156 724
rect 193588 536 193640 542
rect 193588 478 193640 484
rect 170772 400 170824 406
rect 170772 342 170824 348
rect 125232 128 125284 134
rect 125232 70 125284 76
rect 67568 8 67580 64
rect 67636 8 67660 64
rect 67716 8 67740 64
rect 67796 8 67820 64
rect 67876 8 67888 64
rect 67568 -4 67888 8
rect 123760 60 123812 66
rect 123760 2 123812 8
rect 198836 -4 199156 668
rect 199496 304 199816 2150
rect 200408 1902 200436 2246
rect 202708 2106 202736 2246
rect 202696 2100 202748 2106
rect 202696 2042 202748 2048
rect 200396 1896 200448 1902
rect 200396 1838 200448 1844
rect 204916 610 204944 2246
rect 206112 1562 206140 2314
rect 206100 1556 206152 1562
rect 206100 1498 206152 1504
rect 206204 610 206232 2790
rect 206848 1698 206876 2790
rect 207676 2446 207704 5782
rect 208400 5568 208452 5574
rect 208400 5510 208452 5516
rect 208124 4276 208176 4282
rect 208124 4218 208176 4224
rect 208136 2990 208164 4218
rect 208412 3942 208440 5510
rect 208400 3936 208452 3942
rect 208400 3878 208452 3884
rect 208492 3936 208544 3942
rect 208492 3878 208544 3884
rect 208124 2984 208176 2990
rect 208124 2926 208176 2932
rect 208412 2446 208440 3878
rect 208504 3534 208532 3878
rect 208492 3528 208544 3534
rect 208492 3470 208544 3476
rect 208596 2990 208624 6190
rect 209044 5840 209096 5846
rect 209044 5782 209096 5788
rect 208860 5704 208912 5710
rect 208860 5646 208912 5652
rect 208872 3534 208900 5646
rect 209056 4146 209084 5782
rect 208952 4140 209004 4146
rect 208952 4082 209004 4088
rect 209044 4140 209096 4146
rect 209044 4082 209096 4088
rect 208860 3528 208912 3534
rect 208860 3470 208912 3476
rect 208964 3466 208992 4082
rect 209056 3534 209084 4082
rect 209044 3528 209096 3534
rect 209044 3470 209096 3476
rect 208952 3460 209004 3466
rect 208952 3402 209004 3408
rect 208584 2984 208636 2990
rect 208584 2926 208636 2932
rect 209424 2446 209452 6190
rect 212816 5772 212868 5778
rect 212816 5714 212868 5720
rect 209596 5704 209648 5710
rect 209596 5646 209648 5652
rect 209608 3942 209636 5646
rect 210792 5024 210844 5030
rect 210792 4966 210844 4972
rect 211620 5024 211672 5030
rect 211620 4966 211672 4972
rect 210424 4480 210476 4486
rect 210424 4422 210476 4428
rect 210436 4010 210464 4422
rect 210424 4004 210476 4010
rect 210424 3946 210476 3952
rect 209596 3936 209648 3942
rect 209596 3878 209648 3884
rect 209608 3058 209636 3878
rect 210240 3188 210292 3194
rect 210240 3130 210292 3136
rect 209596 3052 209648 3058
rect 209596 2994 209648 3000
rect 210252 2990 210280 3130
rect 210804 3058 210832 4966
rect 211528 4820 211580 4826
rect 211528 4762 211580 4768
rect 211068 4480 211120 4486
rect 211068 4422 211120 4428
rect 211080 4146 211108 4422
rect 211540 4282 211568 4762
rect 211528 4276 211580 4282
rect 211528 4218 211580 4224
rect 211068 4140 211120 4146
rect 211068 4082 211120 4088
rect 210792 3052 210844 3058
rect 210792 2994 210844 3000
rect 210240 2984 210292 2990
rect 210240 2926 210292 2932
rect 207664 2440 207716 2446
rect 207664 2382 207716 2388
rect 208400 2440 208452 2446
rect 208400 2382 208452 2388
rect 209412 2440 209464 2446
rect 209412 2382 209464 2388
rect 208860 2372 208912 2378
rect 208860 2314 208912 2320
rect 210240 2372 210292 2378
rect 210240 2314 210292 2320
rect 206836 1692 206888 1698
rect 206836 1634 206888 1640
rect 208400 1692 208452 1698
rect 208400 1634 208452 1640
rect 204904 604 204956 610
rect 204904 546 204956 552
rect 206192 604 206244 610
rect 206192 546 206244 552
rect 208412 474 208440 1634
rect 208872 1630 208900 2314
rect 208860 1624 208912 1630
rect 208860 1566 208912 1572
rect 210252 1358 210280 2314
rect 210240 1352 210292 1358
rect 210240 1294 210292 1300
rect 210804 950 210832 2994
rect 211080 1086 211108 4082
rect 211436 2984 211488 2990
rect 211436 2926 211488 2932
rect 211068 1080 211120 1086
rect 211068 1022 211120 1028
rect 210792 944 210844 950
rect 210792 886 210844 892
rect 211448 678 211476 2926
rect 211528 2440 211580 2446
rect 211528 2382 211580 2388
rect 211540 1902 211568 2382
rect 211632 2378 211660 4966
rect 211712 4480 211764 4486
rect 211712 4422 211764 4428
rect 212172 4480 212224 4486
rect 212172 4422 212224 4428
rect 211724 3670 211752 4422
rect 211712 3664 211764 3670
rect 211712 3606 211764 3612
rect 211724 3466 211752 3606
rect 212184 3534 212212 4422
rect 212828 4146 212856 5714
rect 213368 5636 213420 5642
rect 213368 5578 213420 5584
rect 213184 4480 213236 4486
rect 213184 4422 213236 4428
rect 212816 4140 212868 4146
rect 212868 4100 212948 4128
rect 212816 4082 212868 4088
rect 212540 3936 212592 3942
rect 212540 3878 212592 3884
rect 212172 3528 212224 3534
rect 212172 3470 212224 3476
rect 211712 3460 211764 3466
rect 211712 3402 211764 3408
rect 211804 2644 211856 2650
rect 211804 2586 211856 2592
rect 211816 2514 211844 2586
rect 211804 2508 211856 2514
rect 211804 2450 211856 2456
rect 211620 2372 211672 2378
rect 211620 2314 211672 2320
rect 211528 1896 211580 1902
rect 211528 1838 211580 1844
rect 212184 1834 212212 3470
rect 212552 2990 212580 3878
rect 212920 3534 212948 4100
rect 212908 3528 212960 3534
rect 212908 3470 212960 3476
rect 212632 3460 212684 3466
rect 212632 3402 212684 3408
rect 212540 2984 212592 2990
rect 212540 2926 212592 2932
rect 212448 2372 212500 2378
rect 212448 2314 212500 2320
rect 212172 1828 212224 1834
rect 212172 1770 212224 1776
rect 212460 678 212488 2314
rect 211436 672 211488 678
rect 211436 614 211488 620
rect 212448 672 212500 678
rect 212448 614 212500 620
rect 208400 468 208452 474
rect 208400 410 208452 416
rect 212644 338 212672 3402
rect 213196 3058 213224 4422
rect 213380 4146 213408 5578
rect 213644 5228 213696 5234
rect 213644 5170 213696 5176
rect 213552 4480 213604 4486
rect 213552 4422 213604 4428
rect 213368 4140 213420 4146
rect 213368 4082 213420 4088
rect 213564 3058 213592 4422
rect 213184 3052 213236 3058
rect 213184 2994 213236 3000
rect 213552 3052 213604 3058
rect 213552 2994 213604 3000
rect 212816 2372 212868 2378
rect 212816 2314 212868 2320
rect 212828 1494 212856 2314
rect 213196 1630 213224 2994
rect 213564 2417 213592 2994
rect 213656 2446 213684 5170
rect 214472 5160 214524 5166
rect 214472 5102 214524 5108
rect 214288 5024 214340 5030
rect 214288 4966 214340 4972
rect 213920 4480 213972 4486
rect 213920 4422 213972 4428
rect 213932 4146 213960 4422
rect 213920 4140 213972 4146
rect 213920 4082 213972 4088
rect 213644 2440 213696 2446
rect 213550 2408 213606 2417
rect 213644 2382 213696 2388
rect 213550 2343 213606 2352
rect 213184 1624 213236 1630
rect 213184 1566 213236 1572
rect 213932 1494 213960 4082
rect 214300 3913 214328 4966
rect 214484 4554 214512 5102
rect 214840 5024 214892 5030
rect 214840 4966 214892 4972
rect 215392 5024 215444 5030
rect 215392 4966 215444 4972
rect 216220 5024 216272 5030
rect 216220 4966 216272 4972
rect 216864 5024 216916 5030
rect 216864 4966 216916 4972
rect 214472 4548 214524 4554
rect 214472 4490 214524 4496
rect 214286 3904 214342 3913
rect 214286 3839 214342 3848
rect 214012 3460 214064 3466
rect 214012 3402 214064 3408
rect 214024 2922 214052 3402
rect 214012 2916 214064 2922
rect 214012 2858 214064 2864
rect 214300 2446 214328 3839
rect 214852 3466 214880 4966
rect 215208 4480 215260 4486
rect 215208 4422 215260 4428
rect 214932 4072 214984 4078
rect 214932 4014 214984 4020
rect 214840 3460 214892 3466
rect 214840 3402 214892 3408
rect 214944 2514 214972 4014
rect 215220 3534 215248 4422
rect 215208 3528 215260 3534
rect 215208 3470 215260 3476
rect 214932 2508 214984 2514
rect 214932 2450 214984 2456
rect 214288 2440 214340 2446
rect 214288 2382 214340 2388
rect 214012 2372 214064 2378
rect 214012 2314 214064 2320
rect 214024 2281 214052 2314
rect 214010 2272 214066 2281
rect 214010 2207 214066 2216
rect 212816 1488 212868 1494
rect 212816 1430 212868 1436
rect 213920 1488 213972 1494
rect 213920 1430 213972 1436
rect 215220 1290 215248 3470
rect 215404 3194 215432 4966
rect 215484 4548 215536 4554
rect 215484 4490 215536 4496
rect 215496 4146 215524 4490
rect 215484 4140 215536 4146
rect 215484 4082 215536 4088
rect 215852 3460 215904 3466
rect 215852 3402 215904 3408
rect 215392 3188 215444 3194
rect 215392 3130 215444 3136
rect 215392 2372 215444 2378
rect 215392 2314 215444 2320
rect 215404 2145 215432 2314
rect 215390 2136 215446 2145
rect 215390 2071 215446 2080
rect 215208 1284 215260 1290
rect 215208 1226 215260 1232
rect 199496 248 199508 304
rect 199564 248 199588 304
rect 199644 248 199668 304
rect 199724 248 199748 304
rect 199804 248 199816 304
rect 212632 332 212684 338
rect 212632 274 212684 280
rect 199496 224 199816 248
rect 199496 168 199508 224
rect 199564 168 199588 224
rect 199644 168 199668 224
rect 199724 168 199748 224
rect 199804 168 199816 224
rect 215864 202 215892 3402
rect 216232 3058 216260 4966
rect 216772 4480 216824 4486
rect 216772 4422 216824 4428
rect 216680 4072 216732 4078
rect 216680 4014 216732 4020
rect 216588 3732 216640 3738
rect 216588 3674 216640 3680
rect 216600 3126 216628 3674
rect 216692 3233 216720 4014
rect 216678 3224 216734 3233
rect 216678 3159 216734 3168
rect 216588 3120 216640 3126
rect 216588 3062 216640 3068
rect 216220 3052 216272 3058
rect 216220 2994 216272 3000
rect 216784 2446 216812 4422
rect 216876 2514 216904 4966
rect 216956 4140 217008 4146
rect 216956 4082 217008 4088
rect 216968 3942 216996 4082
rect 216956 3936 217008 3942
rect 216956 3878 217008 3884
rect 217152 3534 217180 6938
rect 217416 6180 217468 6186
rect 217416 6122 217468 6128
rect 217324 4548 217376 4554
rect 217324 4490 217376 4496
rect 217232 4480 217284 4486
rect 217232 4422 217284 4428
rect 217140 3528 217192 3534
rect 217140 3470 217192 3476
rect 217244 3466 217272 4422
rect 217336 4146 217364 4490
rect 217324 4140 217376 4146
rect 217324 4082 217376 4088
rect 217232 3460 217284 3466
rect 217232 3402 217284 3408
rect 217428 2774 217456 6122
rect 217968 4480 218020 4486
rect 217968 4422 218020 4428
rect 217980 3058 218008 4422
rect 218072 3942 218100 6938
rect 218152 5228 218204 5234
rect 218152 5170 218204 5176
rect 218164 4078 218192 5170
rect 218152 4072 218204 4078
rect 218152 4014 218204 4020
rect 218532 3942 218560 7414
rect 219532 7404 219584 7410
rect 219532 7346 219584 7352
rect 218704 7200 218756 7206
rect 218704 7142 218756 7148
rect 218060 3936 218112 3942
rect 218060 3878 218112 3884
rect 218520 3936 218572 3942
rect 218520 3878 218572 3884
rect 218532 3534 218560 3878
rect 218520 3528 218572 3534
rect 218520 3470 218572 3476
rect 218716 3058 218744 7142
rect 218888 6928 218940 6934
rect 218888 6870 218940 6876
rect 218900 3534 218928 6870
rect 219164 6112 219216 6118
rect 219164 6054 219216 6060
rect 218888 3528 218940 3534
rect 218888 3470 218940 3476
rect 217968 3052 218020 3058
rect 217968 2994 218020 3000
rect 218704 3052 218756 3058
rect 218704 2994 218756 3000
rect 218428 2848 218480 2854
rect 218428 2790 218480 2796
rect 217428 2746 218008 2774
rect 216864 2508 216916 2514
rect 216864 2450 216916 2456
rect 216680 2440 216732 2446
rect 216680 2382 216732 2388
rect 216772 2440 216824 2446
rect 216772 2382 216824 2388
rect 216588 2372 216640 2378
rect 216588 2314 216640 2320
rect 216600 1766 216628 2314
rect 216588 1760 216640 1766
rect 216588 1702 216640 1708
rect 216692 1426 216720 2382
rect 217980 2310 218008 2746
rect 218440 2446 218468 2790
rect 219176 2514 219204 6054
rect 219544 3942 219572 7346
rect 220452 7336 220504 7342
rect 220452 7278 220504 7284
rect 220360 5160 220412 5166
rect 220360 5102 220412 5108
rect 219900 4684 219952 4690
rect 219900 4626 219952 4632
rect 219532 3936 219584 3942
rect 219532 3878 219584 3884
rect 219624 3936 219676 3942
rect 219624 3878 219676 3884
rect 219544 3058 219572 3878
rect 219636 3534 219664 3878
rect 219716 3664 219768 3670
rect 219716 3606 219768 3612
rect 219728 3534 219756 3606
rect 219624 3528 219676 3534
rect 219624 3470 219676 3476
rect 219716 3528 219768 3534
rect 219716 3470 219768 3476
rect 219912 3126 219940 4626
rect 220084 4480 220136 4486
rect 220084 4422 220136 4428
rect 220096 4214 220124 4422
rect 220084 4208 220136 4214
rect 220084 4150 220136 4156
rect 220004 3466 220216 3482
rect 219992 3460 220216 3466
rect 220044 3454 220216 3460
rect 219992 3402 220044 3408
rect 220188 3398 220216 3454
rect 220176 3392 220228 3398
rect 220176 3334 220228 3340
rect 219900 3120 219952 3126
rect 219900 3062 219952 3068
rect 219532 3052 219584 3058
rect 219532 2994 219584 3000
rect 219164 2508 219216 2514
rect 219164 2450 219216 2456
rect 220372 2446 220400 5102
rect 220464 3942 220492 7278
rect 222120 6186 222148 9182
rect 238668 8968 238720 8974
rect 238668 8910 238720 8916
rect 238680 6186 238708 8910
rect 255228 8900 255280 8906
rect 255228 8842 255280 8848
rect 255240 6186 255268 8842
rect 273180 6186 273208 9182
rect 289464 6186 289492 9182
rect 330764 9124 331084 9796
rect 330764 9068 330776 9124
rect 330832 9068 330856 9124
rect 330912 9068 330936 9124
rect 330992 9068 331016 9124
rect 331072 9068 331084 9124
rect 330764 9044 331084 9068
rect 330764 8988 330776 9044
rect 330832 8988 330856 9044
rect 330912 8988 330936 9044
rect 330992 8988 331016 9044
rect 331072 8988 331084 9044
rect 306288 8968 306340 8974
rect 306288 8910 306340 8916
rect 324228 8968 324280 8974
rect 324228 8910 324280 8916
rect 330764 8964 331084 8988
rect 302884 8492 302936 8498
rect 302884 8434 302936 8440
rect 293776 8424 293828 8430
rect 293776 8366 293828 8372
rect 291108 7200 291160 7206
rect 291108 7142 291160 7148
rect 222108 6180 222160 6186
rect 222108 6122 222160 6128
rect 236276 6180 236328 6186
rect 236276 6122 236328 6128
rect 238668 6180 238720 6186
rect 238668 6122 238720 6128
rect 254032 6180 254084 6186
rect 254032 6122 254084 6128
rect 255228 6180 255280 6186
rect 255228 6122 255280 6128
rect 271788 6180 271840 6186
rect 271788 6122 271840 6128
rect 273168 6180 273220 6186
rect 273168 6122 273220 6128
rect 288348 6180 288400 6186
rect 288348 6122 288400 6128
rect 289452 6180 289504 6186
rect 289452 6122 289504 6128
rect 230756 5092 230808 5098
rect 230756 5034 230808 5040
rect 221096 5024 221148 5030
rect 221096 4966 221148 4972
rect 221004 4684 221056 4690
rect 221004 4626 221056 4632
rect 220452 3936 220504 3942
rect 220452 3878 220504 3884
rect 220464 3738 220492 3878
rect 220452 3732 220504 3738
rect 220452 3674 220504 3680
rect 220544 3732 220596 3738
rect 220544 3674 220596 3680
rect 220556 3194 220584 3674
rect 220636 3664 220688 3670
rect 220636 3606 220688 3612
rect 220648 3398 220676 3606
rect 220636 3392 220688 3398
rect 220636 3334 220688 3340
rect 220544 3188 220596 3194
rect 220544 3130 220596 3136
rect 221016 2446 221044 4626
rect 221108 3194 221136 4966
rect 224960 4752 225012 4758
rect 224960 4694 225012 4700
rect 221096 3188 221148 3194
rect 221096 3130 221148 3136
rect 221188 3188 221240 3194
rect 221188 3130 221240 3136
rect 221200 2922 221228 3130
rect 221372 3052 221424 3058
rect 221372 2994 221424 3000
rect 221188 2916 221240 2922
rect 221188 2858 221240 2864
rect 218428 2440 218480 2446
rect 218428 2382 218480 2388
rect 220360 2440 220412 2446
rect 220360 2382 220412 2388
rect 221004 2440 221056 2446
rect 221004 2382 221056 2388
rect 217968 2304 218020 2310
rect 217968 2246 218020 2252
rect 216680 1420 216732 1426
rect 216680 1362 216732 1368
rect 218440 270 218468 2382
rect 221384 2310 221412 2994
rect 221648 2848 221700 2854
rect 221648 2790 221700 2796
rect 221660 2514 221688 2790
rect 221648 2508 221700 2514
rect 221648 2450 221700 2456
rect 224972 2446 225000 4694
rect 230768 2446 230796 5034
rect 224960 2440 225012 2446
rect 224960 2382 225012 2388
rect 230756 2440 230808 2446
rect 230756 2382 230808 2388
rect 223028 2372 223080 2378
rect 223028 2314 223080 2320
rect 226156 2372 226208 2378
rect 226156 2314 226208 2320
rect 231952 2372 232004 2378
rect 231952 2314 232004 2320
rect 221372 2304 221424 2310
rect 221372 2246 221424 2252
rect 223040 2038 223068 2314
rect 224224 2304 224276 2310
rect 224224 2246 224276 2252
rect 224236 2145 224264 2246
rect 224222 2136 224278 2145
rect 226168 2106 226196 2314
rect 224222 2071 224278 2080
rect 226156 2100 226208 2106
rect 226156 2042 226208 2048
rect 231964 2038 231992 2314
rect 236288 2310 236316 6122
rect 239036 5160 239088 5166
rect 239036 5102 239088 5108
rect 237748 4616 237800 4622
rect 237748 4558 237800 4564
rect 237760 2446 237788 4558
rect 239048 2446 239076 5102
rect 254044 3058 254072 6122
rect 262312 5908 262364 5914
rect 262312 5850 262364 5856
rect 263508 5908 263560 5914
rect 263508 5850 263560 5856
rect 260012 4752 260064 4758
rect 260012 4694 260064 4700
rect 259092 3392 259144 3398
rect 259092 3334 259144 3340
rect 259104 3058 259132 3334
rect 254032 3052 254084 3058
rect 254032 2994 254084 3000
rect 259092 3052 259144 3058
rect 259092 2994 259144 3000
rect 247132 2848 247184 2854
rect 247132 2790 247184 2796
rect 251732 2848 251784 2854
rect 251732 2790 251784 2796
rect 247144 2446 247172 2790
rect 251744 2446 251772 2790
rect 254044 2446 254072 2994
rect 260024 2446 260052 4694
rect 260288 3052 260340 3058
rect 260288 2994 260340 3000
rect 260300 2854 260328 2994
rect 260288 2848 260340 2854
rect 260288 2790 260340 2796
rect 237748 2440 237800 2446
rect 237748 2382 237800 2388
rect 239036 2440 239088 2446
rect 239036 2382 239088 2388
rect 247132 2440 247184 2446
rect 247132 2382 247184 2388
rect 251732 2440 251784 2446
rect 251732 2382 251784 2388
rect 254032 2440 254084 2446
rect 254032 2382 254084 2388
rect 255780 2440 255832 2446
rect 255780 2382 255832 2388
rect 260012 2440 260064 2446
rect 260012 2382 260064 2388
rect 244188 2372 244240 2378
rect 244188 2314 244240 2320
rect 246304 2372 246356 2378
rect 246304 2314 246356 2320
rect 236276 2304 236328 2310
rect 236276 2246 236328 2252
rect 237012 2304 237064 2310
rect 237012 2246 237064 2252
rect 223028 2032 223080 2038
rect 223028 1974 223080 1980
rect 231952 2032 232004 2038
rect 231952 1974 232004 1980
rect 237024 1086 237052 2246
rect 244200 1902 244228 2314
rect 244188 1896 244240 1902
rect 244188 1838 244240 1844
rect 246316 1698 246344 2314
rect 246304 1692 246356 1698
rect 246304 1634 246356 1640
rect 237012 1080 237064 1086
rect 237012 1022 237064 1028
rect 247144 338 247172 2382
rect 248052 2304 248104 2310
rect 248052 2246 248104 2252
rect 248064 1970 248092 2246
rect 248052 1964 248104 1970
rect 248052 1906 248104 1912
rect 251744 882 251772 2382
rect 255792 2310 255820 2382
rect 257068 2372 257120 2378
rect 257068 2314 257120 2320
rect 254308 2304 254360 2310
rect 254308 2246 254360 2252
rect 255780 2304 255832 2310
rect 255780 2246 255832 2252
rect 254320 882 254348 2246
rect 255792 1222 255820 2246
rect 255780 1216 255832 1222
rect 255780 1158 255832 1164
rect 251732 876 251784 882
rect 251732 818 251784 824
rect 254308 876 254360 882
rect 254308 818 254360 824
rect 257080 746 257108 2314
rect 258264 2304 258316 2310
rect 258264 2246 258316 2252
rect 258356 2304 258408 2310
rect 258356 2246 258408 2252
rect 257068 740 257120 746
rect 257068 682 257120 688
rect 258276 474 258304 2246
rect 258368 814 258396 2246
rect 260300 2009 260328 2790
rect 262324 2446 262352 5850
rect 263520 2446 263548 5850
rect 262312 2440 262364 2446
rect 262312 2382 262364 2388
rect 263508 2440 263560 2446
rect 263508 2382 263560 2388
rect 264336 2372 264388 2378
rect 264336 2314 264388 2320
rect 260286 2000 260342 2009
rect 260286 1935 260342 1944
rect 258356 808 258408 814
rect 258356 750 258408 756
rect 258264 468 258316 474
rect 258264 410 258316 416
rect 264348 406 264376 2314
rect 271800 2310 271828 6122
rect 287428 4548 287480 4554
rect 287428 4490 287480 4496
rect 273076 4208 273128 4214
rect 273076 4150 273128 4156
rect 273088 2446 273116 4150
rect 287440 2446 287468 4490
rect 273076 2440 273128 2446
rect 273076 2382 273128 2388
rect 287428 2440 287480 2446
rect 287428 2382 287480 2388
rect 277124 2372 277176 2378
rect 277124 2314 277176 2320
rect 285956 2372 286008 2378
rect 285956 2314 286008 2320
rect 265716 2304 265768 2310
rect 265716 2246 265768 2252
rect 271788 2304 271840 2310
rect 271788 2246 271840 2252
rect 265728 814 265756 2246
rect 277136 1154 277164 2314
rect 278320 2304 278372 2310
rect 278320 2246 278372 2252
rect 277124 1148 277176 1154
rect 277124 1090 277176 1096
rect 265716 808 265768 814
rect 265716 750 265768 756
rect 278332 406 278360 2246
rect 285968 542 285996 2314
rect 288360 2310 288388 6122
rect 291120 2514 291148 7142
rect 293788 2514 293816 8366
rect 300216 7404 300268 7410
rect 300216 7346 300268 7352
rect 296536 7268 296588 7274
rect 296536 7210 296588 7216
rect 295432 5024 295484 5030
rect 295432 4966 295484 4972
rect 291108 2508 291160 2514
rect 291108 2450 291160 2456
rect 293776 2508 293828 2514
rect 293776 2450 293828 2456
rect 295444 2446 295472 4966
rect 296548 3058 296576 7210
rect 298652 5636 298704 5642
rect 298652 5578 298704 5584
rect 297364 4276 297416 4282
rect 297364 4218 297416 4224
rect 297376 3058 297404 4218
rect 298664 3058 298692 5578
rect 300228 3058 300256 7346
rect 301412 7336 301464 7342
rect 301412 7278 301464 7284
rect 300860 6316 300912 6322
rect 300860 6258 300912 6264
rect 300872 3466 300900 6258
rect 301136 4820 301188 4826
rect 301136 4762 301188 4768
rect 300860 3460 300912 3466
rect 300860 3402 300912 3408
rect 300308 3392 300360 3398
rect 300308 3334 300360 3340
rect 296536 3052 296588 3058
rect 296536 2994 296588 3000
rect 297364 3052 297416 3058
rect 297364 2994 297416 3000
rect 298652 3052 298704 3058
rect 298652 2994 298704 3000
rect 300216 3052 300268 3058
rect 300216 2994 300268 3000
rect 295800 2848 295852 2854
rect 295800 2790 295852 2796
rect 292580 2440 292632 2446
rect 292580 2382 292632 2388
rect 295432 2440 295484 2446
rect 295432 2382 295484 2388
rect 292592 2310 292620 2382
rect 295812 2378 295840 2790
rect 296548 2446 296576 2994
rect 296994 2544 297050 2553
rect 296994 2479 297050 2488
rect 297008 2446 297036 2479
rect 298664 2446 298692 2994
rect 299572 2848 299624 2854
rect 299572 2790 299624 2796
rect 299584 2446 299612 2790
rect 300320 2446 300348 3334
rect 300872 3058 300900 3402
rect 301148 3058 301176 4762
rect 300860 3052 300912 3058
rect 300860 2994 300912 3000
rect 301136 3052 301188 3058
rect 301136 2994 301188 3000
rect 301228 3052 301280 3058
rect 301228 2994 301280 3000
rect 301148 2854 301176 2994
rect 301240 2922 301268 2994
rect 301228 2916 301280 2922
rect 301228 2858 301280 2864
rect 301136 2848 301188 2854
rect 301136 2790 301188 2796
rect 301424 2650 301452 7278
rect 302792 3392 302844 3398
rect 302792 3334 302844 3340
rect 301412 2644 301464 2650
rect 301412 2586 301464 2592
rect 302804 2582 302832 3334
rect 302896 2650 302924 8434
rect 303436 7268 303488 7274
rect 303436 7210 303488 7216
rect 303448 3534 303476 7210
rect 304724 6928 304776 6934
rect 304724 6870 304776 6876
rect 303804 5840 303856 5846
rect 303804 5782 303856 5788
rect 303436 3528 303488 3534
rect 303436 3470 303488 3476
rect 303448 3058 303476 3470
rect 303436 3052 303488 3058
rect 303436 2994 303488 3000
rect 303816 2990 303844 5782
rect 304172 4480 304224 4486
rect 304172 4422 304224 4428
rect 304184 4078 304212 4422
rect 304172 4072 304224 4078
rect 304172 4014 304224 4020
rect 303988 3936 304040 3942
rect 303988 3878 304040 3884
rect 304000 3534 304028 3878
rect 303988 3528 304040 3534
rect 303988 3470 304040 3476
rect 303804 2984 303856 2990
rect 303804 2926 303856 2932
rect 302884 2644 302936 2650
rect 302884 2586 302936 2592
rect 302792 2576 302844 2582
rect 302792 2518 302844 2524
rect 302804 2446 302832 2518
rect 304184 2446 304212 4014
rect 304356 3052 304408 3058
rect 304356 2994 304408 3000
rect 304368 2854 304396 2994
rect 304356 2848 304408 2854
rect 304356 2790 304408 2796
rect 304736 2650 304764 6870
rect 306104 6248 306156 6254
rect 306104 6190 306156 6196
rect 305000 6180 305052 6186
rect 305000 6122 305052 6128
rect 304816 6112 304868 6118
rect 304816 6054 304868 6060
rect 304828 4078 304856 6054
rect 304816 4072 304868 4078
rect 304816 4014 304868 4020
rect 304828 3534 304856 4014
rect 304816 3528 304868 3534
rect 304816 3470 304868 3476
rect 304724 2644 304776 2650
rect 304724 2586 304776 2592
rect 296536 2440 296588 2446
rect 296536 2382 296588 2388
rect 296996 2440 297048 2446
rect 296996 2382 297048 2388
rect 298652 2440 298704 2446
rect 298652 2382 298704 2388
rect 299572 2440 299624 2446
rect 299572 2382 299624 2388
rect 300308 2440 300360 2446
rect 300308 2382 300360 2388
rect 302792 2440 302844 2446
rect 302792 2382 302844 2388
rect 304172 2440 304224 2446
rect 304172 2382 304224 2388
rect 295800 2372 295852 2378
rect 295800 2314 295852 2320
rect 299020 2372 299072 2378
rect 299020 2314 299072 2320
rect 288348 2304 288400 2310
rect 288348 2246 288400 2252
rect 292580 2304 292632 2310
rect 292580 2246 292632 2252
rect 292592 1018 292620 2246
rect 292580 1012 292632 1018
rect 292580 954 292632 960
rect 295812 542 295840 2314
rect 299032 610 299060 2314
rect 299584 1018 299612 2382
rect 300320 1562 300348 2382
rect 300768 2372 300820 2378
rect 300768 2314 300820 2320
rect 303988 2372 304040 2378
rect 303988 2314 304040 2320
rect 300780 2281 300808 2314
rect 300766 2272 300822 2281
rect 300766 2207 300822 2216
rect 304000 1873 304028 2314
rect 305012 2310 305040 6122
rect 305276 5704 305328 5710
rect 305276 5646 305328 5652
rect 305184 4072 305236 4078
rect 305184 4014 305236 4020
rect 305000 2304 305052 2310
rect 305000 2246 305052 2252
rect 303986 1864 304042 1873
rect 303986 1799 304042 1808
rect 300308 1556 300360 1562
rect 300308 1498 300360 1504
rect 299572 1012 299624 1018
rect 299572 954 299624 960
rect 305196 950 305224 4014
rect 305288 3534 305316 5646
rect 305368 5568 305420 5574
rect 305368 5510 305420 5516
rect 305276 3528 305328 3534
rect 305276 3470 305328 3476
rect 305380 2990 305408 5510
rect 306012 5024 306064 5030
rect 306012 4966 306064 4972
rect 305552 4480 305604 4486
rect 305552 4422 305604 4428
rect 305460 3936 305512 3942
rect 305460 3878 305512 3884
rect 305368 2984 305420 2990
rect 305368 2926 305420 2932
rect 305472 2854 305500 3878
rect 305564 3534 305592 4422
rect 305552 3528 305604 3534
rect 305552 3470 305604 3476
rect 305460 2848 305512 2854
rect 305460 2790 305512 2796
rect 305472 2514 305500 2790
rect 305460 2508 305512 2514
rect 305460 2450 305512 2456
rect 305460 2372 305512 2378
rect 305460 2314 305512 2320
rect 305184 944 305236 950
rect 305184 886 305236 892
rect 305472 678 305500 2314
rect 305564 1698 305592 3470
rect 306024 2446 306052 4966
rect 306116 3534 306144 6190
rect 306300 6186 306328 8910
rect 308404 8356 308456 8362
rect 308404 8298 308456 8304
rect 306656 7472 306708 7478
rect 306656 7414 306708 7420
rect 306288 6180 306340 6186
rect 306288 6122 306340 6128
rect 306196 4480 306248 4486
rect 306196 4422 306248 4428
rect 306380 4480 306432 4486
rect 306380 4422 306432 4428
rect 306104 3528 306156 3534
rect 306104 3470 306156 3476
rect 306208 3058 306236 4422
rect 306392 3516 306420 4422
rect 306472 4140 306524 4146
rect 306472 4082 306524 4088
rect 306564 4140 306616 4146
rect 306564 4082 306616 4088
rect 306484 3942 306512 4082
rect 306472 3936 306524 3942
rect 306472 3878 306524 3884
rect 306472 3528 306524 3534
rect 306392 3488 306472 3516
rect 306472 3470 306524 3476
rect 306196 3052 306248 3058
rect 306196 2994 306248 3000
rect 306208 2774 306236 2994
rect 306116 2746 306236 2774
rect 306012 2440 306064 2446
rect 306012 2382 306064 2388
rect 305552 1692 305604 1698
rect 305552 1634 305604 1640
rect 306024 1290 306052 2382
rect 306116 1562 306144 2746
rect 306196 2100 306248 2106
rect 306196 2042 306248 2048
rect 306104 1556 306156 1562
rect 306104 1498 306156 1504
rect 306012 1284 306064 1290
rect 306012 1226 306064 1232
rect 306208 1222 306236 2042
rect 306484 2038 306512 3470
rect 306576 3058 306604 4082
rect 306564 3052 306616 3058
rect 306564 2994 306616 3000
rect 306668 2922 306696 7414
rect 308128 5772 308180 5778
rect 308128 5714 308180 5720
rect 306748 5024 306800 5030
rect 306748 4966 306800 4972
rect 307576 5024 307628 5030
rect 307576 4966 307628 4972
rect 307852 5024 307904 5030
rect 307852 4966 307904 4972
rect 306656 2916 306708 2922
rect 306656 2858 306708 2864
rect 306760 2446 306788 4966
rect 306840 4480 306892 4486
rect 306840 4422 306892 4428
rect 306852 3058 306880 4422
rect 307024 3936 307076 3942
rect 307024 3878 307076 3884
rect 306840 3052 306892 3058
rect 306840 2994 306892 3000
rect 306748 2440 306800 2446
rect 306748 2382 306800 2388
rect 306288 2032 306340 2038
rect 306288 1974 306340 1980
rect 306472 2032 306524 2038
rect 306472 1974 306524 1980
rect 306300 1358 306328 1974
rect 306288 1352 306340 1358
rect 306288 1294 306340 1300
rect 306196 1216 306248 1222
rect 306196 1158 306248 1164
rect 306760 882 306788 2382
rect 307036 1766 307064 3878
rect 307588 3466 307616 4966
rect 307760 4616 307812 4622
rect 307760 4558 307812 4564
rect 307668 4480 307720 4486
rect 307668 4422 307720 4428
rect 307680 4146 307708 4422
rect 307668 4140 307720 4146
rect 307668 4082 307720 4088
rect 307668 3936 307720 3942
rect 307668 3878 307720 3884
rect 307116 3460 307168 3466
rect 307116 3402 307168 3408
rect 307576 3460 307628 3466
rect 307576 3402 307628 3408
rect 307128 1834 307156 3402
rect 307392 3392 307444 3398
rect 307392 3334 307444 3340
rect 307404 3126 307432 3334
rect 307392 3120 307444 3126
rect 307392 3062 307444 3068
rect 307392 2984 307444 2990
rect 307392 2926 307444 2932
rect 307300 2372 307352 2378
rect 307300 2314 307352 2320
rect 307116 1828 307168 1834
rect 307116 1770 307168 1776
rect 307024 1760 307076 1766
rect 307024 1702 307076 1708
rect 306748 876 306800 882
rect 306748 818 306800 824
rect 307312 678 307340 2314
rect 307404 1630 307432 2926
rect 307392 1624 307444 1630
rect 307392 1566 307444 1572
rect 305460 672 305512 678
rect 305460 614 305512 620
rect 307300 672 307352 678
rect 307300 614 307352 620
rect 299020 604 299072 610
rect 299020 546 299072 552
rect 285956 536 286008 542
rect 285956 478 286008 484
rect 295800 536 295852 542
rect 307680 513 307708 3878
rect 307772 2854 307800 4558
rect 307864 3058 307892 4966
rect 308140 3534 308168 5714
rect 308128 3528 308180 3534
rect 308128 3470 308180 3476
rect 307852 3052 307904 3058
rect 307852 2994 307904 3000
rect 307760 2848 307812 2854
rect 307760 2790 307812 2796
rect 307864 2106 307892 2994
rect 308416 2650 308444 8298
rect 319628 7540 319680 7546
rect 319628 7482 319680 7488
rect 314752 7472 314804 7478
rect 314752 7414 314804 7420
rect 310704 7336 310756 7342
rect 310704 7278 310756 7284
rect 308496 5092 308548 5098
rect 308496 5034 308548 5040
rect 308508 4826 308536 5034
rect 308588 5024 308640 5030
rect 308588 4966 308640 4972
rect 308496 4820 308548 4826
rect 308496 4762 308548 4768
rect 308496 3664 308548 3670
rect 308496 3606 308548 3612
rect 308508 2990 308536 3606
rect 308600 3058 308628 4966
rect 309232 4480 309284 4486
rect 309232 4422 309284 4428
rect 309600 4480 309652 4486
rect 309600 4422 309652 4428
rect 310428 4480 310480 4486
rect 310428 4422 310480 4428
rect 309244 4078 309272 4422
rect 308680 4072 308732 4078
rect 308680 4014 308732 4020
rect 309232 4072 309284 4078
rect 309232 4014 309284 4020
rect 308692 3670 308720 4014
rect 308680 3664 308732 3670
rect 308680 3606 308732 3612
rect 309244 3534 309272 4014
rect 309612 3534 309640 4422
rect 310440 4146 310468 4422
rect 309692 4140 309744 4146
rect 309692 4082 309744 4088
rect 310428 4140 310480 4146
rect 310428 4082 310480 4088
rect 310612 4140 310664 4146
rect 310612 4082 310664 4088
rect 309704 3942 309732 4082
rect 309692 3936 309744 3942
rect 309692 3878 309744 3884
rect 309784 3936 309836 3942
rect 309784 3878 309836 3884
rect 309704 3670 309732 3878
rect 309692 3664 309744 3670
rect 309692 3606 309744 3612
rect 309232 3528 309284 3534
rect 309232 3470 309284 3476
rect 309600 3528 309652 3534
rect 309600 3470 309652 3476
rect 309796 3466 309824 3878
rect 309784 3460 309836 3466
rect 309784 3402 309836 3408
rect 309416 3392 309468 3398
rect 309416 3334 309468 3340
rect 309428 3126 309456 3334
rect 309416 3120 309468 3126
rect 309416 3062 309468 3068
rect 308588 3052 308640 3058
rect 308588 2994 308640 3000
rect 308496 2984 308548 2990
rect 308496 2926 308548 2932
rect 308600 2650 308628 2994
rect 309048 2848 309100 2854
rect 309048 2790 309100 2796
rect 308404 2644 308456 2650
rect 308404 2586 308456 2592
rect 308588 2644 308640 2650
rect 308588 2586 308640 2592
rect 309060 2582 309088 2790
rect 309048 2576 309100 2582
rect 309048 2518 309100 2524
rect 309232 2372 309284 2378
rect 309232 2314 309284 2320
rect 307852 2100 307904 2106
rect 307852 2042 307904 2048
rect 307760 1896 307812 1902
rect 307760 1838 307812 1844
rect 307772 950 307800 1838
rect 309244 1494 309272 2314
rect 309232 1488 309284 1494
rect 309232 1430 309284 1436
rect 307760 944 307812 950
rect 307760 886 307812 892
rect 295800 478 295852 484
rect 307666 504 307722 513
rect 307666 439 307722 448
rect 264336 400 264388 406
rect 264336 342 264388 348
rect 278320 400 278372 406
rect 278320 342 278372 348
rect 247132 332 247184 338
rect 247132 274 247184 280
rect 218428 264 218480 270
rect 218428 206 218480 212
rect 310440 202 310468 4082
rect 310624 4010 310652 4082
rect 310716 4010 310744 7278
rect 314292 6996 314344 7002
rect 314292 6938 314344 6944
rect 314016 4684 314068 4690
rect 314016 4626 314068 4632
rect 311440 4140 311492 4146
rect 311440 4082 311492 4088
rect 310612 4004 310664 4010
rect 310612 3946 310664 3952
rect 310704 4004 310756 4010
rect 310704 3946 310756 3952
rect 311452 3942 311480 4082
rect 311348 3936 311400 3942
rect 310886 3904 310942 3913
rect 311348 3878 311400 3884
rect 311440 3936 311492 3942
rect 311440 3878 311492 3884
rect 310886 3839 310942 3848
rect 310704 3732 310756 3738
rect 310704 3674 310756 3680
rect 310716 3126 310744 3674
rect 310900 3534 310928 3839
rect 310888 3528 310940 3534
rect 310888 3470 310940 3476
rect 311164 3528 311216 3534
rect 311164 3470 311216 3476
rect 311176 3194 311204 3470
rect 311164 3188 311216 3194
rect 311164 3130 311216 3136
rect 310704 3120 310756 3126
rect 310704 3062 310756 3068
rect 310900 2514 311204 2530
rect 310888 2508 311216 2514
rect 310940 2502 311164 2508
rect 310888 2450 310940 2456
rect 311164 2450 311216 2456
rect 310612 2440 310664 2446
rect 310704 2440 310756 2446
rect 310612 2382 310664 2388
rect 310702 2408 310704 2417
rect 310756 2408 310758 2417
rect 310624 2310 310652 2382
rect 310702 2343 310758 2352
rect 311360 2310 311388 3878
rect 312728 3732 312780 3738
rect 312728 3674 312780 3680
rect 312268 3392 312320 3398
rect 312268 3334 312320 3340
rect 312280 2582 312308 3334
rect 312740 3058 312768 3674
rect 314028 3058 314056 4626
rect 312728 3052 312780 3058
rect 312728 2994 312780 3000
rect 314016 3052 314068 3058
rect 314016 2994 314068 3000
rect 313372 2848 313424 2854
rect 313372 2790 313424 2796
rect 312268 2576 312320 2582
rect 312268 2518 312320 2524
rect 313188 2576 313240 2582
rect 313188 2518 313240 2524
rect 310612 2304 310664 2310
rect 310612 2246 310664 2252
rect 311348 2304 311400 2310
rect 311348 2246 311400 2252
rect 311532 2304 311584 2310
rect 311532 2246 311584 2252
rect 311360 1834 311388 2246
rect 311348 1828 311400 1834
rect 311348 1770 311400 1776
rect 311544 1426 311572 2246
rect 313200 1902 313228 2518
rect 313280 2372 313332 2378
rect 313280 2314 313332 2320
rect 313188 1896 313240 1902
rect 313188 1838 313240 1844
rect 311532 1420 311584 1426
rect 311532 1362 311584 1368
rect 313292 270 313320 2314
rect 313384 2310 313412 2790
rect 314304 2650 314332 6938
rect 314764 3194 314792 7414
rect 315948 7404 316000 7410
rect 315948 7346 316000 7352
rect 314660 3188 314712 3194
rect 314660 3130 314712 3136
rect 314752 3188 314804 3194
rect 314752 3130 314804 3136
rect 314292 2644 314344 2650
rect 314292 2586 314344 2592
rect 313372 2304 313424 2310
rect 314672 2292 314700 3130
rect 315764 2984 315816 2990
rect 315764 2926 315816 2932
rect 315776 2378 315804 2926
rect 315960 2446 315988 7346
rect 318340 6996 318392 7002
rect 318340 6938 318392 6944
rect 317880 4276 317932 4282
rect 317880 4218 317932 4224
rect 316776 4004 316828 4010
rect 316776 3946 316828 3952
rect 316788 3466 316816 3946
rect 316776 3460 316828 3466
rect 316776 3402 316828 3408
rect 317892 3194 317920 4218
rect 317880 3188 317932 3194
rect 317880 3130 317932 3136
rect 317892 3058 317920 3130
rect 317880 3052 317932 3058
rect 317880 2994 317932 3000
rect 318352 2650 318380 6938
rect 318984 2848 319036 2854
rect 318984 2790 319036 2796
rect 319444 2848 319496 2854
rect 319444 2790 319496 2796
rect 318340 2644 318392 2650
rect 318340 2586 318392 2592
rect 318352 2446 318380 2586
rect 318996 2446 319024 2790
rect 319456 2446 319484 2790
rect 319640 2650 319668 7482
rect 324240 6254 324268 8910
rect 330764 8908 330776 8964
rect 330832 8908 330856 8964
rect 330912 8908 330936 8964
rect 330992 8908 331016 8964
rect 331072 8908 331084 8964
rect 330764 8884 331084 8908
rect 330764 8828 330776 8884
rect 330832 8828 330856 8884
rect 330912 8828 330936 8884
rect 330992 8828 331016 8884
rect 331072 8828 331084 8884
rect 330764 7098 331084 8828
rect 330764 7046 330770 7098
rect 330822 7080 330834 7098
rect 330886 7080 330898 7098
rect 330950 7080 330962 7098
rect 331014 7080 331026 7098
rect 330832 7046 330834 7080
rect 331014 7046 331016 7080
rect 331078 7046 331084 7098
rect 330764 7024 330776 7046
rect 330832 7024 330856 7046
rect 330912 7024 330936 7046
rect 330992 7024 331016 7046
rect 331072 7024 331084 7046
rect 330764 7000 331084 7024
rect 330764 6944 330776 7000
rect 330832 6944 330856 7000
rect 330912 6944 330936 7000
rect 330992 6944 331016 7000
rect 331072 6944 331084 7000
rect 330764 6920 331084 6944
rect 330764 6864 330776 6920
rect 330832 6864 330856 6920
rect 330912 6864 330936 6920
rect 330992 6864 331016 6920
rect 331072 6864 331084 6920
rect 330764 6840 331084 6864
rect 330764 6784 330776 6840
rect 330832 6784 330856 6840
rect 330912 6784 330936 6840
rect 330992 6784 331016 6840
rect 331072 6784 331084 6840
rect 324228 6248 324280 6254
rect 324228 6190 324280 6196
rect 326436 6180 326488 6186
rect 326436 6122 326488 6128
rect 325332 4684 325384 4690
rect 325332 4626 325384 4632
rect 319996 3664 320048 3670
rect 319996 3606 320048 3612
rect 319628 2644 319680 2650
rect 319628 2586 319680 2592
rect 319720 2644 319772 2650
rect 319720 2586 319772 2592
rect 315948 2440 316000 2446
rect 315948 2382 316000 2388
rect 316592 2440 316644 2446
rect 316592 2382 316644 2388
rect 318340 2440 318392 2446
rect 318340 2382 318392 2388
rect 318984 2440 319036 2446
rect 318984 2382 319036 2388
rect 319444 2440 319496 2446
rect 319444 2382 319496 2388
rect 315764 2372 315816 2378
rect 315764 2314 315816 2320
rect 314752 2304 314804 2310
rect 314672 2264 314752 2292
rect 313372 2246 313424 2252
rect 314752 2246 314804 2252
rect 313384 882 313412 2246
rect 313372 876 313424 882
rect 313372 818 313424 824
rect 313280 264 313332 270
rect 313280 206 313332 212
rect 199496 144 199816 168
rect 199496 88 199508 144
rect 199564 88 199588 144
rect 199644 88 199668 144
rect 199724 88 199748 144
rect 199804 88 199816 144
rect 215852 196 215904 202
rect 215852 138 215904 144
rect 310428 196 310480 202
rect 310428 138 310480 144
rect 199496 64 199816 88
rect 315776 66 315804 2314
rect 316604 2106 316632 2382
rect 317052 2372 317104 2378
rect 317052 2314 317104 2320
rect 317064 2145 317092 2314
rect 317050 2136 317106 2145
rect 316592 2100 316644 2106
rect 317050 2071 317106 2080
rect 316592 2042 316644 2048
rect 318996 1154 319024 2382
rect 319456 1222 319484 2382
rect 319732 2378 319760 2586
rect 319720 2372 319772 2378
rect 319720 2314 319772 2320
rect 320008 1766 320036 3606
rect 324504 3596 324556 3602
rect 324504 3538 324556 3544
rect 323400 2984 323452 2990
rect 323400 2926 323452 2932
rect 323412 2310 323440 2926
rect 323768 2848 323820 2854
rect 323768 2790 323820 2796
rect 323780 2310 323808 2790
rect 324516 2310 324544 3538
rect 324688 2848 324740 2854
rect 324688 2790 324740 2796
rect 325148 2848 325200 2854
rect 325148 2790 325200 2796
rect 324700 2446 324728 2790
rect 325160 2446 325188 2790
rect 325344 2582 325372 4626
rect 325240 2576 325292 2582
rect 325240 2518 325292 2524
rect 325332 2576 325384 2582
rect 325332 2518 325384 2524
rect 325424 2576 325476 2582
rect 325424 2518 325476 2524
rect 324688 2440 324740 2446
rect 324688 2382 324740 2388
rect 325148 2440 325200 2446
rect 325148 2382 325200 2388
rect 323400 2304 323452 2310
rect 323400 2246 323452 2252
rect 323768 2304 323820 2310
rect 323768 2246 323820 2252
rect 324504 2304 324556 2310
rect 324504 2246 324556 2252
rect 319996 1760 320048 1766
rect 319996 1702 320048 1708
rect 323780 1222 323808 2246
rect 319444 1216 319496 1222
rect 319444 1158 319496 1164
rect 323768 1216 323820 1222
rect 323768 1158 323820 1164
rect 318984 1148 319036 1154
rect 318984 1090 319036 1096
rect 324700 610 324728 2382
rect 325160 1358 325188 2382
rect 325252 2292 325280 2518
rect 325436 2292 325464 2518
rect 326448 2310 326476 6122
rect 330764 6010 331084 6784
rect 330764 5958 330770 6010
rect 330822 5958 330834 6010
rect 330886 5958 330898 6010
rect 330950 5958 330962 6010
rect 331014 5958 331026 6010
rect 331078 5958 331084 6010
rect 330764 5721 331084 5958
rect 330764 5665 330776 5721
rect 330832 5665 330856 5721
rect 330912 5665 330936 5721
rect 330992 5665 331016 5721
rect 331072 5665 331084 5721
rect 330764 5641 331084 5665
rect 330764 5585 330776 5641
rect 330832 5585 330856 5641
rect 330912 5585 330936 5641
rect 330992 5585 331016 5641
rect 331072 5585 331084 5641
rect 327172 5568 327224 5574
rect 327172 5510 327224 5516
rect 330764 5561 331084 5585
rect 327184 2446 327212 5510
rect 330764 5505 330776 5561
rect 330832 5505 330856 5561
rect 330912 5505 330936 5561
rect 330992 5505 331016 5561
rect 331072 5505 331084 5561
rect 330764 5481 331084 5505
rect 330764 5425 330776 5481
rect 330832 5425 330856 5481
rect 330912 5425 330936 5481
rect 330992 5425 331016 5481
rect 331072 5425 331084 5481
rect 330764 4922 331084 5425
rect 330764 4870 330770 4922
rect 330822 4870 330834 4922
rect 330886 4870 330898 4922
rect 330950 4870 330962 4922
rect 331014 4870 331026 4922
rect 331078 4870 331084 4922
rect 330024 4616 330076 4622
rect 330024 4558 330076 4564
rect 330036 2446 330064 4558
rect 330764 4362 331084 4870
rect 330764 4306 330776 4362
rect 330832 4306 330856 4362
rect 330912 4306 330936 4362
rect 330992 4306 331016 4362
rect 331072 4306 331084 4362
rect 330764 4282 331084 4306
rect 330764 4226 330776 4282
rect 330832 4226 330856 4282
rect 330912 4226 330936 4282
rect 330992 4226 331016 4282
rect 331072 4226 331084 4282
rect 330764 4202 331084 4226
rect 330764 4146 330776 4202
rect 330832 4146 330856 4202
rect 330912 4146 330936 4202
rect 330992 4146 331016 4202
rect 331072 4146 331084 4202
rect 330764 4122 331084 4146
rect 330764 4066 330776 4122
rect 330832 4066 330856 4122
rect 330912 4066 330936 4122
rect 330992 4066 331016 4122
rect 331072 4066 331084 4122
rect 330764 3834 331084 4066
rect 330764 3782 330770 3834
rect 330822 3782 330834 3834
rect 330886 3782 330898 3834
rect 330950 3782 330962 3834
rect 331014 3782 331026 3834
rect 331078 3782 331084 3834
rect 330764 3003 331084 3782
rect 331424 9784 331744 9796
rect 331424 9728 331436 9784
rect 331492 9728 331516 9784
rect 331572 9728 331596 9784
rect 331652 9728 331676 9784
rect 331732 9728 331744 9784
rect 331424 9704 331744 9728
rect 331424 9648 331436 9704
rect 331492 9648 331516 9704
rect 331572 9648 331596 9704
rect 331652 9648 331676 9704
rect 331732 9648 331744 9704
rect 331424 9624 331744 9648
rect 331424 9568 331436 9624
rect 331492 9568 331516 9624
rect 331572 9568 331596 9624
rect 331652 9568 331676 9624
rect 331732 9568 331744 9624
rect 331424 9544 331744 9568
rect 331424 9488 331436 9544
rect 331492 9488 331516 9544
rect 331572 9488 331596 9544
rect 331652 9488 331676 9544
rect 331732 9488 331744 9544
rect 331424 7740 331744 9488
rect 340788 9240 340840 9246
rect 340788 9182 340840 9188
rect 357256 9240 357308 9246
rect 357256 9182 357308 9188
rect 375288 9240 375340 9246
rect 375288 9182 375340 9188
rect 426348 9240 426400 9246
rect 426348 9182 426400 9188
rect 442908 9240 442960 9246
rect 442908 9182 442960 9188
rect 331424 7684 331436 7740
rect 331492 7684 331516 7740
rect 331572 7684 331596 7740
rect 331652 7684 331676 7740
rect 331732 7684 331744 7740
rect 331424 7660 331744 7684
rect 331424 7642 331436 7660
rect 331492 7642 331516 7660
rect 331572 7642 331596 7660
rect 331652 7642 331676 7660
rect 331732 7642 331744 7660
rect 331424 7590 331430 7642
rect 331492 7604 331494 7642
rect 331674 7604 331676 7642
rect 331482 7590 331494 7604
rect 331546 7590 331558 7604
rect 331610 7590 331622 7604
rect 331674 7590 331686 7604
rect 331738 7590 331744 7642
rect 331424 7580 331744 7590
rect 331424 7524 331436 7580
rect 331492 7524 331516 7580
rect 331572 7524 331596 7580
rect 331652 7524 331676 7580
rect 331732 7524 331744 7580
rect 331424 7500 331744 7524
rect 331424 7444 331436 7500
rect 331492 7444 331516 7500
rect 331572 7444 331596 7500
rect 331652 7444 331676 7500
rect 331732 7444 331744 7500
rect 331424 6554 331744 7444
rect 331424 6502 331430 6554
rect 331482 6502 331494 6554
rect 331546 6502 331558 6554
rect 331610 6502 331622 6554
rect 331674 6502 331686 6554
rect 331738 6502 331744 6554
rect 331424 6381 331744 6502
rect 331424 6325 331436 6381
rect 331492 6325 331516 6381
rect 331572 6325 331596 6381
rect 331652 6325 331676 6381
rect 331732 6325 331744 6381
rect 331424 6301 331744 6325
rect 331424 6245 331436 6301
rect 331492 6245 331516 6301
rect 331572 6245 331596 6301
rect 331652 6245 331676 6301
rect 331732 6245 331744 6301
rect 331424 6221 331744 6245
rect 331424 6165 331436 6221
rect 331492 6165 331516 6221
rect 331572 6165 331596 6221
rect 331652 6165 331676 6221
rect 331732 6165 331744 6221
rect 340800 6186 340828 9182
rect 351920 6316 351972 6322
rect 351920 6258 351972 6264
rect 341984 6248 342036 6254
rect 341984 6190 342036 6196
rect 331424 6141 331744 6165
rect 331424 6085 331436 6141
rect 331492 6085 331516 6141
rect 331572 6085 331596 6141
rect 331652 6085 331676 6141
rect 331732 6085 331744 6141
rect 340788 6180 340840 6186
rect 340788 6122 340840 6128
rect 331424 5466 331744 6085
rect 340880 5908 340932 5914
rect 340880 5850 340932 5856
rect 338028 5772 338080 5778
rect 338028 5714 338080 5720
rect 332508 5704 332560 5710
rect 332508 5646 332560 5652
rect 331424 5414 331430 5466
rect 331482 5414 331494 5466
rect 331546 5414 331558 5466
rect 331610 5414 331622 5466
rect 331674 5414 331686 5466
rect 331738 5414 331744 5466
rect 331424 5022 331744 5414
rect 332324 5160 332376 5166
rect 332324 5102 332376 5108
rect 331424 4966 331436 5022
rect 331492 4966 331516 5022
rect 331572 4966 331596 5022
rect 331652 4966 331676 5022
rect 331732 4966 331744 5022
rect 331424 4942 331744 4966
rect 331424 4886 331436 4942
rect 331492 4886 331516 4942
rect 331572 4886 331596 4942
rect 331652 4886 331676 4942
rect 331732 4886 331744 4942
rect 331424 4862 331744 4886
rect 331424 4806 331436 4862
rect 331492 4806 331516 4862
rect 331572 4806 331596 4862
rect 331652 4806 331676 4862
rect 331732 4806 331744 4862
rect 331424 4782 331744 4806
rect 331424 4726 331436 4782
rect 331492 4726 331516 4782
rect 331572 4726 331596 4782
rect 331652 4726 331676 4782
rect 331732 4726 331744 4782
rect 331424 4378 331744 4726
rect 331424 4326 331430 4378
rect 331482 4326 331494 4378
rect 331546 4326 331558 4378
rect 331610 4326 331622 4378
rect 331674 4326 331686 4378
rect 331738 4326 331744 4378
rect 331424 3663 331744 4326
rect 331424 3607 331436 3663
rect 331492 3607 331516 3663
rect 331572 3607 331596 3663
rect 331652 3607 331676 3663
rect 331732 3607 331744 3663
rect 331312 3596 331364 3602
rect 331312 3538 331364 3544
rect 331424 3583 331744 3607
rect 331324 3194 331352 3538
rect 331424 3527 331436 3583
rect 331492 3527 331516 3583
rect 331572 3527 331596 3583
rect 331652 3527 331676 3583
rect 331732 3527 331744 3583
rect 331424 3503 331744 3527
rect 331424 3447 331436 3503
rect 331492 3447 331516 3503
rect 331572 3447 331596 3503
rect 331652 3447 331676 3503
rect 331732 3447 331744 3503
rect 331424 3423 331744 3447
rect 331424 3367 331436 3423
rect 331492 3367 331516 3423
rect 331572 3367 331596 3423
rect 331652 3367 331676 3423
rect 331732 3367 331744 3423
rect 331424 3290 331744 3367
rect 331424 3238 331430 3290
rect 331482 3238 331494 3290
rect 331546 3238 331558 3290
rect 331610 3238 331622 3290
rect 331674 3238 331686 3290
rect 331738 3238 331744 3290
rect 331312 3188 331364 3194
rect 331312 3130 331364 3136
rect 330764 2947 330776 3003
rect 330832 2947 330856 3003
rect 330912 2947 330936 3003
rect 330992 2947 331016 3003
rect 331072 2947 331084 3003
rect 330764 2923 331084 2947
rect 330764 2867 330776 2923
rect 330832 2867 330856 2923
rect 330912 2867 330936 2923
rect 330992 2867 331016 2923
rect 331072 2867 331084 2923
rect 330764 2843 331084 2867
rect 330764 2787 330776 2843
rect 330832 2787 330856 2843
rect 330912 2787 330936 2843
rect 330992 2787 331016 2843
rect 331072 2787 331084 2843
rect 330764 2763 331084 2787
rect 330764 2746 330776 2763
rect 330832 2746 330856 2763
rect 330912 2746 330936 2763
rect 330992 2746 331016 2763
rect 331072 2746 331084 2763
rect 330764 2694 330770 2746
rect 330832 2707 330834 2746
rect 331014 2707 331016 2746
rect 330822 2694 330834 2707
rect 330886 2694 330898 2707
rect 330950 2694 330962 2707
rect 331014 2694 331026 2707
rect 331078 2694 331084 2746
rect 327172 2440 327224 2446
rect 327172 2382 327224 2388
rect 330024 2440 330076 2446
rect 330024 2382 330076 2388
rect 325252 2264 325464 2292
rect 326436 2304 326488 2310
rect 326436 2246 326488 2252
rect 329288 2304 329340 2310
rect 329288 2246 329340 2252
rect 329300 1766 329328 2246
rect 329288 1760 329340 1766
rect 329288 1702 329340 1708
rect 325148 1352 325200 1358
rect 325148 1294 325200 1300
rect 330764 964 331084 2694
rect 331220 2372 331272 2378
rect 331220 2314 331272 2320
rect 331232 1086 331260 2314
rect 331424 2202 331744 3238
rect 332336 2446 332364 5102
rect 332324 2440 332376 2446
rect 332324 2382 332376 2388
rect 332520 2310 332548 5646
rect 336372 3596 336424 3602
rect 336372 3538 336424 3544
rect 332784 2848 332836 2854
rect 332784 2790 332836 2796
rect 332796 2378 332824 2790
rect 336384 2446 336412 3538
rect 337292 2848 337344 2854
rect 337292 2790 337344 2796
rect 337844 2848 337896 2854
rect 337844 2790 337896 2796
rect 336372 2440 336424 2446
rect 336372 2382 336424 2388
rect 337304 2378 337332 2790
rect 337856 2446 337884 2790
rect 337844 2440 337896 2446
rect 337844 2382 337896 2388
rect 332784 2372 332836 2378
rect 332784 2314 332836 2320
rect 335268 2372 335320 2378
rect 335268 2314 335320 2320
rect 337292 2372 337344 2378
rect 337292 2314 337344 2320
rect 332508 2304 332560 2310
rect 332508 2246 332560 2252
rect 331424 2150 331430 2202
rect 331482 2150 331494 2202
rect 331546 2150 331558 2202
rect 331610 2150 331622 2202
rect 331674 2150 331686 2202
rect 331738 2150 331744 2202
rect 331220 1080 331272 1086
rect 331220 1022 331272 1028
rect 330764 908 330776 964
rect 330832 908 330856 964
rect 330912 908 330936 964
rect 330992 908 331016 964
rect 331072 908 331084 964
rect 330764 884 331084 908
rect 330764 828 330776 884
rect 330832 828 330856 884
rect 330912 828 330936 884
rect 330992 828 331016 884
rect 331072 828 331084 884
rect 330764 804 331084 828
rect 330764 748 330776 804
rect 330832 748 330856 804
rect 330912 748 330936 804
rect 330992 748 331016 804
rect 331072 748 331084 804
rect 330764 724 331084 748
rect 330764 668 330776 724
rect 330832 668 330856 724
rect 330912 668 330936 724
rect 330992 668 331016 724
rect 331072 668 331084 724
rect 324688 604 324740 610
rect 324688 546 324740 552
rect 199496 8 199508 64
rect 199564 8 199588 64
rect 199644 8 199668 64
rect 199724 8 199748 64
rect 199804 8 199816 64
rect 199496 -4 199816 8
rect 315764 60 315816 66
rect 315764 2 315816 8
rect 330764 -4 331084 668
rect 331424 304 331744 2150
rect 332600 1488 332652 1494
rect 332600 1430 332652 1436
rect 332612 678 332640 1430
rect 332796 678 332824 2314
rect 335280 1970 335308 2314
rect 337200 2304 337252 2310
rect 337200 2246 337252 2252
rect 337212 2038 337240 2246
rect 337200 2032 337252 2038
rect 337200 1974 337252 1980
rect 335268 1964 335320 1970
rect 335268 1906 335320 1912
rect 332600 672 332652 678
rect 332600 614 332652 620
rect 332784 672 332836 678
rect 332784 614 332836 620
rect 331424 248 331436 304
rect 331492 248 331516 304
rect 331572 248 331596 304
rect 331652 248 331676 304
rect 331732 248 331744 304
rect 331424 224 331744 248
rect 331424 168 331436 224
rect 331492 168 331516 224
rect 331572 168 331596 224
rect 331652 168 331676 224
rect 331732 168 331744 224
rect 331424 144 331744 168
rect 331424 88 331436 144
rect 331492 88 331516 144
rect 331572 88 331596 144
rect 331652 88 331676 144
rect 331732 88 331744 144
rect 337304 134 337332 2314
rect 337856 950 337884 2382
rect 338040 2310 338068 5714
rect 340052 4072 340104 4078
rect 340052 4014 340104 4020
rect 340064 3194 340092 4014
rect 340052 3188 340104 3194
rect 340052 3130 340104 3136
rect 340892 2990 340920 5850
rect 340880 2984 340932 2990
rect 340880 2926 340932 2932
rect 341524 2848 341576 2854
rect 341524 2790 341576 2796
rect 341536 2446 341564 2790
rect 341524 2440 341576 2446
rect 341524 2382 341576 2388
rect 339960 2372 340012 2378
rect 339960 2314 340012 2320
rect 338028 2304 338080 2310
rect 338028 2246 338080 2252
rect 338028 1760 338080 1766
rect 338028 1702 338080 1708
rect 337844 944 337896 950
rect 337844 886 337896 892
rect 338040 542 338068 1702
rect 338028 536 338080 542
rect 338028 478 338080 484
rect 339972 338 340000 2314
rect 341536 1086 341564 2382
rect 341996 2378 342024 6190
rect 342352 5840 342404 5846
rect 342352 5782 342404 5788
rect 342168 3120 342220 3126
rect 342168 3062 342220 3068
rect 342076 2848 342128 2854
rect 342076 2790 342128 2796
rect 342088 2582 342116 2790
rect 342076 2576 342128 2582
rect 342076 2518 342128 2524
rect 342088 2446 342116 2518
rect 342180 2446 342208 3062
rect 342076 2440 342128 2446
rect 342076 2382 342128 2388
rect 342168 2440 342220 2446
rect 342168 2382 342220 2388
rect 341984 2372 342036 2378
rect 341984 2314 342036 2320
rect 342364 2310 342392 5782
rect 350540 4820 350592 4826
rect 350540 4762 350592 4768
rect 349804 4480 349856 4486
rect 349804 4422 349856 4428
rect 348240 3528 348292 3534
rect 348240 3470 348292 3476
rect 344284 3460 344336 3466
rect 344284 3402 344336 3408
rect 344296 3194 344324 3402
rect 348252 3194 348280 3470
rect 344284 3188 344336 3194
rect 344284 3130 344336 3136
rect 348240 3188 348292 3194
rect 348240 3130 348292 3136
rect 349816 2922 349844 4422
rect 350552 3738 350580 4762
rect 350724 4752 350776 4758
rect 350724 4694 350776 4700
rect 350540 3732 350592 3738
rect 350540 3674 350592 3680
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 349804 2916 349856 2922
rect 349804 2858 349856 2864
rect 345572 2848 345624 2854
rect 345572 2790 345624 2796
rect 346676 2848 346728 2854
rect 346676 2790 346728 2796
rect 348424 2848 348476 2854
rect 348424 2790 348476 2796
rect 349712 2848 349764 2854
rect 349712 2790 349764 2796
rect 345584 2446 345612 2790
rect 345572 2440 345624 2446
rect 345572 2382 345624 2388
rect 346216 2440 346268 2446
rect 346216 2382 346268 2388
rect 346584 2440 346636 2446
rect 346584 2382 346636 2388
rect 342352 2304 342404 2310
rect 342352 2246 342404 2252
rect 345664 2304 345716 2310
rect 345664 2246 345716 2252
rect 345676 1698 345704 2246
rect 345664 1692 345716 1698
rect 345664 1634 345716 1640
rect 346228 1358 346256 2382
rect 346308 1896 346360 1902
rect 346308 1838 346360 1844
rect 346216 1352 346268 1358
rect 346216 1294 346268 1300
rect 341524 1080 341576 1086
rect 341524 1022 341576 1028
rect 346320 746 346348 1838
rect 346308 740 346360 746
rect 346308 682 346360 688
rect 346596 474 346624 2382
rect 346688 2378 346716 2790
rect 348436 2378 348464 2790
rect 349724 2378 349752 2790
rect 350460 2650 350488 3334
rect 350736 3194 350764 4694
rect 351932 3670 351960 6258
rect 357268 6254 357296 9182
rect 362500 7744 362552 7750
rect 362500 7686 362552 7692
rect 357256 6248 357308 6254
rect 357256 6190 357308 6196
rect 362224 6180 362276 6186
rect 362224 6122 362276 6128
rect 355784 6112 355836 6118
rect 355784 6054 355836 6060
rect 355140 5908 355192 5914
rect 355140 5850 355192 5856
rect 353300 4752 353352 4758
rect 353300 4694 353352 4700
rect 351920 3664 351972 3670
rect 351920 3606 351972 3612
rect 350724 3188 350776 3194
rect 350724 3130 350776 3136
rect 353312 3058 353340 4694
rect 353944 3732 353996 3738
rect 353944 3674 353996 3680
rect 353956 3194 353984 3674
rect 354036 3664 354088 3670
rect 354036 3606 354088 3612
rect 353944 3188 353996 3194
rect 353944 3130 353996 3136
rect 353300 3052 353352 3058
rect 353300 2994 353352 3000
rect 354048 2990 354076 3606
rect 354036 2984 354088 2990
rect 354036 2926 354088 2932
rect 350632 2848 350684 2854
rect 350632 2790 350684 2796
rect 352380 2848 352432 2854
rect 352380 2790 352432 2796
rect 353668 2848 353720 2854
rect 353668 2790 353720 2796
rect 354496 2848 354548 2854
rect 354496 2790 354548 2796
rect 350448 2644 350500 2650
rect 350448 2586 350500 2592
rect 350644 2446 350672 2790
rect 350632 2440 350684 2446
rect 350632 2382 350684 2388
rect 346676 2372 346728 2378
rect 346676 2314 346728 2320
rect 348424 2372 348476 2378
rect 348424 2314 348476 2320
rect 349712 2372 349764 2378
rect 349712 2314 349764 2320
rect 346688 1834 346716 2314
rect 346768 2304 346820 2310
rect 346768 2246 346820 2252
rect 346676 1828 346728 1834
rect 346676 1770 346728 1776
rect 346584 468 346636 474
rect 346584 410 346636 416
rect 339960 332 340012 338
rect 339960 274 340012 280
rect 346780 202 346808 2246
rect 348436 270 348464 2314
rect 349620 2304 349672 2310
rect 349620 2246 349672 2252
rect 349632 2106 349660 2246
rect 349620 2100 349672 2106
rect 349620 2042 349672 2048
rect 349724 338 349752 2314
rect 350540 2032 350592 2038
rect 350540 1974 350592 1980
rect 349804 1964 349856 1970
rect 349804 1906 349856 1912
rect 349816 406 349844 1906
rect 350552 678 350580 1974
rect 350644 1902 350672 2382
rect 352392 2378 352420 2790
rect 353680 2446 353708 2790
rect 353668 2440 353720 2446
rect 353668 2382 353720 2388
rect 352380 2372 352432 2378
rect 352380 2314 352432 2320
rect 353300 2372 353352 2378
rect 353300 2314 353352 2320
rect 352288 2304 352340 2310
rect 352288 2246 352340 2252
rect 350632 1896 350684 1902
rect 350632 1838 350684 1844
rect 352300 1630 352328 2246
rect 352288 1624 352340 1630
rect 352288 1566 352340 1572
rect 350540 672 350592 678
rect 350540 614 350592 620
rect 352392 406 352420 2314
rect 353312 2009 353340 2314
rect 354404 2304 354456 2310
rect 354404 2246 354456 2252
rect 353298 2000 353354 2009
rect 353298 1935 353354 1944
rect 354416 1562 354444 2246
rect 354508 1698 354536 2790
rect 355152 2650 355180 5850
rect 355796 2650 355824 6054
rect 355876 5092 355928 5098
rect 355876 5034 355928 5040
rect 355888 3670 355916 5034
rect 357440 5024 357492 5030
rect 357440 4966 357492 4972
rect 355876 3664 355928 3670
rect 355876 3606 355928 3612
rect 357452 3482 357480 4966
rect 356992 3466 357480 3482
rect 356980 3460 357480 3466
rect 357032 3454 357480 3460
rect 356980 3402 357032 3408
rect 357164 3392 357216 3398
rect 357164 3334 357216 3340
rect 357176 3058 357204 3334
rect 362236 3126 362264 6122
rect 362224 3120 362276 3126
rect 362224 3062 362276 3068
rect 357164 3052 357216 3058
rect 357164 2994 357216 3000
rect 359556 2916 359608 2922
rect 359556 2858 359608 2864
rect 356060 2848 356112 2854
rect 356060 2790 356112 2796
rect 358176 2848 358228 2854
rect 358176 2790 358228 2796
rect 355140 2644 355192 2650
rect 355140 2586 355192 2592
rect 355784 2644 355836 2650
rect 355784 2586 355836 2592
rect 355152 2378 355180 2586
rect 356072 2446 356100 2790
rect 358188 2446 358216 2790
rect 359568 2650 359596 2858
rect 359556 2644 359608 2650
rect 359556 2586 359608 2592
rect 359568 2446 359596 2586
rect 362236 2446 362264 3062
rect 362512 2650 362540 7686
rect 375300 6186 375328 9182
rect 391848 8968 391900 8974
rect 391848 8910 391900 8916
rect 408408 8968 408460 8974
rect 408408 8910 408460 8916
rect 387156 8424 387208 8430
rect 387156 8366 387208 8372
rect 385316 7200 385368 7206
rect 385316 7142 385368 7148
rect 380532 6248 380584 6254
rect 380532 6190 380584 6196
rect 375288 6180 375340 6186
rect 375288 6122 375340 6128
rect 367284 4208 367336 4214
rect 367284 4150 367336 4156
rect 362500 2644 362552 2650
rect 362500 2586 362552 2592
rect 367296 2514 367324 4150
rect 380544 2650 380572 6190
rect 381268 4548 381320 4554
rect 381268 4490 381320 4496
rect 380900 2848 380952 2854
rect 380900 2790 380952 2796
rect 380532 2644 380584 2650
rect 380532 2586 380584 2592
rect 367284 2508 367336 2514
rect 367284 2450 367336 2456
rect 380912 2446 380940 2790
rect 381280 2446 381308 4490
rect 382740 3188 382792 3194
rect 382740 3130 382792 3136
rect 382752 2650 382780 3130
rect 382740 2644 382792 2650
rect 382740 2586 382792 2592
rect 382752 2446 382780 2586
rect 385328 2514 385356 7142
rect 387168 2650 387196 8366
rect 391860 6254 391888 8910
rect 395620 8492 395672 8498
rect 395620 8434 395672 8440
rect 391848 6248 391900 6254
rect 391848 6190 391900 6196
rect 390192 5636 390244 5642
rect 390192 5578 390244 5584
rect 388444 4208 388496 4214
rect 388444 4150 388496 4156
rect 387156 2644 387208 2650
rect 387156 2586 387208 2592
rect 385316 2508 385368 2514
rect 385316 2450 385368 2456
rect 387168 2446 387196 2586
rect 388456 2446 388484 4150
rect 390204 3058 390232 5578
rect 393596 3392 393648 3398
rect 393596 3334 393648 3340
rect 394240 3392 394292 3398
rect 394240 3334 394292 3340
rect 394700 3392 394752 3398
rect 394700 3334 394752 3340
rect 390192 3052 390244 3058
rect 390192 2994 390244 3000
rect 390560 3052 390612 3058
rect 390560 2994 390612 3000
rect 390572 2854 390600 2994
rect 393608 2990 393636 3334
rect 394252 3058 394280 3334
rect 394240 3052 394292 3058
rect 394240 2994 394292 3000
rect 394424 3052 394476 3058
rect 394424 2994 394476 3000
rect 391112 2984 391164 2990
rect 391112 2926 391164 2932
rect 393596 2984 393648 2990
rect 393596 2926 393648 2932
rect 390560 2848 390612 2854
rect 390560 2790 390612 2796
rect 391124 2553 391152 2926
rect 391110 2544 391166 2553
rect 391110 2479 391166 2488
rect 391124 2446 391152 2479
rect 356060 2440 356112 2446
rect 356060 2382 356112 2388
rect 358176 2440 358228 2446
rect 358176 2382 358228 2388
rect 359556 2440 359608 2446
rect 359556 2382 359608 2388
rect 362224 2440 362276 2446
rect 380900 2440 380952 2446
rect 362224 2382 362276 2388
rect 372434 2408 372490 2417
rect 355140 2372 355192 2378
rect 355140 2314 355192 2320
rect 355966 2136 356022 2145
rect 355966 2071 356022 2080
rect 354496 1692 354548 1698
rect 354496 1634 354548 1640
rect 354404 1556 354456 1562
rect 354404 1498 354456 1504
rect 355980 1358 356008 2071
rect 355968 1352 356020 1358
rect 355968 1294 356020 1300
rect 356072 474 356100 2382
rect 357900 2372 357952 2378
rect 357900 2314 357952 2320
rect 357912 814 357940 2314
rect 358188 1358 358216 2382
rect 371148 2372 371200 2378
rect 380900 2382 380952 2388
rect 381268 2440 381320 2446
rect 381268 2382 381320 2388
rect 382740 2440 382792 2446
rect 382740 2382 382792 2388
rect 387156 2440 387208 2446
rect 387156 2382 387208 2388
rect 388444 2440 388496 2446
rect 388444 2382 388496 2388
rect 391112 2440 391164 2446
rect 391112 2382 391164 2388
rect 372434 2343 372436 2352
rect 371148 2314 371200 2320
rect 372488 2343 372490 2352
rect 372436 2314 372488 2320
rect 371160 1970 371188 2314
rect 371148 1964 371200 1970
rect 371148 1906 371200 1912
rect 380912 1630 380940 2382
rect 389272 2372 389324 2378
rect 389272 2314 389324 2320
rect 391664 2372 391716 2378
rect 391664 2314 391716 2320
rect 393872 2372 393924 2378
rect 393872 2314 393924 2320
rect 386512 2304 386564 2310
rect 386512 2246 386564 2252
rect 386524 2106 386552 2246
rect 386512 2100 386564 2106
rect 386512 2042 386564 2048
rect 389180 1896 389232 1902
rect 389180 1838 389232 1844
rect 380900 1624 380952 1630
rect 380900 1566 380952 1572
rect 358176 1352 358228 1358
rect 358176 1294 358228 1300
rect 389192 1290 389220 1838
rect 389284 1766 389312 2314
rect 390468 2304 390520 2310
rect 390468 2246 390520 2252
rect 390480 1970 390508 2246
rect 390558 2000 390614 2009
rect 390468 1964 390520 1970
rect 390558 1935 390614 1944
rect 390468 1906 390520 1912
rect 389272 1760 389324 1766
rect 389272 1702 389324 1708
rect 389180 1284 389232 1290
rect 389180 1226 389232 1232
rect 390572 1086 390600 1935
rect 390560 1080 390612 1086
rect 390560 1022 390612 1028
rect 391676 950 391704 2314
rect 393884 1018 393912 2314
rect 394436 2281 394464 2994
rect 394712 2446 394740 3334
rect 395632 2650 395660 8434
rect 403992 8356 404044 8362
rect 403992 8298 404044 8304
rect 403716 7472 403768 7478
rect 403716 7414 403768 7420
rect 403072 7336 403124 7342
rect 403072 7278 403124 7284
rect 396724 7268 396776 7274
rect 396724 7210 396776 7216
rect 396736 3058 396764 7210
rect 402060 6928 402112 6934
rect 402060 6870 402112 6876
rect 398564 6180 398616 6186
rect 398564 6122 398616 6128
rect 396908 3392 396960 3398
rect 396908 3334 396960 3340
rect 397368 3392 397420 3398
rect 397368 3334 397420 3340
rect 396080 3052 396132 3058
rect 396080 2994 396132 3000
rect 396724 3052 396776 3058
rect 396724 2994 396776 3000
rect 395988 2848 396040 2854
rect 395988 2790 396040 2796
rect 395620 2644 395672 2650
rect 395620 2586 395672 2592
rect 394700 2440 394752 2446
rect 394700 2382 394752 2388
rect 394422 2272 394478 2281
rect 394422 2207 394478 2216
rect 394712 1290 394740 2382
rect 394700 1284 394752 1290
rect 394700 1226 394752 1232
rect 393872 1012 393924 1018
rect 393872 954 393924 960
rect 391664 944 391716 950
rect 391664 886 391716 892
rect 357900 808 357952 814
rect 357900 750 357952 756
rect 396000 678 396028 2790
rect 396092 2553 396120 2994
rect 396172 2848 396224 2854
rect 396172 2790 396224 2796
rect 396078 2544 396134 2553
rect 396078 2479 396134 2488
rect 396184 2378 396212 2790
rect 396920 2446 396948 3334
rect 397380 2446 397408 3334
rect 398576 2650 398604 6122
rect 401508 4004 401560 4010
rect 401508 3946 401560 3952
rect 401232 3664 401284 3670
rect 401232 3606 401284 3612
rect 399392 3528 399444 3534
rect 399392 3470 399444 3476
rect 398932 2848 398984 2854
rect 398932 2790 398984 2796
rect 398564 2644 398616 2650
rect 398564 2586 398616 2592
rect 398944 2446 398972 2790
rect 399404 2774 399432 3470
rect 399852 2848 399904 2854
rect 399852 2790 399904 2796
rect 401140 2848 401192 2854
rect 401140 2790 401192 2796
rect 399404 2746 399524 2774
rect 396908 2440 396960 2446
rect 396908 2382 396960 2388
rect 397368 2440 397420 2446
rect 397368 2382 397420 2388
rect 398932 2440 398984 2446
rect 398932 2382 398984 2388
rect 396172 2372 396224 2378
rect 396172 2314 396224 2320
rect 396920 1873 396948 2382
rect 399300 2372 399352 2378
rect 399300 2314 399352 2320
rect 397828 1964 397880 1970
rect 397828 1906 397880 1912
rect 396906 1864 396962 1873
rect 396906 1799 396962 1808
rect 397840 814 397868 1906
rect 399312 1902 399340 2314
rect 399496 1902 399524 2746
rect 399864 2446 399892 2790
rect 400770 2544 400826 2553
rect 400770 2479 400826 2488
rect 399852 2440 399904 2446
rect 399852 2382 399904 2388
rect 399300 1896 399352 1902
rect 399300 1838 399352 1844
rect 399484 1896 399536 1902
rect 399484 1838 399536 1844
rect 399864 1766 399892 2382
rect 399852 1760 399904 1766
rect 399482 1728 399538 1737
rect 399852 1702 399904 1708
rect 399482 1663 399538 1672
rect 399298 1592 399354 1601
rect 399298 1527 399354 1536
rect 398010 1456 398066 1465
rect 398010 1391 398066 1400
rect 399022 1456 399078 1465
rect 399022 1391 399078 1400
rect 398024 1290 398052 1391
rect 398838 1320 398894 1329
rect 398012 1284 398064 1290
rect 398012 1226 398064 1232
rect 398104 1284 398156 1290
rect 399036 1290 399064 1391
rect 398838 1255 398894 1264
rect 399024 1284 399076 1290
rect 398104 1226 398156 1232
rect 397920 1080 397972 1086
rect 397920 1022 397972 1028
rect 397828 808 397880 814
rect 397828 750 397880 756
rect 395988 672 396040 678
rect 395988 614 396040 620
rect 397932 610 397960 1022
rect 398012 944 398064 950
rect 398012 886 398064 892
rect 397920 604 397972 610
rect 397920 546 397972 552
rect 398024 474 398052 886
rect 356060 468 356112 474
rect 356060 410 356112 416
rect 398012 468 398064 474
rect 398012 410 398064 416
rect 349804 400 349856 406
rect 349804 342 349856 348
rect 352380 400 352432 406
rect 352380 342 352432 348
rect 398116 338 398144 1226
rect 398852 1222 398880 1255
rect 399024 1226 399076 1232
rect 398840 1216 398892 1222
rect 398840 1158 398892 1164
rect 398196 876 398248 882
rect 398196 818 398248 824
rect 398208 406 398236 818
rect 399312 746 399340 1527
rect 399300 740 399352 746
rect 399300 682 399352 688
rect 398196 400 398248 406
rect 398196 342 398248 348
rect 349712 332 349764 338
rect 349712 274 349764 280
rect 398104 332 398156 338
rect 398104 274 398156 280
rect 348424 264 348476 270
rect 348424 206 348476 212
rect 399496 202 399524 1663
rect 399576 1556 399628 1562
rect 399576 1498 399628 1504
rect 399588 1086 399616 1498
rect 399666 1320 399722 1329
rect 399666 1255 399722 1264
rect 399680 1154 399708 1255
rect 399850 1184 399906 1193
rect 399668 1148 399720 1154
rect 399850 1119 399906 1128
rect 399668 1090 399720 1096
rect 399576 1080 399628 1086
rect 399576 1022 399628 1028
rect 399760 1080 399812 1086
rect 399760 1022 399812 1028
rect 346768 196 346820 202
rect 346768 138 346820 144
rect 399484 196 399536 202
rect 399484 138 399536 144
rect 399772 134 399800 1022
rect 399864 270 399892 1119
rect 400784 814 400812 2479
rect 401152 2446 401180 2790
rect 401244 2774 401272 3606
rect 401520 2774 401548 3946
rect 401784 3052 401836 3058
rect 401784 2994 401836 3000
rect 401244 2746 401456 2774
rect 401520 2746 401640 2774
rect 401140 2440 401192 2446
rect 401140 2382 401192 2388
rect 400864 2304 400916 2310
rect 400864 2246 400916 2252
rect 400772 808 400824 814
rect 400876 796 400904 2246
rect 401152 1494 401180 2382
rect 401140 1488 401192 1494
rect 401140 1430 401192 1436
rect 400956 1420 401008 1426
rect 400956 1362 401008 1368
rect 400968 1086 400996 1362
rect 401048 1216 401100 1222
rect 401048 1158 401100 1164
rect 401140 1216 401192 1222
rect 401140 1158 401192 1164
rect 400956 1080 401008 1086
rect 400956 1022 401008 1028
rect 401060 898 401088 1158
rect 401152 1018 401180 1158
rect 401140 1012 401192 1018
rect 401140 954 401192 960
rect 401324 944 401376 950
rect 401060 892 401324 898
rect 401060 886 401376 892
rect 401060 870 401364 886
rect 400956 808 401008 814
rect 400876 768 400956 796
rect 400772 750 400824 756
rect 400956 750 401008 756
rect 401324 808 401376 814
rect 401428 796 401456 2746
rect 401508 2372 401560 2378
rect 401508 2314 401560 2320
rect 401520 1562 401548 2314
rect 401508 1556 401560 1562
rect 401508 1498 401560 1504
rect 401612 882 401640 2746
rect 401600 876 401652 882
rect 401600 818 401652 824
rect 401796 814 401824 2994
rect 402072 814 402100 6870
rect 402336 5024 402388 5030
rect 402336 4966 402388 4972
rect 402348 814 402376 4966
rect 402610 1592 402666 1601
rect 402610 1527 402666 1536
rect 402624 814 402652 1527
rect 402704 1420 402756 1426
rect 402704 1362 402756 1368
rect 402716 1154 402744 1362
rect 402704 1148 402756 1154
rect 402704 1090 402756 1096
rect 401376 768 401456 796
rect 401784 808 401836 814
rect 401324 750 401376 756
rect 401784 750 401836 756
rect 402060 808 402112 814
rect 402060 750 402112 756
rect 402336 808 402388 814
rect 402336 750 402388 756
rect 402612 808 402664 814
rect 403084 796 403112 7278
rect 403728 814 403756 7414
rect 403808 4820 403860 4826
rect 403808 4762 403860 4768
rect 403164 808 403216 814
rect 403084 768 403164 796
rect 402612 750 402664 756
rect 403164 750 403216 756
rect 403716 808 403768 814
rect 403716 750 403768 756
rect 399944 672 399996 678
rect 400220 672 400272 678
rect 399996 632 400220 660
rect 399944 614 399996 620
rect 400220 614 400272 620
rect 403440 672 403492 678
rect 403820 626 403848 4762
rect 403900 4276 403952 4282
rect 403900 4218 403952 4224
rect 403912 796 403940 4218
rect 404004 2514 404032 8298
rect 408316 7744 408368 7750
rect 408316 7686 408368 7692
rect 404544 7540 404596 7546
rect 404544 7482 404596 7488
rect 403992 2508 404044 2514
rect 403992 2450 404044 2456
rect 404266 1320 404322 1329
rect 404266 1255 404322 1264
rect 404280 814 404308 1255
rect 404556 814 404584 7482
rect 407212 7404 407264 7410
rect 407212 7346 407264 7352
rect 407120 5772 407172 5778
rect 407120 5714 407172 5720
rect 406108 5704 406160 5710
rect 406108 5646 406160 5652
rect 405280 4684 405332 4690
rect 405280 4626 405332 4632
rect 405188 2372 405240 2378
rect 405188 2314 405240 2320
rect 405096 1488 405148 1494
rect 404818 1456 404874 1465
rect 405096 1430 405148 1436
rect 404818 1391 404874 1400
rect 404832 814 404860 1391
rect 405108 814 405136 1430
rect 405200 1426 405228 2314
rect 405188 1420 405240 1426
rect 405188 1362 405240 1368
rect 403992 808 404044 814
rect 403912 768 403992 796
rect 403992 750 404044 756
rect 404268 808 404320 814
rect 404268 750 404320 756
rect 404544 808 404596 814
rect 404544 750 404596 756
rect 404820 808 404872 814
rect 404820 750 404872 756
rect 405096 808 405148 814
rect 405292 796 405320 4626
rect 405924 4616 405976 4622
rect 405924 4558 405976 4564
rect 405936 814 405964 4558
rect 405372 808 405424 814
rect 405292 768 405372 796
rect 405096 750 405148 756
rect 405372 750 405424 756
rect 405924 808 405976 814
rect 406120 796 406148 5646
rect 406200 4480 406252 4486
rect 406200 4422 406252 4428
rect 406212 2774 406240 4422
rect 406476 3596 406528 3602
rect 406476 3538 406528 3544
rect 406212 2746 406332 2774
rect 406200 808 406252 814
rect 406120 768 406200 796
rect 405924 750 405976 756
rect 406200 750 406252 756
rect 403492 620 403848 626
rect 403440 614 403848 620
rect 403452 598 403848 614
rect 403440 536 403492 542
rect 400494 504 400550 513
rect 400678 504 400734 513
rect 400494 439 400496 448
rect 400548 439 400550 448
rect 400600 462 400678 490
rect 400496 410 400548 416
rect 400600 354 400628 462
rect 400678 439 400734 448
rect 403438 504 403440 513
rect 406200 536 406252 542
rect 403492 504 403494 513
rect 406304 490 406332 2746
rect 406384 944 406436 950
rect 406384 886 406436 892
rect 406396 513 406424 886
rect 406488 814 406516 3538
rect 406936 1488 406988 1494
rect 406936 1430 406988 1436
rect 406752 1148 406804 1154
rect 406752 1090 406804 1096
rect 406764 814 406792 1090
rect 406948 1086 406976 1430
rect 406936 1080 406988 1086
rect 406936 1022 406988 1028
rect 406476 808 406528 814
rect 406476 750 406528 756
rect 406752 808 406804 814
rect 407132 796 407160 5714
rect 407224 2514 407252 7346
rect 407764 5840 407816 5846
rect 407764 5782 407816 5788
rect 407304 4752 407356 4758
rect 407304 4694 407356 4700
rect 407212 2508 407264 2514
rect 407212 2450 407264 2456
rect 407212 1420 407264 1426
rect 407212 1362 407264 1368
rect 407224 1018 407252 1362
rect 407212 1012 407264 1018
rect 407212 954 407264 960
rect 407316 814 407344 4694
rect 407672 2304 407724 2310
rect 407672 2246 407724 2252
rect 407684 1562 407712 2246
rect 407580 1556 407632 1562
rect 407580 1498 407632 1504
rect 407672 1556 407724 1562
rect 407672 1498 407724 1504
rect 407488 1352 407540 1358
rect 407486 1320 407488 1329
rect 407540 1320 407542 1329
rect 407486 1255 407542 1264
rect 407486 1184 407542 1193
rect 407486 1119 407488 1128
rect 407540 1119 407542 1128
rect 407488 1090 407540 1096
rect 407592 1018 407620 1498
rect 407580 1012 407632 1018
rect 407580 954 407632 960
rect 407776 814 407804 5782
rect 407856 2644 407908 2650
rect 407856 2586 407908 2592
rect 407212 808 407264 814
rect 407132 768 407212 796
rect 406752 750 406804 756
rect 407212 750 407264 756
rect 407304 808 407356 814
rect 407304 750 407356 756
rect 407764 808 407816 814
rect 407764 750 407816 756
rect 407764 672 407816 678
rect 407868 626 407896 2586
rect 408328 2446 408356 7686
rect 408420 6186 408448 8910
rect 411812 6996 411864 7002
rect 411812 6938 411864 6944
rect 408408 6180 408460 6186
rect 408408 6122 408460 6128
rect 409972 5908 410024 5914
rect 409972 5850 410024 5856
rect 409420 3460 409472 3466
rect 409420 3402 409472 3408
rect 408500 2848 408552 2854
rect 408500 2790 408552 2796
rect 408512 2650 408540 2790
rect 408500 2644 408552 2650
rect 408500 2586 408552 2592
rect 408512 2514 408540 2586
rect 408500 2508 408552 2514
rect 408500 2450 408552 2456
rect 408316 2440 408368 2446
rect 408316 2382 408368 2388
rect 408040 1896 408092 1902
rect 408040 1838 408092 1844
rect 408052 814 408080 1838
rect 408316 1828 408368 1834
rect 408316 1770 408368 1776
rect 408328 814 408356 1770
rect 408408 1760 408460 1766
rect 408408 1702 408460 1708
rect 408590 1728 408646 1737
rect 408420 1358 408448 1702
rect 408590 1663 408646 1672
rect 408408 1352 408460 1358
rect 408408 1294 408460 1300
rect 408604 814 408632 1663
rect 408868 1148 408920 1154
rect 408868 1090 408920 1096
rect 408880 814 408908 1090
rect 409432 814 409460 3402
rect 409696 2372 409748 2378
rect 409696 2314 409748 2320
rect 409708 882 409736 2314
rect 409696 876 409748 882
rect 409696 818 409748 824
rect 409984 814 410012 5850
rect 410248 3732 410300 3738
rect 410248 3674 410300 3680
rect 410260 814 410288 3674
rect 411076 3120 411128 3126
rect 411076 3062 411128 3068
rect 410524 1488 410576 1494
rect 410524 1430 410576 1436
rect 410536 814 410564 1430
rect 410798 1320 410854 1329
rect 410798 1255 410854 1264
rect 410812 814 410840 1255
rect 411088 814 411116 3062
rect 411824 2514 411852 6938
rect 426360 6254 426388 9182
rect 416320 6248 416372 6254
rect 416320 6190 416372 6196
rect 426348 6248 426400 6254
rect 426348 6190 426400 6196
rect 442816 6248 442868 6254
rect 442816 6190 442868 6196
rect 416332 3126 416360 6190
rect 434628 6180 434680 6186
rect 434628 6122 434680 6128
rect 421380 5568 421432 5574
rect 421380 5510 421432 5516
rect 416320 3120 416372 3126
rect 416320 3062 416372 3068
rect 411812 2508 411864 2514
rect 411812 2450 411864 2456
rect 416332 2446 416360 3062
rect 421392 2446 421420 5510
rect 422576 3120 422628 3126
rect 422576 3062 422628 3068
rect 422588 2582 422616 3062
rect 434640 2582 434668 6122
rect 442828 4826 442856 6190
rect 442920 6186 442948 9182
rect 462692 9124 463012 9796
rect 462692 9068 462704 9124
rect 462760 9068 462784 9124
rect 462840 9068 462864 9124
rect 462920 9068 462944 9124
rect 463000 9068 463012 9124
rect 462692 9044 463012 9068
rect 462692 8988 462704 9044
rect 462760 8988 462784 9044
rect 462840 8988 462864 9044
rect 462920 8988 462944 9044
rect 463000 8988 463012 9044
rect 462692 8964 463012 8988
rect 462692 8908 462704 8964
rect 462760 8908 462784 8964
rect 462840 8908 462864 8964
rect 462920 8908 462944 8964
rect 463000 8908 463012 8964
rect 462692 8884 463012 8908
rect 462692 8828 462704 8884
rect 462760 8828 462784 8884
rect 462840 8828 462864 8884
rect 462920 8828 462944 8884
rect 463000 8828 463012 8884
rect 462692 7098 463012 8828
rect 462692 7046 462698 7098
rect 462750 7080 462762 7098
rect 462814 7080 462826 7098
rect 462878 7080 462890 7098
rect 462942 7080 462954 7098
rect 462760 7046 462762 7080
rect 462942 7046 462944 7080
rect 463006 7046 463012 7098
rect 462692 7024 462704 7046
rect 462760 7024 462784 7046
rect 462840 7024 462864 7046
rect 462920 7024 462944 7046
rect 463000 7024 463012 7046
rect 462692 7000 463012 7024
rect 462692 6944 462704 7000
rect 462760 6944 462784 7000
rect 462840 6944 462864 7000
rect 462920 6944 462944 7000
rect 463000 6944 463012 7000
rect 462692 6920 463012 6944
rect 462692 6864 462704 6920
rect 462760 6864 462784 6920
rect 462840 6864 462864 6920
rect 462920 6864 462944 6920
rect 463000 6864 463012 6920
rect 462692 6840 463012 6864
rect 462692 6784 462704 6840
rect 462760 6784 462784 6840
rect 462840 6784 462864 6840
rect 462920 6784 462944 6840
rect 463000 6784 463012 6840
rect 442908 6180 442960 6186
rect 442908 6122 442960 6128
rect 462692 6010 463012 6784
rect 462692 5958 462698 6010
rect 462750 5958 462762 6010
rect 462814 5958 462826 6010
rect 462878 5958 462890 6010
rect 462942 5958 462954 6010
rect 463006 5958 463012 6010
rect 462692 5721 463012 5958
rect 462692 5665 462704 5721
rect 462760 5665 462784 5721
rect 462840 5665 462864 5721
rect 462920 5665 462944 5721
rect 463000 5665 463012 5721
rect 462692 5641 463012 5665
rect 462692 5585 462704 5641
rect 462760 5585 462784 5641
rect 462840 5585 462864 5641
rect 462920 5585 462944 5641
rect 463000 5585 463012 5641
rect 462692 5561 463012 5585
rect 462692 5505 462704 5561
rect 462760 5505 462784 5561
rect 462840 5505 462864 5561
rect 462920 5505 462944 5561
rect 463000 5505 463012 5561
rect 462692 5481 463012 5505
rect 462692 5425 462704 5481
rect 462760 5425 462784 5481
rect 462840 5425 462864 5481
rect 462920 5425 462944 5481
rect 463000 5425 463012 5481
rect 462692 4922 463012 5425
rect 462692 4870 462698 4922
rect 462750 4870 462762 4922
rect 462814 4870 462826 4922
rect 462878 4870 462890 4922
rect 462942 4870 462954 4922
rect 463006 4870 463012 4922
rect 442816 4820 442868 4826
rect 442816 4762 442868 4768
rect 452660 4820 452712 4826
rect 452660 4762 452712 4768
rect 434996 2848 435048 2854
rect 434996 2790 435048 2796
rect 435732 2848 435784 2854
rect 435732 2790 435784 2796
rect 435008 2582 435036 2790
rect 422576 2576 422628 2582
rect 422576 2518 422628 2524
rect 434628 2576 434680 2582
rect 434628 2518 434680 2524
rect 434996 2576 435048 2582
rect 434996 2518 435048 2524
rect 422588 2446 422616 2518
rect 435008 2446 435036 2518
rect 435744 2446 435772 2790
rect 416320 2440 416372 2446
rect 416320 2382 416372 2388
rect 421380 2440 421432 2446
rect 421380 2382 421432 2388
rect 422576 2440 422628 2446
rect 422576 2382 422628 2388
rect 434996 2440 435048 2446
rect 434996 2382 435048 2388
rect 435732 2440 435784 2446
rect 435732 2382 435784 2388
rect 425152 2372 425204 2378
rect 425152 2314 425204 2320
rect 435456 2372 435508 2378
rect 435456 2314 435508 2320
rect 413008 2304 413060 2310
rect 413008 2246 413060 2252
rect 416596 2304 416648 2310
rect 416596 2246 416648 2252
rect 413020 1222 413048 2246
rect 413008 1216 413060 1222
rect 413008 1158 413060 1164
rect 416608 1154 416636 2246
rect 425164 2038 425192 2314
rect 426532 2304 426584 2310
rect 426532 2246 426584 2252
rect 426544 2038 426572 2246
rect 425152 2032 425204 2038
rect 425152 1974 425204 1980
rect 426532 2032 426584 2038
rect 435468 2009 435496 2314
rect 426532 1974 426584 1980
rect 435454 2000 435510 2009
rect 435454 1935 435510 1944
rect 435744 1358 435772 2382
rect 439412 2372 439464 2378
rect 439412 2314 439464 2320
rect 447784 2372 447836 2378
rect 447784 2314 447836 2320
rect 439424 2145 439452 2314
rect 440608 2304 440660 2310
rect 440608 2246 440660 2252
rect 439410 2136 439466 2145
rect 439410 2071 439466 2080
rect 440620 1970 440648 2246
rect 440608 1964 440660 1970
rect 440608 1906 440660 1912
rect 447796 1698 447824 2314
rect 452672 2310 452700 4762
rect 462692 4362 463012 4870
rect 462692 4306 462704 4362
rect 462760 4306 462784 4362
rect 462840 4306 462864 4362
rect 462920 4306 462944 4362
rect 463000 4306 463012 4362
rect 462692 4282 463012 4306
rect 462692 4226 462704 4282
rect 462760 4226 462784 4282
rect 462840 4226 462864 4282
rect 462920 4226 462944 4282
rect 463000 4226 463012 4282
rect 462692 4202 463012 4226
rect 462692 4146 462704 4202
rect 462760 4146 462784 4202
rect 462840 4146 462864 4202
rect 462920 4146 462944 4202
rect 463000 4146 463012 4202
rect 462692 4122 463012 4146
rect 462692 4066 462704 4122
rect 462760 4066 462784 4122
rect 462840 4066 462864 4122
rect 462920 4066 462944 4122
rect 463000 4066 463012 4122
rect 462692 3834 463012 4066
rect 462692 3782 462698 3834
rect 462750 3782 462762 3834
rect 462814 3782 462826 3834
rect 462878 3782 462890 3834
rect 462942 3782 462954 3834
rect 463006 3782 463012 3834
rect 462692 3003 463012 3782
rect 462692 2947 462704 3003
rect 462760 2947 462784 3003
rect 462840 2947 462864 3003
rect 462920 2947 462944 3003
rect 463000 2947 463012 3003
rect 462692 2923 463012 2947
rect 462692 2867 462704 2923
rect 462760 2867 462784 2923
rect 462840 2867 462864 2923
rect 462920 2867 462944 2923
rect 463000 2867 463012 2923
rect 462692 2843 463012 2867
rect 462692 2787 462704 2843
rect 462760 2787 462784 2843
rect 462840 2787 462864 2843
rect 462920 2787 462944 2843
rect 463000 2787 463012 2843
rect 462692 2763 463012 2787
rect 462692 2746 462704 2763
rect 462760 2746 462784 2763
rect 462840 2746 462864 2763
rect 462920 2746 462944 2763
rect 463000 2746 463012 2763
rect 462692 2694 462698 2746
rect 462760 2707 462762 2746
rect 462942 2707 462944 2746
rect 462750 2694 462762 2707
rect 462814 2694 462826 2707
rect 462878 2694 462890 2707
rect 462942 2694 462954 2707
rect 463006 2694 463012 2746
rect 448612 2304 448664 2310
rect 448612 2246 448664 2252
rect 452660 2304 452712 2310
rect 452660 2246 452712 2252
rect 453396 2304 453448 2310
rect 453396 2246 453448 2252
rect 461860 2304 461912 2310
rect 461860 2246 461912 2252
rect 448624 1902 448652 2246
rect 448612 1896 448664 1902
rect 448612 1838 448664 1844
rect 453408 1834 453436 2246
rect 453396 1828 453448 1834
rect 453396 1770 453448 1776
rect 447784 1692 447836 1698
rect 447784 1634 447836 1640
rect 461872 1562 461900 2246
rect 461860 1556 461912 1562
rect 461860 1498 461912 1504
rect 435732 1352 435784 1358
rect 435732 1294 435784 1300
rect 416596 1148 416648 1154
rect 416596 1090 416648 1096
rect 411444 1080 411496 1086
rect 411444 1022 411496 1028
rect 411456 882 411484 1022
rect 462692 964 463012 2694
rect 462692 908 462704 964
rect 462760 908 462784 964
rect 462840 908 462864 964
rect 462920 908 462944 964
rect 463000 908 463012 964
rect 462692 884 463012 908
rect 411444 876 411496 882
rect 411444 818 411496 824
rect 462692 828 462704 884
rect 462760 828 462784 884
rect 462840 828 462864 884
rect 462920 828 462944 884
rect 463000 828 463012 884
rect 408040 808 408092 814
rect 408040 750 408092 756
rect 408316 808 408368 814
rect 408316 750 408368 756
rect 408592 808 408644 814
rect 408592 750 408644 756
rect 408868 808 408920 814
rect 408868 750 408920 756
rect 409420 808 409472 814
rect 409420 750 409472 756
rect 409972 808 410024 814
rect 409972 750 410024 756
rect 410248 808 410300 814
rect 410248 750 410300 756
rect 410524 808 410576 814
rect 410524 750 410576 756
rect 410800 808 410852 814
rect 410800 750 410852 756
rect 411076 808 411128 814
rect 411076 750 411128 756
rect 462692 804 463012 828
rect 407816 620 407896 626
rect 407764 614 407896 620
rect 407776 598 407896 614
rect 462692 748 462704 804
rect 462760 748 462784 804
rect 462840 748 462864 804
rect 462920 748 462944 804
rect 463000 748 463012 804
rect 462692 724 463012 748
rect 462692 668 462704 724
rect 462760 668 462784 724
rect 462840 668 462864 724
rect 462920 668 462944 724
rect 463000 668 463012 724
rect 409696 536 409748 542
rect 406252 484 406332 490
rect 406200 478 406332 484
rect 406212 462 406332 478
rect 406382 504 406438 513
rect 403438 439 403494 448
rect 406382 439 406438 448
rect 409694 504 409696 513
rect 409748 504 409750 513
rect 409694 439 409750 448
rect 399956 326 400628 354
rect 399852 264 399904 270
rect 399852 206 399904 212
rect 331424 64 331744 88
rect 337292 128 337344 134
rect 337292 70 337344 76
rect 399760 128 399812 134
rect 399760 70 399812 76
rect 399956 66 399984 326
rect 331424 8 331436 64
rect 331492 8 331516 64
rect 331572 8 331596 64
rect 331652 8 331676 64
rect 331732 8 331744 64
rect 331424 -4 331744 8
rect 399944 60 399996 66
rect 399944 2 399996 8
rect 462692 -4 463012 668
rect 463352 9784 463672 9796
rect 463352 9728 463364 9784
rect 463420 9728 463444 9784
rect 463500 9728 463524 9784
rect 463580 9728 463604 9784
rect 463660 9728 463672 9784
rect 463352 9704 463672 9728
rect 463352 9648 463364 9704
rect 463420 9648 463444 9704
rect 463500 9648 463524 9704
rect 463580 9648 463604 9704
rect 463660 9648 463672 9704
rect 463352 9624 463672 9648
rect 463352 9568 463364 9624
rect 463420 9568 463444 9624
rect 463500 9568 463524 9624
rect 463580 9568 463604 9624
rect 463660 9568 463672 9624
rect 463352 9544 463672 9568
rect 463352 9488 463364 9544
rect 463420 9488 463444 9544
rect 463500 9488 463524 9544
rect 463580 9488 463604 9544
rect 463660 9488 463672 9544
rect 463352 7740 463672 9488
rect 530676 9784 530996 9796
rect 530676 9728 530688 9784
rect 530744 9728 530768 9784
rect 530824 9728 530848 9784
rect 530904 9728 530928 9784
rect 530984 9728 530996 9784
rect 530676 9704 530996 9728
rect 530676 9648 530688 9704
rect 530744 9648 530768 9704
rect 530824 9648 530848 9704
rect 530904 9648 530928 9704
rect 530984 9648 530996 9704
rect 530676 9624 530996 9648
rect 530676 9568 530688 9624
rect 530744 9568 530768 9624
rect 530824 9568 530848 9624
rect 530904 9568 530928 9624
rect 530984 9568 530996 9624
rect 530676 9544 530996 9568
rect 530676 9488 530688 9544
rect 530744 9488 530768 9544
rect 530824 9488 530848 9544
rect 530904 9488 530928 9544
rect 530984 9488 530996 9544
rect 463352 7684 463364 7740
rect 463420 7684 463444 7740
rect 463500 7684 463524 7740
rect 463580 7684 463604 7740
rect 463660 7684 463672 7740
rect 463352 7660 463672 7684
rect 463352 7642 463364 7660
rect 463420 7642 463444 7660
rect 463500 7642 463524 7660
rect 463580 7642 463604 7660
rect 463660 7642 463672 7660
rect 463352 7590 463358 7642
rect 463420 7604 463422 7642
rect 463602 7604 463604 7642
rect 463410 7590 463422 7604
rect 463474 7590 463486 7604
rect 463538 7590 463550 7604
rect 463602 7590 463614 7604
rect 463666 7590 463672 7642
rect 463352 7580 463672 7590
rect 463352 7524 463364 7580
rect 463420 7524 463444 7580
rect 463500 7524 463524 7580
rect 463580 7524 463604 7580
rect 463660 7524 463672 7580
rect 463352 7500 463672 7524
rect 463352 7444 463364 7500
rect 463420 7444 463444 7500
rect 463500 7444 463524 7500
rect 463580 7444 463604 7500
rect 463660 7444 463672 7500
rect 463352 6554 463672 7444
rect 463352 6502 463358 6554
rect 463410 6502 463422 6554
rect 463474 6502 463486 6554
rect 463538 6502 463550 6554
rect 463602 6502 463614 6554
rect 463666 6502 463672 6554
rect 463352 6381 463672 6502
rect 463352 6325 463364 6381
rect 463420 6325 463444 6381
rect 463500 6325 463524 6381
rect 463580 6325 463604 6381
rect 463660 6325 463672 6381
rect 463352 6301 463672 6325
rect 463352 6245 463364 6301
rect 463420 6245 463444 6301
rect 463500 6245 463524 6301
rect 463580 6245 463604 6301
rect 463660 6245 463672 6301
rect 463352 6221 463672 6245
rect 463352 6165 463364 6221
rect 463420 6165 463444 6221
rect 463500 6165 463524 6221
rect 463580 6165 463604 6221
rect 463660 6165 463672 6221
rect 530016 9124 530336 9136
rect 530016 9068 530028 9124
rect 530084 9068 530108 9124
rect 530164 9068 530188 9124
rect 530244 9068 530268 9124
rect 530324 9068 530336 9124
rect 530016 9044 530336 9068
rect 530016 8988 530028 9044
rect 530084 8988 530108 9044
rect 530164 8988 530188 9044
rect 530244 8988 530268 9044
rect 530324 8988 530336 9044
rect 530016 8964 530336 8988
rect 530016 8908 530028 8964
rect 530084 8908 530108 8964
rect 530164 8908 530188 8964
rect 530244 8908 530268 8964
rect 530324 8908 530336 8964
rect 530016 8884 530336 8908
rect 530016 8828 530028 8884
rect 530084 8828 530108 8884
rect 530164 8828 530188 8884
rect 530244 8828 530268 8884
rect 530324 8828 530336 8884
rect 530016 7080 530336 8828
rect 530016 7024 530028 7080
rect 530084 7024 530108 7080
rect 530164 7024 530188 7080
rect 530244 7024 530268 7080
rect 530324 7024 530336 7080
rect 530016 7000 530336 7024
rect 530016 6944 530028 7000
rect 530084 6944 530108 7000
rect 530164 6944 530188 7000
rect 530244 6944 530268 7000
rect 530324 6944 530336 7000
rect 530016 6920 530336 6944
rect 530016 6864 530028 6920
rect 530084 6864 530108 6920
rect 530164 6864 530188 6920
rect 530244 6864 530268 6920
rect 530324 6864 530336 6920
rect 530016 6840 530336 6864
rect 530016 6784 530028 6840
rect 530084 6784 530108 6840
rect 530164 6784 530188 6840
rect 530244 6784 530268 6840
rect 530324 6784 530336 6840
rect 463352 6141 463672 6165
rect 463352 6085 463364 6141
rect 463420 6085 463444 6141
rect 463500 6085 463524 6141
rect 463580 6085 463604 6141
rect 463660 6085 463672 6141
rect 470416 6180 470468 6186
rect 470416 6122 470468 6128
rect 463352 5466 463672 6085
rect 463352 5414 463358 5466
rect 463410 5414 463422 5466
rect 463474 5414 463486 5466
rect 463538 5414 463550 5466
rect 463602 5414 463614 5466
rect 463666 5414 463672 5466
rect 463352 5022 463672 5414
rect 463352 4966 463364 5022
rect 463420 4966 463444 5022
rect 463500 4966 463524 5022
rect 463580 4966 463604 5022
rect 463660 4966 463672 5022
rect 463352 4942 463672 4966
rect 463352 4886 463364 4942
rect 463420 4886 463444 4942
rect 463500 4886 463524 4942
rect 463580 4886 463604 4942
rect 463660 4886 463672 4942
rect 463352 4862 463672 4886
rect 463352 4806 463364 4862
rect 463420 4806 463444 4862
rect 463500 4806 463524 4862
rect 463580 4806 463604 4862
rect 463660 4806 463672 4862
rect 463352 4782 463672 4806
rect 463352 4726 463364 4782
rect 463420 4726 463444 4782
rect 463500 4726 463524 4782
rect 463580 4726 463604 4782
rect 463660 4726 463672 4782
rect 463352 4378 463672 4726
rect 463352 4326 463358 4378
rect 463410 4326 463422 4378
rect 463474 4326 463486 4378
rect 463538 4326 463550 4378
rect 463602 4326 463614 4378
rect 463666 4326 463672 4378
rect 463352 3663 463672 4326
rect 463352 3607 463364 3663
rect 463420 3607 463444 3663
rect 463500 3607 463524 3663
rect 463580 3607 463604 3663
rect 463660 3607 463672 3663
rect 463352 3583 463672 3607
rect 463352 3527 463364 3583
rect 463420 3527 463444 3583
rect 463500 3527 463524 3583
rect 463580 3527 463604 3583
rect 463660 3527 463672 3583
rect 463352 3503 463672 3527
rect 463352 3447 463364 3503
rect 463420 3447 463444 3503
rect 463500 3447 463524 3503
rect 463580 3447 463604 3503
rect 463660 3447 463672 3503
rect 463352 3423 463672 3447
rect 463352 3367 463364 3423
rect 463420 3367 463444 3423
rect 463500 3367 463524 3423
rect 463580 3367 463604 3423
rect 463660 3367 463672 3423
rect 463352 3290 463672 3367
rect 463352 3238 463358 3290
rect 463410 3238 463422 3290
rect 463474 3238 463486 3290
rect 463538 3238 463550 3290
rect 463602 3238 463614 3290
rect 463666 3238 463672 3290
rect 463352 2202 463672 3238
rect 470428 2922 470456 6122
rect 530016 5721 530336 6784
rect 530016 5665 530028 5721
rect 530084 5665 530108 5721
rect 530164 5665 530188 5721
rect 530244 5665 530268 5721
rect 530324 5665 530336 5721
rect 530016 5641 530336 5665
rect 530016 5585 530028 5641
rect 530084 5585 530108 5641
rect 530164 5585 530188 5641
rect 530244 5585 530268 5641
rect 530324 5585 530336 5641
rect 530016 5561 530336 5585
rect 530016 5505 530028 5561
rect 530084 5505 530108 5561
rect 530164 5505 530188 5561
rect 530244 5505 530268 5561
rect 530324 5505 530336 5561
rect 530016 5481 530336 5505
rect 530016 5425 530028 5481
rect 530084 5425 530108 5481
rect 530164 5425 530188 5481
rect 530244 5425 530268 5481
rect 530324 5425 530336 5481
rect 530016 4362 530336 5425
rect 530016 4306 530028 4362
rect 530084 4306 530108 4362
rect 530164 4306 530188 4362
rect 530244 4306 530268 4362
rect 530324 4306 530336 4362
rect 530016 4282 530336 4306
rect 530016 4226 530028 4282
rect 530084 4226 530108 4282
rect 530164 4226 530188 4282
rect 530244 4226 530268 4282
rect 530324 4226 530336 4282
rect 481640 4208 481692 4214
rect 481640 4150 481692 4156
rect 530016 4202 530336 4226
rect 478880 3188 478932 3194
rect 478880 3130 478932 3136
rect 470416 2916 470468 2922
rect 470416 2858 470468 2864
rect 470428 2446 470456 2858
rect 465724 2440 465776 2446
rect 465722 2408 465724 2417
rect 470416 2440 470468 2446
rect 465776 2408 465778 2417
rect 470416 2382 470468 2388
rect 465722 2343 465778 2352
rect 474372 2372 474424 2378
rect 474372 2314 474424 2320
rect 466552 2304 466604 2310
rect 466552 2246 466604 2252
rect 470692 2304 470744 2310
rect 470692 2246 470744 2252
rect 463352 2150 463358 2202
rect 463410 2150 463422 2202
rect 463474 2150 463486 2202
rect 463538 2150 463550 2202
rect 463602 2150 463614 2202
rect 463666 2150 463672 2202
rect 463352 304 463672 2150
rect 466564 1698 466592 2246
rect 466552 1692 466604 1698
rect 466552 1634 466604 1640
rect 463352 248 463364 304
rect 463420 248 463444 304
rect 463500 248 463524 304
rect 463580 248 463604 304
rect 463660 248 463672 304
rect 463352 224 463672 248
rect 463352 168 463364 224
rect 463420 168 463444 224
rect 463500 168 463524 224
rect 463580 168 463604 224
rect 463660 168 463672 224
rect 463352 144 463672 168
rect 463352 88 463364 144
rect 463420 88 463444 144
rect 463500 88 463524 144
rect 463580 88 463604 144
rect 463660 88 463672 144
rect 463352 64 463672 88
rect 470704 66 470732 2246
rect 474384 1630 474412 2314
rect 475476 2304 475528 2310
rect 475476 2246 475528 2252
rect 475488 1766 475516 2246
rect 475476 1760 475528 1766
rect 475476 1702 475528 1708
rect 474372 1624 474424 1630
rect 474372 1566 474424 1572
rect 478432 1426 478828 1442
rect 478420 1420 478840 1426
rect 478472 1414 478788 1420
rect 478420 1362 478472 1368
rect 478788 1362 478840 1368
rect 478892 814 478920 3130
rect 478972 2372 479024 2378
rect 478972 2314 479024 2320
rect 478984 2106 479012 2314
rect 479800 2304 479852 2310
rect 479800 2246 479852 2252
rect 478972 2100 479024 2106
rect 478972 2042 479024 2048
rect 479812 1630 479840 2246
rect 479800 1624 479852 1630
rect 479800 1566 479852 1572
rect 480996 1488 481048 1494
rect 480996 1430 481048 1436
rect 479616 1352 479668 1358
rect 479616 1294 479668 1300
rect 479628 950 479656 1294
rect 480352 1284 480404 1290
rect 480352 1226 480404 1232
rect 480904 1284 480956 1290
rect 480904 1226 480956 1232
rect 479616 944 479668 950
rect 479616 886 479668 892
rect 479708 944 479760 950
rect 479708 886 479760 892
rect 478880 808 478932 814
rect 478880 750 478932 756
rect 479720 610 479748 886
rect 480364 814 480392 1226
rect 480916 1086 480944 1226
rect 481008 1086 481036 1430
rect 480904 1080 480956 1086
rect 480904 1022 480956 1028
rect 480996 1080 481048 1086
rect 480996 1022 481048 1028
rect 481652 814 481680 4150
rect 530016 4146 530028 4202
rect 530084 4146 530108 4202
rect 530164 4146 530188 4202
rect 530244 4146 530268 4202
rect 530324 4146 530336 4202
rect 530016 4122 530336 4146
rect 530016 4066 530028 4122
rect 530084 4066 530108 4122
rect 530164 4066 530188 4122
rect 530244 4066 530268 4122
rect 530324 4066 530336 4122
rect 491300 3392 491352 3398
rect 491300 3334 491352 3340
rect 484584 3052 484636 3058
rect 484584 2994 484636 3000
rect 482560 1080 482612 1086
rect 482560 1022 482612 1028
rect 482652 1080 482704 1086
rect 482652 1022 482704 1028
rect 482572 814 482600 1022
rect 480352 808 480404 814
rect 480352 750 480404 756
rect 481640 808 481692 814
rect 481640 750 481692 756
rect 482560 808 482612 814
rect 482560 750 482612 756
rect 479708 604 479760 610
rect 479708 546 479760 552
rect 482664 513 482692 1022
rect 484596 814 484624 2994
rect 488632 2984 488684 2990
rect 488632 2926 488684 2932
rect 488540 1964 488592 1970
rect 488540 1906 488592 1912
rect 485872 1896 485924 1902
rect 485872 1838 485924 1844
rect 484768 1828 484820 1834
rect 484768 1770 484820 1776
rect 484780 1358 484808 1770
rect 484676 1352 484728 1358
rect 484676 1294 484728 1300
rect 484768 1352 484820 1358
rect 484768 1294 484820 1300
rect 484688 814 484716 1294
rect 485884 1290 485912 1838
rect 485780 1284 485832 1290
rect 485780 1226 485832 1232
rect 485872 1284 485924 1290
rect 485872 1226 485924 1232
rect 485792 814 485820 1226
rect 488552 1222 488580 1906
rect 486884 1216 486936 1222
rect 486884 1158 486936 1164
rect 488540 1216 488592 1222
rect 488540 1158 488592 1164
rect 486896 814 486924 1158
rect 488644 814 488672 2926
rect 489828 1692 489880 1698
rect 489828 1634 489880 1640
rect 488816 1284 488868 1290
rect 488816 1226 488868 1232
rect 488828 814 488856 1226
rect 489840 898 489868 1634
rect 489840 870 489960 898
rect 489932 814 489960 870
rect 491312 814 491340 3334
rect 499764 3120 499816 3126
rect 499764 3062 499816 3068
rect 492680 2644 492732 2650
rect 492680 2586 492732 2592
rect 492128 2304 492180 2310
rect 492128 2246 492180 2252
rect 492140 1426 492168 2246
rect 492128 1420 492180 1426
rect 492128 1362 492180 1368
rect 492692 814 492720 2586
rect 494060 2032 494112 2038
rect 494060 1974 494112 1980
rect 494072 814 494100 1974
rect 496636 1624 496688 1630
rect 496636 1566 496688 1572
rect 495624 1556 495676 1562
rect 495624 1498 495676 1504
rect 494704 1352 494756 1358
rect 494704 1294 494756 1300
rect 494716 1086 494744 1294
rect 494704 1080 494756 1086
rect 494704 1022 494756 1028
rect 494520 1012 494572 1018
rect 494520 954 494572 960
rect 484584 808 484636 814
rect 484584 750 484636 756
rect 484676 808 484728 814
rect 484676 750 484728 756
rect 485780 808 485832 814
rect 485780 750 485832 756
rect 486884 808 486936 814
rect 486884 750 486936 756
rect 488632 808 488684 814
rect 488632 750 488684 756
rect 488816 808 488868 814
rect 488816 750 488868 756
rect 489920 808 489972 814
rect 489920 750 489972 756
rect 491300 808 491352 814
rect 491300 750 491352 756
rect 492680 808 492732 814
rect 492680 750 492732 756
rect 494060 808 494112 814
rect 494060 750 494112 756
rect 494532 746 494560 954
rect 495636 814 495664 1498
rect 496648 814 496676 1566
rect 499776 814 499804 3062
rect 530016 3003 530336 4066
rect 530016 2947 530028 3003
rect 530084 2947 530108 3003
rect 530164 2947 530188 3003
rect 530244 2947 530268 3003
rect 530324 2947 530336 3003
rect 530016 2923 530336 2947
rect 530016 2867 530028 2923
rect 530084 2867 530108 2923
rect 530164 2867 530188 2923
rect 530244 2867 530268 2923
rect 530324 2867 530336 2923
rect 530016 2843 530336 2867
rect 530016 2787 530028 2843
rect 530084 2787 530108 2843
rect 530164 2787 530188 2843
rect 530244 2787 530268 2843
rect 530324 2787 530336 2843
rect 530016 2763 530336 2787
rect 530016 2707 530028 2763
rect 530084 2707 530108 2763
rect 530164 2707 530188 2763
rect 530244 2707 530268 2763
rect 530324 2707 530336 2763
rect 505376 2576 505428 2582
rect 505376 2518 505428 2524
rect 500868 2304 500920 2310
rect 500868 2246 500920 2252
rect 500132 1216 500184 1222
rect 500132 1158 500184 1164
rect 500144 814 500172 1158
rect 500880 882 500908 2246
rect 502340 1760 502392 1766
rect 502340 1702 502392 1708
rect 500868 876 500920 882
rect 500868 818 500920 824
rect 502352 814 502380 1702
rect 505388 814 505416 2518
rect 530016 964 530336 2707
rect 530016 908 530028 964
rect 530084 908 530108 964
rect 530164 908 530188 964
rect 530244 908 530268 964
rect 530324 908 530336 964
rect 530016 884 530336 908
rect 530016 828 530028 884
rect 530084 828 530108 884
rect 530164 828 530188 884
rect 530244 828 530268 884
rect 530324 828 530336 884
rect 495624 808 495676 814
rect 495624 750 495676 756
rect 496636 808 496688 814
rect 496636 750 496688 756
rect 499764 808 499816 814
rect 499764 750 499816 756
rect 500132 808 500184 814
rect 500132 750 500184 756
rect 502340 808 502392 814
rect 502340 750 502392 756
rect 505376 808 505428 814
rect 505376 750 505428 756
rect 530016 804 530336 828
rect 530016 748 530028 804
rect 530084 748 530108 804
rect 530164 748 530188 804
rect 530244 748 530268 804
rect 530324 748 530336 804
rect 494520 740 494572 746
rect 494520 682 494572 688
rect 530016 724 530336 748
rect 530016 668 530028 724
rect 530084 668 530108 724
rect 530164 668 530188 724
rect 530244 668 530268 724
rect 530324 668 530336 724
rect 530016 656 530336 668
rect 530676 7740 530996 9488
rect 530676 7684 530688 7740
rect 530744 7684 530768 7740
rect 530824 7684 530848 7740
rect 530904 7684 530928 7740
rect 530984 7684 530996 7740
rect 530676 7660 530996 7684
rect 530676 7604 530688 7660
rect 530744 7604 530768 7660
rect 530824 7604 530848 7660
rect 530904 7604 530928 7660
rect 530984 7604 530996 7660
rect 530676 7580 530996 7604
rect 530676 7524 530688 7580
rect 530744 7524 530768 7580
rect 530824 7524 530848 7580
rect 530904 7524 530928 7580
rect 530984 7524 530996 7580
rect 530676 7500 530996 7524
rect 530676 7444 530688 7500
rect 530744 7444 530768 7500
rect 530824 7444 530848 7500
rect 530904 7444 530928 7500
rect 530984 7444 530996 7500
rect 530676 6381 530996 7444
rect 530676 6325 530688 6381
rect 530744 6325 530768 6381
rect 530824 6325 530848 6381
rect 530904 6325 530928 6381
rect 530984 6325 530996 6381
rect 530676 6301 530996 6325
rect 530676 6245 530688 6301
rect 530744 6245 530768 6301
rect 530824 6245 530848 6301
rect 530904 6245 530928 6301
rect 530984 6245 530996 6301
rect 530676 6221 530996 6245
rect 530676 6165 530688 6221
rect 530744 6165 530768 6221
rect 530824 6165 530848 6221
rect 530904 6165 530928 6221
rect 530984 6165 530996 6221
rect 530676 6141 530996 6165
rect 530676 6085 530688 6141
rect 530744 6085 530768 6141
rect 530824 6085 530848 6141
rect 530904 6085 530928 6141
rect 530984 6085 530996 6141
rect 530676 5022 530996 6085
rect 530676 4966 530688 5022
rect 530744 4966 530768 5022
rect 530824 4966 530848 5022
rect 530904 4966 530928 5022
rect 530984 4966 530996 5022
rect 530676 4942 530996 4966
rect 530676 4886 530688 4942
rect 530744 4886 530768 4942
rect 530824 4886 530848 4942
rect 530904 4886 530928 4942
rect 530984 4886 530996 4942
rect 530676 4862 530996 4886
rect 530676 4806 530688 4862
rect 530744 4806 530768 4862
rect 530824 4806 530848 4862
rect 530904 4806 530928 4862
rect 530984 4806 530996 4862
rect 530676 4782 530996 4806
rect 530676 4726 530688 4782
rect 530744 4726 530768 4782
rect 530824 4726 530848 4782
rect 530904 4726 530928 4782
rect 530984 4726 530996 4782
rect 530676 3663 530996 4726
rect 530676 3607 530688 3663
rect 530744 3607 530768 3663
rect 530824 3607 530848 3663
rect 530904 3607 530928 3663
rect 530984 3607 530996 3663
rect 530676 3583 530996 3607
rect 530676 3527 530688 3583
rect 530744 3527 530768 3583
rect 530824 3527 530848 3583
rect 530904 3527 530928 3583
rect 530984 3527 530996 3583
rect 530676 3503 530996 3527
rect 530676 3447 530688 3503
rect 530744 3447 530768 3503
rect 530824 3447 530848 3503
rect 530904 3447 530928 3503
rect 530984 3447 530996 3503
rect 530676 3423 530996 3447
rect 530676 3367 530688 3423
rect 530744 3367 530768 3423
rect 530824 3367 530848 3423
rect 530904 3367 530928 3423
rect 530984 3367 530996 3423
rect 479706 504 479762 513
rect 479706 439 479762 448
rect 482650 504 482706 513
rect 482650 439 482706 448
rect 479720 66 479748 439
rect 530676 304 530996 3367
rect 530676 248 530688 304
rect 530744 248 530768 304
rect 530824 248 530848 304
rect 530904 248 530928 304
rect 530984 248 530996 304
rect 530676 224 530996 248
rect 530676 168 530688 224
rect 530744 168 530768 224
rect 530824 168 530848 224
rect 530904 168 530928 224
rect 530984 168 530996 224
rect 530676 144 530996 168
rect 530676 88 530688 144
rect 530744 88 530768 144
rect 530824 88 530848 144
rect 530904 88 530928 144
rect 530984 88 530996 144
rect 463352 8 463364 64
rect 463420 8 463444 64
rect 463500 8 463524 64
rect 463580 8 463604 64
rect 463660 8 463672 64
rect 463352 -4 463672 8
rect 470692 60 470744 66
rect 470692 2 470744 8
rect 479708 60 479760 66
rect 479708 2 479760 8
rect 530676 64 530996 88
rect 530676 8 530688 64
rect 530744 8 530768 64
rect 530824 8 530848 64
rect 530904 8 530928 64
rect 530984 8 530996 64
rect 530676 -4 530996 8
<< via2 >>
rect -1064 9728 -1008 9784
rect -984 9728 -928 9784
rect -904 9728 -848 9784
rect -824 9728 -768 9784
rect -1064 9648 -1008 9704
rect -984 9648 -928 9704
rect -904 9648 -848 9704
rect -824 9648 -768 9704
rect -1064 9568 -1008 9624
rect -984 9568 -928 9624
rect -904 9568 -848 9624
rect -824 9568 -768 9624
rect -1064 9488 -1008 9544
rect -984 9488 -928 9544
rect -904 9488 -848 9544
rect -824 9488 -768 9544
rect -1064 7684 -1008 7740
rect -984 7684 -928 7740
rect -904 7684 -848 7740
rect -824 7684 -768 7740
rect -1064 7604 -1008 7660
rect -984 7604 -928 7660
rect -904 7604 -848 7660
rect -824 7604 -768 7660
rect -1064 7524 -1008 7580
rect -984 7524 -928 7580
rect -904 7524 -848 7580
rect -824 7524 -768 7580
rect -1064 7444 -1008 7500
rect -984 7444 -928 7500
rect -904 7444 -848 7500
rect -824 7444 -768 7500
rect -1064 6325 -1008 6381
rect -984 6325 -928 6381
rect -904 6325 -848 6381
rect -824 6325 -768 6381
rect -1064 6245 -1008 6301
rect -984 6245 -928 6301
rect -904 6245 -848 6301
rect -824 6245 -768 6301
rect -1064 6165 -1008 6221
rect -984 6165 -928 6221
rect -904 6165 -848 6221
rect -824 6165 -768 6221
rect -1064 6085 -1008 6141
rect -984 6085 -928 6141
rect -904 6085 -848 6141
rect -824 6085 -768 6141
rect -1064 4966 -1008 5022
rect -984 4966 -928 5022
rect -904 4966 -848 5022
rect -824 4966 -768 5022
rect -1064 4886 -1008 4942
rect -984 4886 -928 4942
rect -904 4886 -848 4942
rect -824 4886 -768 4942
rect -1064 4806 -1008 4862
rect -984 4806 -928 4862
rect -904 4806 -848 4862
rect -824 4806 -768 4862
rect -1064 4726 -1008 4782
rect -984 4726 -928 4782
rect -904 4726 -848 4782
rect -824 4726 -768 4782
rect -1064 3607 -1008 3663
rect -984 3607 -928 3663
rect -904 3607 -848 3663
rect -824 3607 -768 3663
rect -1064 3527 -1008 3583
rect -984 3527 -928 3583
rect -904 3527 -848 3583
rect -824 3527 -768 3583
rect -1064 3447 -1008 3503
rect -984 3447 -928 3503
rect -904 3447 -848 3503
rect -824 3447 -768 3503
rect -1064 3367 -1008 3423
rect -984 3367 -928 3423
rect -904 3367 -848 3423
rect -824 3367 -768 3423
rect -404 9068 -348 9124
rect -324 9068 -268 9124
rect -244 9068 -188 9124
rect -164 9068 -108 9124
rect -404 8988 -348 9044
rect -324 8988 -268 9044
rect -244 8988 -188 9044
rect -164 8988 -108 9044
rect -404 8908 -348 8964
rect -324 8908 -268 8964
rect -244 8908 -188 8964
rect -164 8908 -108 8964
rect -404 8828 -348 8884
rect -324 8828 -268 8884
rect -244 8828 -188 8884
rect -164 8828 -108 8884
rect -404 7024 -348 7080
rect -324 7024 -268 7080
rect -244 7024 -188 7080
rect -164 7024 -108 7080
rect -404 6944 -348 7000
rect -324 6944 -268 7000
rect -244 6944 -188 7000
rect -164 6944 -108 7000
rect -404 6864 -348 6920
rect -324 6864 -268 6920
rect -244 6864 -188 6920
rect -164 6864 -108 6920
rect -404 6784 -348 6840
rect -324 6784 -268 6840
rect -244 6784 -188 6840
rect -164 6784 -108 6840
rect -404 5665 -348 5721
rect -324 5665 -268 5721
rect -244 5665 -188 5721
rect -164 5665 -108 5721
rect -404 5585 -348 5641
rect -324 5585 -268 5641
rect -244 5585 -188 5641
rect -164 5585 -108 5641
rect -404 5505 -348 5561
rect -324 5505 -268 5561
rect -244 5505 -188 5561
rect -164 5505 -108 5561
rect -404 5425 -348 5481
rect -324 5425 -268 5481
rect -244 5425 -188 5481
rect -164 5425 -108 5481
rect -404 4306 -348 4362
rect -324 4306 -268 4362
rect -244 4306 -188 4362
rect -164 4306 -108 4362
rect -404 4226 -348 4282
rect -324 4226 -268 4282
rect -244 4226 -188 4282
rect -164 4226 -108 4282
rect -404 4146 -348 4202
rect -324 4146 -268 4202
rect -244 4146 -188 4202
rect -164 4146 -108 4202
rect -404 4066 -348 4122
rect -324 4066 -268 4122
rect -244 4066 -188 4122
rect -164 4066 -108 4122
rect -404 2947 -348 3003
rect -324 2947 -268 3003
rect -244 2947 -188 3003
rect -164 2947 -108 3003
rect -404 2867 -348 2923
rect -324 2867 -268 2923
rect -244 2867 -188 2923
rect -164 2867 -108 2923
rect -404 2787 -348 2843
rect -324 2787 -268 2843
rect -244 2787 -188 2843
rect -164 2787 -108 2843
rect -404 2707 -348 2763
rect -324 2707 -268 2763
rect -244 2707 -188 2763
rect -164 2707 -108 2763
rect -404 908 -348 964
rect -324 908 -268 964
rect -244 908 -188 964
rect -164 908 -108 964
rect -404 828 -348 884
rect -324 828 -268 884
rect -244 828 -188 884
rect -164 828 -108 884
rect -404 748 -348 804
rect -324 748 -268 804
rect -244 748 -188 804
rect -164 748 -108 804
rect -404 668 -348 724
rect -324 668 -268 724
rect -244 668 -188 724
rect -164 668 -108 724
rect 26054 1536 26110 1592
rect 26974 1400 27030 1456
rect 28538 1148 28594 1184
rect 28538 1128 28540 1148
rect 28540 1128 28592 1148
rect 28592 1128 28594 1148
rect 29090 1808 29146 1864
rect 31206 1672 31262 1728
rect 28630 468 28686 504
rect 28630 448 28632 468
rect 28632 448 28684 468
rect 28684 448 28686 468
rect -1064 248 -1008 304
rect -984 248 -928 304
rect -904 248 -848 304
rect -824 248 -768 304
rect -1064 168 -1008 224
rect -984 168 -928 224
rect -904 168 -848 224
rect -824 168 -768 224
rect 31206 1284 31262 1320
rect 31206 1264 31208 1284
rect 31208 1264 31260 1284
rect 31260 1264 31262 1284
rect 66920 9068 66976 9124
rect 67000 9068 67056 9124
rect 67080 9068 67136 9124
rect 67160 9068 67216 9124
rect 66920 8988 66976 9044
rect 67000 8988 67056 9044
rect 67080 8988 67136 9044
rect 67160 8988 67216 9044
rect 66920 8908 66976 8964
rect 67000 8908 67056 8964
rect 67080 8908 67136 8964
rect 67160 8908 67216 8964
rect 66920 8828 66976 8884
rect 67000 8828 67056 8884
rect 67080 8828 67136 8884
rect 67160 8828 67216 8884
rect 66920 7046 66966 7080
rect 66966 7046 66976 7080
rect 67000 7046 67030 7080
rect 67030 7046 67042 7080
rect 67042 7046 67056 7080
rect 67080 7046 67094 7080
rect 67094 7046 67106 7080
rect 67106 7046 67136 7080
rect 67160 7046 67170 7080
rect 67170 7046 67216 7080
rect 66920 7024 66976 7046
rect 67000 7024 67056 7046
rect 67080 7024 67136 7046
rect 67160 7024 67216 7046
rect 66920 6944 66976 7000
rect 67000 6944 67056 7000
rect 67080 6944 67136 7000
rect 67160 6944 67216 7000
rect 66920 6864 66976 6920
rect 67000 6864 67056 6920
rect 67080 6864 67136 6920
rect 67160 6864 67216 6920
rect 66920 6784 66976 6840
rect 67000 6784 67056 6840
rect 67080 6784 67136 6840
rect 67160 6784 67216 6840
rect 66920 5665 66976 5721
rect 67000 5665 67056 5721
rect 67080 5665 67136 5721
rect 67160 5665 67216 5721
rect 66920 5585 66976 5641
rect 67000 5585 67056 5641
rect 67080 5585 67136 5641
rect 67160 5585 67216 5641
rect 66920 5505 66976 5561
rect 67000 5505 67056 5561
rect 67080 5505 67136 5561
rect 67160 5505 67216 5561
rect 66920 5425 66976 5481
rect 67000 5425 67056 5481
rect 67080 5425 67136 5481
rect 67160 5425 67216 5481
rect 54666 2488 54722 2544
rect 36726 1944 36782 2000
rect 66920 4306 66976 4362
rect 67000 4306 67056 4362
rect 67080 4306 67136 4362
rect 67160 4306 67216 4362
rect 66920 4226 66976 4282
rect 67000 4226 67056 4282
rect 67080 4226 67136 4282
rect 67160 4226 67216 4282
rect 66920 4146 66976 4202
rect 67000 4146 67056 4202
rect 67080 4146 67136 4202
rect 67160 4146 67216 4202
rect 66920 4066 66976 4122
rect 67000 4066 67056 4122
rect 67080 4066 67136 4122
rect 67160 4066 67216 4122
rect 66920 2947 66976 3003
rect 67000 2947 67056 3003
rect 67080 2947 67136 3003
rect 67160 2947 67216 3003
rect 66920 2867 66976 2923
rect 67000 2867 67056 2923
rect 67080 2867 67136 2923
rect 67160 2867 67216 2923
rect 66920 2787 66976 2843
rect 67000 2787 67056 2843
rect 67080 2787 67136 2843
rect 67160 2787 67216 2843
rect 66920 2746 66976 2763
rect 67000 2746 67056 2763
rect 67080 2746 67136 2763
rect 67160 2746 67216 2763
rect 66920 2707 66966 2746
rect 66966 2707 66976 2746
rect 67000 2707 67030 2746
rect 67030 2707 67042 2746
rect 67042 2707 67056 2746
rect 67080 2707 67094 2746
rect 67094 2707 67106 2746
rect 67106 2707 67136 2746
rect 67160 2707 67170 2746
rect 67170 2707 67216 2746
rect 36542 1808 36598 1864
rect 33782 1672 33838 1728
rect 32862 1536 32918 1592
rect 31850 1400 31906 1456
rect 31758 1264 31814 1320
rect 31574 1128 31630 1184
rect -1064 88 -1008 144
rect -984 88 -928 144
rect -904 88 -848 144
rect -824 88 -768 144
rect 66920 908 66976 964
rect 67000 908 67056 964
rect 67080 908 67136 964
rect 67160 908 67216 964
rect 66920 828 66976 884
rect 67000 828 67056 884
rect 67080 828 67136 884
rect 67160 828 67216 884
rect 66920 748 66976 804
rect 67000 748 67056 804
rect 67080 748 67136 804
rect 67160 748 67216 804
rect 66920 668 66976 724
rect 67000 668 67056 724
rect 67080 668 67136 724
rect 67160 668 67216 724
rect -1064 8 -1008 64
rect -984 8 -928 64
rect -904 8 -848 64
rect -824 8 -768 64
rect 67580 9728 67636 9784
rect 67660 9728 67716 9784
rect 67740 9728 67796 9784
rect 67820 9728 67876 9784
rect 67580 9648 67636 9704
rect 67660 9648 67716 9704
rect 67740 9648 67796 9704
rect 67820 9648 67876 9704
rect 67580 9568 67636 9624
rect 67660 9568 67716 9624
rect 67740 9568 67796 9624
rect 67820 9568 67876 9624
rect 67580 9488 67636 9544
rect 67660 9488 67716 9544
rect 67740 9488 67796 9544
rect 67820 9488 67876 9544
rect 67580 7684 67636 7740
rect 67660 7684 67716 7740
rect 67740 7684 67796 7740
rect 67820 7684 67876 7740
rect 67580 7642 67636 7660
rect 67660 7642 67716 7660
rect 67740 7642 67796 7660
rect 67820 7642 67876 7660
rect 67580 7604 67626 7642
rect 67626 7604 67636 7642
rect 67660 7604 67690 7642
rect 67690 7604 67702 7642
rect 67702 7604 67716 7642
rect 67740 7604 67754 7642
rect 67754 7604 67766 7642
rect 67766 7604 67796 7642
rect 67820 7604 67830 7642
rect 67830 7604 67876 7642
rect 67580 7524 67636 7580
rect 67660 7524 67716 7580
rect 67740 7524 67796 7580
rect 67820 7524 67876 7580
rect 67580 7444 67636 7500
rect 67660 7444 67716 7500
rect 67740 7444 67796 7500
rect 67820 7444 67876 7500
rect 67580 6325 67636 6381
rect 67660 6325 67716 6381
rect 67740 6325 67796 6381
rect 67820 6325 67876 6381
rect 67580 6245 67636 6301
rect 67660 6245 67716 6301
rect 67740 6245 67796 6301
rect 67820 6245 67876 6301
rect 67580 6165 67636 6221
rect 67660 6165 67716 6221
rect 67740 6165 67796 6221
rect 67820 6165 67876 6221
rect 67580 6085 67636 6141
rect 67660 6085 67716 6141
rect 67740 6085 67796 6141
rect 67820 6085 67876 6141
rect 67580 4966 67636 5022
rect 67660 4966 67716 5022
rect 67740 4966 67796 5022
rect 67820 4966 67876 5022
rect 67580 4886 67636 4942
rect 67660 4886 67716 4942
rect 67740 4886 67796 4942
rect 67820 4886 67876 4942
rect 67580 4806 67636 4862
rect 67660 4806 67716 4862
rect 67740 4806 67796 4862
rect 67820 4806 67876 4862
rect 67580 4726 67636 4782
rect 67660 4726 67716 4782
rect 67740 4726 67796 4782
rect 67820 4726 67876 4782
rect 67580 3607 67636 3663
rect 67660 3607 67716 3663
rect 67740 3607 67796 3663
rect 67820 3607 67876 3663
rect 67580 3527 67636 3583
rect 67660 3527 67716 3583
rect 67740 3527 67796 3583
rect 67820 3527 67876 3583
rect 67580 3447 67636 3503
rect 67660 3447 67716 3503
rect 67740 3447 67796 3503
rect 67820 3447 67876 3503
rect 67580 3367 67636 3423
rect 67660 3367 67716 3423
rect 67740 3367 67796 3423
rect 67820 3367 67876 3423
rect 107658 2388 107660 2408
rect 107660 2388 107712 2408
rect 107712 2388 107714 2408
rect 107658 2352 107714 2388
rect 67580 248 67636 304
rect 67660 248 67716 304
rect 67740 248 67796 304
rect 67820 248 67876 304
rect 67580 168 67636 224
rect 67660 168 67716 224
rect 67740 168 67796 224
rect 67820 168 67876 224
rect 122562 3168 122618 3224
rect 122654 2216 122710 2272
rect 123206 2080 123262 2136
rect 122930 448 122986 504
rect 67580 88 67636 144
rect 67660 88 67716 144
rect 67740 88 67796 144
rect 67820 88 67876 144
rect 198848 9068 198904 9124
rect 198928 9068 198984 9124
rect 199008 9068 199064 9124
rect 199088 9068 199144 9124
rect 198848 8988 198904 9044
rect 198928 8988 198984 9044
rect 199008 8988 199064 9044
rect 199088 8988 199144 9044
rect 198848 8908 198904 8964
rect 198928 8908 198984 8964
rect 199008 8908 199064 8964
rect 199088 8908 199144 8964
rect 198848 8828 198904 8884
rect 198928 8828 198984 8884
rect 199008 8828 199064 8884
rect 199088 8828 199144 8884
rect 198848 7046 198894 7080
rect 198894 7046 198904 7080
rect 198928 7046 198958 7080
rect 198958 7046 198970 7080
rect 198970 7046 198984 7080
rect 199008 7046 199022 7080
rect 199022 7046 199034 7080
rect 199034 7046 199064 7080
rect 199088 7046 199098 7080
rect 199098 7046 199144 7080
rect 198848 7024 198904 7046
rect 198928 7024 198984 7046
rect 199008 7024 199064 7046
rect 199088 7024 199144 7046
rect 198848 6944 198904 7000
rect 198928 6944 198984 7000
rect 199008 6944 199064 7000
rect 199088 6944 199144 7000
rect 198848 6864 198904 6920
rect 198928 6864 198984 6920
rect 199008 6864 199064 6920
rect 199088 6864 199144 6920
rect 198848 6784 198904 6840
rect 198928 6784 198984 6840
rect 199008 6784 199064 6840
rect 199088 6784 199144 6840
rect 148230 2524 148232 2544
rect 148232 2524 148284 2544
rect 148284 2524 148286 2544
rect 148230 2488 148286 2524
rect 130198 1944 130254 2000
rect 198848 5665 198904 5721
rect 198928 5665 198984 5721
rect 199008 5665 199064 5721
rect 199088 5665 199144 5721
rect 198848 5585 198904 5641
rect 198928 5585 198984 5641
rect 199008 5585 199064 5641
rect 199088 5585 199144 5641
rect 198848 5505 198904 5561
rect 198928 5505 198984 5561
rect 199008 5505 199064 5561
rect 199088 5505 199144 5561
rect 198848 5425 198904 5481
rect 198928 5425 198984 5481
rect 199008 5425 199064 5481
rect 199088 5425 199144 5481
rect 198848 4306 198904 4362
rect 198928 4306 198984 4362
rect 199008 4306 199064 4362
rect 199088 4306 199144 4362
rect 198848 4226 198904 4282
rect 198928 4226 198984 4282
rect 199008 4226 199064 4282
rect 199088 4226 199144 4282
rect 198848 4146 198904 4202
rect 198928 4146 198984 4202
rect 199008 4146 199064 4202
rect 199088 4146 199144 4202
rect 198848 4066 198904 4122
rect 198928 4066 198984 4122
rect 199008 4066 199064 4122
rect 199088 4066 199144 4122
rect 198848 2947 198904 3003
rect 198928 2947 198984 3003
rect 199008 2947 199064 3003
rect 199088 2947 199144 3003
rect 198848 2867 198904 2923
rect 198928 2867 198984 2923
rect 199008 2867 199064 2923
rect 199088 2867 199144 2923
rect 198848 2787 198904 2843
rect 198928 2787 198984 2843
rect 199008 2787 199064 2843
rect 199088 2787 199144 2843
rect 198848 2746 198904 2763
rect 198928 2746 198984 2763
rect 199008 2746 199064 2763
rect 199088 2746 199144 2763
rect 198848 2707 198894 2746
rect 198894 2707 198904 2746
rect 198928 2707 198958 2746
rect 198958 2707 198970 2746
rect 198970 2707 198984 2746
rect 199008 2707 199022 2746
rect 199022 2707 199034 2746
rect 199034 2707 199064 2746
rect 199088 2707 199098 2746
rect 199098 2707 199144 2746
rect 199508 9728 199564 9784
rect 199588 9728 199644 9784
rect 199668 9728 199724 9784
rect 199748 9728 199804 9784
rect 199508 9648 199564 9704
rect 199588 9648 199644 9704
rect 199668 9648 199724 9704
rect 199748 9648 199804 9704
rect 199508 9568 199564 9624
rect 199588 9568 199644 9624
rect 199668 9568 199724 9624
rect 199748 9568 199804 9624
rect 199508 9488 199564 9544
rect 199588 9488 199644 9544
rect 199668 9488 199724 9544
rect 199748 9488 199804 9544
rect 199508 7684 199564 7740
rect 199588 7684 199644 7740
rect 199668 7684 199724 7740
rect 199748 7684 199804 7740
rect 199508 7642 199564 7660
rect 199588 7642 199644 7660
rect 199668 7642 199724 7660
rect 199748 7642 199804 7660
rect 199508 7604 199554 7642
rect 199554 7604 199564 7642
rect 199588 7604 199618 7642
rect 199618 7604 199630 7642
rect 199630 7604 199644 7642
rect 199668 7604 199682 7642
rect 199682 7604 199694 7642
rect 199694 7604 199724 7642
rect 199748 7604 199758 7642
rect 199758 7604 199804 7642
rect 199508 7524 199564 7580
rect 199588 7524 199644 7580
rect 199668 7524 199724 7580
rect 199748 7524 199804 7580
rect 199508 7444 199564 7500
rect 199588 7444 199644 7500
rect 199668 7444 199724 7500
rect 199748 7444 199804 7500
rect 199508 6325 199564 6381
rect 199588 6325 199644 6381
rect 199668 6325 199724 6381
rect 199748 6325 199804 6381
rect 199508 6245 199564 6301
rect 199588 6245 199644 6301
rect 199668 6245 199724 6301
rect 199748 6245 199804 6301
rect 199508 6165 199564 6221
rect 199588 6165 199644 6221
rect 199668 6165 199724 6221
rect 199748 6165 199804 6221
rect 199508 6085 199564 6141
rect 199588 6085 199644 6141
rect 199668 6085 199724 6141
rect 199748 6085 199804 6141
rect 199508 4966 199564 5022
rect 199588 4966 199644 5022
rect 199668 4966 199724 5022
rect 199748 4966 199804 5022
rect 199508 4886 199564 4942
rect 199588 4886 199644 4942
rect 199668 4886 199724 4942
rect 199748 4886 199804 4942
rect 199508 4806 199564 4862
rect 199588 4806 199644 4862
rect 199668 4806 199724 4862
rect 199748 4806 199804 4862
rect 199508 4726 199564 4782
rect 199588 4726 199644 4782
rect 199668 4726 199724 4782
rect 199748 4726 199804 4782
rect 199508 3607 199564 3663
rect 199588 3607 199644 3663
rect 199668 3607 199724 3663
rect 199748 3607 199804 3663
rect 199508 3527 199564 3583
rect 199588 3527 199644 3583
rect 199668 3527 199724 3583
rect 199748 3527 199804 3583
rect 199508 3447 199564 3503
rect 199588 3447 199644 3503
rect 199668 3447 199724 3503
rect 199748 3447 199804 3503
rect 199508 3367 199564 3423
rect 199588 3367 199644 3423
rect 199668 3367 199724 3423
rect 199748 3367 199804 3423
rect 201682 2352 201738 2408
rect 198848 908 198904 964
rect 198928 908 198984 964
rect 199008 908 199064 964
rect 199088 908 199144 964
rect 198848 828 198904 884
rect 198928 828 198984 884
rect 199008 828 199064 884
rect 199088 828 199144 884
rect 198848 748 198904 804
rect 198928 748 198984 804
rect 199008 748 199064 804
rect 199088 748 199144 804
rect 198848 668 198904 724
rect 198928 668 198984 724
rect 199008 668 199064 724
rect 199088 668 199144 724
rect 67580 8 67636 64
rect 67660 8 67716 64
rect 67740 8 67796 64
rect 67820 8 67876 64
rect 213550 2352 213606 2408
rect 214286 3848 214342 3904
rect 214010 2216 214066 2272
rect 215390 2080 215446 2136
rect 199508 248 199564 304
rect 199588 248 199644 304
rect 199668 248 199724 304
rect 199748 248 199804 304
rect 199508 168 199564 224
rect 199588 168 199644 224
rect 199668 168 199724 224
rect 199748 168 199804 224
rect 216678 3168 216734 3224
rect 330776 9068 330832 9124
rect 330856 9068 330912 9124
rect 330936 9068 330992 9124
rect 331016 9068 331072 9124
rect 330776 8988 330832 9044
rect 330856 8988 330912 9044
rect 330936 8988 330992 9044
rect 331016 8988 331072 9044
rect 224222 2080 224278 2136
rect 260286 1944 260342 2000
rect 296994 2488 297050 2544
rect 300766 2216 300822 2272
rect 303986 1808 304042 1864
rect 307666 448 307722 504
rect 310886 3848 310942 3904
rect 310702 2388 310704 2408
rect 310704 2388 310756 2408
rect 310756 2388 310758 2408
rect 310702 2352 310758 2388
rect 330776 8908 330832 8964
rect 330856 8908 330912 8964
rect 330936 8908 330992 8964
rect 331016 8908 331072 8964
rect 330776 8828 330832 8884
rect 330856 8828 330912 8884
rect 330936 8828 330992 8884
rect 331016 8828 331072 8884
rect 330776 7046 330822 7080
rect 330822 7046 330832 7080
rect 330856 7046 330886 7080
rect 330886 7046 330898 7080
rect 330898 7046 330912 7080
rect 330936 7046 330950 7080
rect 330950 7046 330962 7080
rect 330962 7046 330992 7080
rect 331016 7046 331026 7080
rect 331026 7046 331072 7080
rect 330776 7024 330832 7046
rect 330856 7024 330912 7046
rect 330936 7024 330992 7046
rect 331016 7024 331072 7046
rect 330776 6944 330832 7000
rect 330856 6944 330912 7000
rect 330936 6944 330992 7000
rect 331016 6944 331072 7000
rect 330776 6864 330832 6920
rect 330856 6864 330912 6920
rect 330936 6864 330992 6920
rect 331016 6864 331072 6920
rect 330776 6784 330832 6840
rect 330856 6784 330912 6840
rect 330936 6784 330992 6840
rect 331016 6784 331072 6840
rect 199508 88 199564 144
rect 199588 88 199644 144
rect 199668 88 199724 144
rect 199748 88 199804 144
rect 317050 2080 317106 2136
rect 330776 5665 330832 5721
rect 330856 5665 330912 5721
rect 330936 5665 330992 5721
rect 331016 5665 331072 5721
rect 330776 5585 330832 5641
rect 330856 5585 330912 5641
rect 330936 5585 330992 5641
rect 331016 5585 331072 5641
rect 330776 5505 330832 5561
rect 330856 5505 330912 5561
rect 330936 5505 330992 5561
rect 331016 5505 331072 5561
rect 330776 5425 330832 5481
rect 330856 5425 330912 5481
rect 330936 5425 330992 5481
rect 331016 5425 331072 5481
rect 330776 4306 330832 4362
rect 330856 4306 330912 4362
rect 330936 4306 330992 4362
rect 331016 4306 331072 4362
rect 330776 4226 330832 4282
rect 330856 4226 330912 4282
rect 330936 4226 330992 4282
rect 331016 4226 331072 4282
rect 330776 4146 330832 4202
rect 330856 4146 330912 4202
rect 330936 4146 330992 4202
rect 331016 4146 331072 4202
rect 330776 4066 330832 4122
rect 330856 4066 330912 4122
rect 330936 4066 330992 4122
rect 331016 4066 331072 4122
rect 331436 9728 331492 9784
rect 331516 9728 331572 9784
rect 331596 9728 331652 9784
rect 331676 9728 331732 9784
rect 331436 9648 331492 9704
rect 331516 9648 331572 9704
rect 331596 9648 331652 9704
rect 331676 9648 331732 9704
rect 331436 9568 331492 9624
rect 331516 9568 331572 9624
rect 331596 9568 331652 9624
rect 331676 9568 331732 9624
rect 331436 9488 331492 9544
rect 331516 9488 331572 9544
rect 331596 9488 331652 9544
rect 331676 9488 331732 9544
rect 331436 7684 331492 7740
rect 331516 7684 331572 7740
rect 331596 7684 331652 7740
rect 331676 7684 331732 7740
rect 331436 7642 331492 7660
rect 331516 7642 331572 7660
rect 331596 7642 331652 7660
rect 331676 7642 331732 7660
rect 331436 7604 331482 7642
rect 331482 7604 331492 7642
rect 331516 7604 331546 7642
rect 331546 7604 331558 7642
rect 331558 7604 331572 7642
rect 331596 7604 331610 7642
rect 331610 7604 331622 7642
rect 331622 7604 331652 7642
rect 331676 7604 331686 7642
rect 331686 7604 331732 7642
rect 331436 7524 331492 7580
rect 331516 7524 331572 7580
rect 331596 7524 331652 7580
rect 331676 7524 331732 7580
rect 331436 7444 331492 7500
rect 331516 7444 331572 7500
rect 331596 7444 331652 7500
rect 331676 7444 331732 7500
rect 331436 6325 331492 6381
rect 331516 6325 331572 6381
rect 331596 6325 331652 6381
rect 331676 6325 331732 6381
rect 331436 6245 331492 6301
rect 331516 6245 331572 6301
rect 331596 6245 331652 6301
rect 331676 6245 331732 6301
rect 331436 6165 331492 6221
rect 331516 6165 331572 6221
rect 331596 6165 331652 6221
rect 331676 6165 331732 6221
rect 331436 6085 331492 6141
rect 331516 6085 331572 6141
rect 331596 6085 331652 6141
rect 331676 6085 331732 6141
rect 331436 4966 331492 5022
rect 331516 4966 331572 5022
rect 331596 4966 331652 5022
rect 331676 4966 331732 5022
rect 331436 4886 331492 4942
rect 331516 4886 331572 4942
rect 331596 4886 331652 4942
rect 331676 4886 331732 4942
rect 331436 4806 331492 4862
rect 331516 4806 331572 4862
rect 331596 4806 331652 4862
rect 331676 4806 331732 4862
rect 331436 4726 331492 4782
rect 331516 4726 331572 4782
rect 331596 4726 331652 4782
rect 331676 4726 331732 4782
rect 331436 3607 331492 3663
rect 331516 3607 331572 3663
rect 331596 3607 331652 3663
rect 331676 3607 331732 3663
rect 331436 3527 331492 3583
rect 331516 3527 331572 3583
rect 331596 3527 331652 3583
rect 331676 3527 331732 3583
rect 331436 3447 331492 3503
rect 331516 3447 331572 3503
rect 331596 3447 331652 3503
rect 331676 3447 331732 3503
rect 331436 3367 331492 3423
rect 331516 3367 331572 3423
rect 331596 3367 331652 3423
rect 331676 3367 331732 3423
rect 330776 2947 330832 3003
rect 330856 2947 330912 3003
rect 330936 2947 330992 3003
rect 331016 2947 331072 3003
rect 330776 2867 330832 2923
rect 330856 2867 330912 2923
rect 330936 2867 330992 2923
rect 331016 2867 331072 2923
rect 330776 2787 330832 2843
rect 330856 2787 330912 2843
rect 330936 2787 330992 2843
rect 331016 2787 331072 2843
rect 330776 2746 330832 2763
rect 330856 2746 330912 2763
rect 330936 2746 330992 2763
rect 331016 2746 331072 2763
rect 330776 2707 330822 2746
rect 330822 2707 330832 2746
rect 330856 2707 330886 2746
rect 330886 2707 330898 2746
rect 330898 2707 330912 2746
rect 330936 2707 330950 2746
rect 330950 2707 330962 2746
rect 330962 2707 330992 2746
rect 331016 2707 331026 2746
rect 331026 2707 331072 2746
rect 330776 908 330832 964
rect 330856 908 330912 964
rect 330936 908 330992 964
rect 331016 908 331072 964
rect 330776 828 330832 884
rect 330856 828 330912 884
rect 330936 828 330992 884
rect 331016 828 331072 884
rect 330776 748 330832 804
rect 330856 748 330912 804
rect 330936 748 330992 804
rect 331016 748 331072 804
rect 330776 668 330832 724
rect 330856 668 330912 724
rect 330936 668 330992 724
rect 331016 668 331072 724
rect 199508 8 199564 64
rect 199588 8 199644 64
rect 199668 8 199724 64
rect 199748 8 199804 64
rect 331436 248 331492 304
rect 331516 248 331572 304
rect 331596 248 331652 304
rect 331676 248 331732 304
rect 331436 168 331492 224
rect 331516 168 331572 224
rect 331596 168 331652 224
rect 331676 168 331732 224
rect 331436 88 331492 144
rect 331516 88 331572 144
rect 331596 88 331652 144
rect 331676 88 331732 144
rect 353298 1944 353354 2000
rect 391110 2488 391166 2544
rect 355966 2080 356022 2136
rect 372434 2372 372490 2408
rect 372434 2352 372436 2372
rect 372436 2352 372488 2372
rect 372488 2352 372490 2372
rect 390558 1944 390614 2000
rect 394422 2216 394478 2272
rect 396078 2488 396134 2544
rect 396906 1808 396962 1864
rect 400770 2488 400826 2544
rect 399482 1672 399538 1728
rect 399298 1536 399354 1592
rect 398010 1400 398066 1456
rect 399022 1400 399078 1456
rect 398838 1264 398894 1320
rect 399666 1264 399722 1320
rect 399850 1128 399906 1184
rect 402610 1536 402666 1592
rect 404266 1264 404322 1320
rect 404818 1400 404874 1456
rect 400494 468 400550 504
rect 400494 448 400496 468
rect 400496 448 400548 468
rect 400548 448 400550 468
rect 400678 448 400734 504
rect 403438 484 403440 504
rect 403440 484 403492 504
rect 403492 484 403494 504
rect 403438 448 403494 484
rect 407486 1300 407488 1320
rect 407488 1300 407540 1320
rect 407540 1300 407542 1320
rect 407486 1264 407542 1300
rect 407486 1148 407542 1184
rect 407486 1128 407488 1148
rect 407488 1128 407540 1148
rect 407540 1128 407542 1148
rect 408590 1672 408646 1728
rect 410798 1264 410854 1320
rect 462704 9068 462760 9124
rect 462784 9068 462840 9124
rect 462864 9068 462920 9124
rect 462944 9068 463000 9124
rect 462704 8988 462760 9044
rect 462784 8988 462840 9044
rect 462864 8988 462920 9044
rect 462944 8988 463000 9044
rect 462704 8908 462760 8964
rect 462784 8908 462840 8964
rect 462864 8908 462920 8964
rect 462944 8908 463000 8964
rect 462704 8828 462760 8884
rect 462784 8828 462840 8884
rect 462864 8828 462920 8884
rect 462944 8828 463000 8884
rect 462704 7046 462750 7080
rect 462750 7046 462760 7080
rect 462784 7046 462814 7080
rect 462814 7046 462826 7080
rect 462826 7046 462840 7080
rect 462864 7046 462878 7080
rect 462878 7046 462890 7080
rect 462890 7046 462920 7080
rect 462944 7046 462954 7080
rect 462954 7046 463000 7080
rect 462704 7024 462760 7046
rect 462784 7024 462840 7046
rect 462864 7024 462920 7046
rect 462944 7024 463000 7046
rect 462704 6944 462760 7000
rect 462784 6944 462840 7000
rect 462864 6944 462920 7000
rect 462944 6944 463000 7000
rect 462704 6864 462760 6920
rect 462784 6864 462840 6920
rect 462864 6864 462920 6920
rect 462944 6864 463000 6920
rect 462704 6784 462760 6840
rect 462784 6784 462840 6840
rect 462864 6784 462920 6840
rect 462944 6784 463000 6840
rect 462704 5665 462760 5721
rect 462784 5665 462840 5721
rect 462864 5665 462920 5721
rect 462944 5665 463000 5721
rect 462704 5585 462760 5641
rect 462784 5585 462840 5641
rect 462864 5585 462920 5641
rect 462944 5585 463000 5641
rect 462704 5505 462760 5561
rect 462784 5505 462840 5561
rect 462864 5505 462920 5561
rect 462944 5505 463000 5561
rect 462704 5425 462760 5481
rect 462784 5425 462840 5481
rect 462864 5425 462920 5481
rect 462944 5425 463000 5481
rect 435454 1944 435510 2000
rect 439410 2080 439466 2136
rect 462704 4306 462760 4362
rect 462784 4306 462840 4362
rect 462864 4306 462920 4362
rect 462944 4306 463000 4362
rect 462704 4226 462760 4282
rect 462784 4226 462840 4282
rect 462864 4226 462920 4282
rect 462944 4226 463000 4282
rect 462704 4146 462760 4202
rect 462784 4146 462840 4202
rect 462864 4146 462920 4202
rect 462944 4146 463000 4202
rect 462704 4066 462760 4122
rect 462784 4066 462840 4122
rect 462864 4066 462920 4122
rect 462944 4066 463000 4122
rect 462704 2947 462760 3003
rect 462784 2947 462840 3003
rect 462864 2947 462920 3003
rect 462944 2947 463000 3003
rect 462704 2867 462760 2923
rect 462784 2867 462840 2923
rect 462864 2867 462920 2923
rect 462944 2867 463000 2923
rect 462704 2787 462760 2843
rect 462784 2787 462840 2843
rect 462864 2787 462920 2843
rect 462944 2787 463000 2843
rect 462704 2746 462760 2763
rect 462784 2746 462840 2763
rect 462864 2746 462920 2763
rect 462944 2746 463000 2763
rect 462704 2707 462750 2746
rect 462750 2707 462760 2746
rect 462784 2707 462814 2746
rect 462814 2707 462826 2746
rect 462826 2707 462840 2746
rect 462864 2707 462878 2746
rect 462878 2707 462890 2746
rect 462890 2707 462920 2746
rect 462944 2707 462954 2746
rect 462954 2707 463000 2746
rect 462704 908 462760 964
rect 462784 908 462840 964
rect 462864 908 462920 964
rect 462944 908 463000 964
rect 462704 828 462760 884
rect 462784 828 462840 884
rect 462864 828 462920 884
rect 462944 828 463000 884
rect 462704 748 462760 804
rect 462784 748 462840 804
rect 462864 748 462920 804
rect 462944 748 463000 804
rect 462704 668 462760 724
rect 462784 668 462840 724
rect 462864 668 462920 724
rect 462944 668 463000 724
rect 406382 448 406438 504
rect 409694 484 409696 504
rect 409696 484 409748 504
rect 409748 484 409750 504
rect 409694 448 409750 484
rect 331436 8 331492 64
rect 331516 8 331572 64
rect 331596 8 331652 64
rect 331676 8 331732 64
rect 463364 9728 463420 9784
rect 463444 9728 463500 9784
rect 463524 9728 463580 9784
rect 463604 9728 463660 9784
rect 463364 9648 463420 9704
rect 463444 9648 463500 9704
rect 463524 9648 463580 9704
rect 463604 9648 463660 9704
rect 463364 9568 463420 9624
rect 463444 9568 463500 9624
rect 463524 9568 463580 9624
rect 463604 9568 463660 9624
rect 463364 9488 463420 9544
rect 463444 9488 463500 9544
rect 463524 9488 463580 9544
rect 463604 9488 463660 9544
rect 530688 9728 530744 9784
rect 530768 9728 530824 9784
rect 530848 9728 530904 9784
rect 530928 9728 530984 9784
rect 530688 9648 530744 9704
rect 530768 9648 530824 9704
rect 530848 9648 530904 9704
rect 530928 9648 530984 9704
rect 530688 9568 530744 9624
rect 530768 9568 530824 9624
rect 530848 9568 530904 9624
rect 530928 9568 530984 9624
rect 530688 9488 530744 9544
rect 530768 9488 530824 9544
rect 530848 9488 530904 9544
rect 530928 9488 530984 9544
rect 463364 7684 463420 7740
rect 463444 7684 463500 7740
rect 463524 7684 463580 7740
rect 463604 7684 463660 7740
rect 463364 7642 463420 7660
rect 463444 7642 463500 7660
rect 463524 7642 463580 7660
rect 463604 7642 463660 7660
rect 463364 7604 463410 7642
rect 463410 7604 463420 7642
rect 463444 7604 463474 7642
rect 463474 7604 463486 7642
rect 463486 7604 463500 7642
rect 463524 7604 463538 7642
rect 463538 7604 463550 7642
rect 463550 7604 463580 7642
rect 463604 7604 463614 7642
rect 463614 7604 463660 7642
rect 463364 7524 463420 7580
rect 463444 7524 463500 7580
rect 463524 7524 463580 7580
rect 463604 7524 463660 7580
rect 463364 7444 463420 7500
rect 463444 7444 463500 7500
rect 463524 7444 463580 7500
rect 463604 7444 463660 7500
rect 463364 6325 463420 6381
rect 463444 6325 463500 6381
rect 463524 6325 463580 6381
rect 463604 6325 463660 6381
rect 463364 6245 463420 6301
rect 463444 6245 463500 6301
rect 463524 6245 463580 6301
rect 463604 6245 463660 6301
rect 463364 6165 463420 6221
rect 463444 6165 463500 6221
rect 463524 6165 463580 6221
rect 463604 6165 463660 6221
rect 530028 9068 530084 9124
rect 530108 9068 530164 9124
rect 530188 9068 530244 9124
rect 530268 9068 530324 9124
rect 530028 8988 530084 9044
rect 530108 8988 530164 9044
rect 530188 8988 530244 9044
rect 530268 8988 530324 9044
rect 530028 8908 530084 8964
rect 530108 8908 530164 8964
rect 530188 8908 530244 8964
rect 530268 8908 530324 8964
rect 530028 8828 530084 8884
rect 530108 8828 530164 8884
rect 530188 8828 530244 8884
rect 530268 8828 530324 8884
rect 530028 7024 530084 7080
rect 530108 7024 530164 7080
rect 530188 7024 530244 7080
rect 530268 7024 530324 7080
rect 530028 6944 530084 7000
rect 530108 6944 530164 7000
rect 530188 6944 530244 7000
rect 530268 6944 530324 7000
rect 530028 6864 530084 6920
rect 530108 6864 530164 6920
rect 530188 6864 530244 6920
rect 530268 6864 530324 6920
rect 530028 6784 530084 6840
rect 530108 6784 530164 6840
rect 530188 6784 530244 6840
rect 530268 6784 530324 6840
rect 463364 6085 463420 6141
rect 463444 6085 463500 6141
rect 463524 6085 463580 6141
rect 463604 6085 463660 6141
rect 463364 4966 463420 5022
rect 463444 4966 463500 5022
rect 463524 4966 463580 5022
rect 463604 4966 463660 5022
rect 463364 4886 463420 4942
rect 463444 4886 463500 4942
rect 463524 4886 463580 4942
rect 463604 4886 463660 4942
rect 463364 4806 463420 4862
rect 463444 4806 463500 4862
rect 463524 4806 463580 4862
rect 463604 4806 463660 4862
rect 463364 4726 463420 4782
rect 463444 4726 463500 4782
rect 463524 4726 463580 4782
rect 463604 4726 463660 4782
rect 463364 3607 463420 3663
rect 463444 3607 463500 3663
rect 463524 3607 463580 3663
rect 463604 3607 463660 3663
rect 463364 3527 463420 3583
rect 463444 3527 463500 3583
rect 463524 3527 463580 3583
rect 463604 3527 463660 3583
rect 463364 3447 463420 3503
rect 463444 3447 463500 3503
rect 463524 3447 463580 3503
rect 463604 3447 463660 3503
rect 463364 3367 463420 3423
rect 463444 3367 463500 3423
rect 463524 3367 463580 3423
rect 463604 3367 463660 3423
rect 530028 5665 530084 5721
rect 530108 5665 530164 5721
rect 530188 5665 530244 5721
rect 530268 5665 530324 5721
rect 530028 5585 530084 5641
rect 530108 5585 530164 5641
rect 530188 5585 530244 5641
rect 530268 5585 530324 5641
rect 530028 5505 530084 5561
rect 530108 5505 530164 5561
rect 530188 5505 530244 5561
rect 530268 5505 530324 5561
rect 530028 5425 530084 5481
rect 530108 5425 530164 5481
rect 530188 5425 530244 5481
rect 530268 5425 530324 5481
rect 530028 4306 530084 4362
rect 530108 4306 530164 4362
rect 530188 4306 530244 4362
rect 530268 4306 530324 4362
rect 530028 4226 530084 4282
rect 530108 4226 530164 4282
rect 530188 4226 530244 4282
rect 530268 4226 530324 4282
rect 465722 2388 465724 2408
rect 465724 2388 465776 2408
rect 465776 2388 465778 2408
rect 465722 2352 465778 2388
rect 463364 248 463420 304
rect 463444 248 463500 304
rect 463524 248 463580 304
rect 463604 248 463660 304
rect 463364 168 463420 224
rect 463444 168 463500 224
rect 463524 168 463580 224
rect 463604 168 463660 224
rect 463364 88 463420 144
rect 463444 88 463500 144
rect 463524 88 463580 144
rect 463604 88 463660 144
rect 530028 4146 530084 4202
rect 530108 4146 530164 4202
rect 530188 4146 530244 4202
rect 530268 4146 530324 4202
rect 530028 4066 530084 4122
rect 530108 4066 530164 4122
rect 530188 4066 530244 4122
rect 530268 4066 530324 4122
rect 530028 2947 530084 3003
rect 530108 2947 530164 3003
rect 530188 2947 530244 3003
rect 530268 2947 530324 3003
rect 530028 2867 530084 2923
rect 530108 2867 530164 2923
rect 530188 2867 530244 2923
rect 530268 2867 530324 2923
rect 530028 2787 530084 2843
rect 530108 2787 530164 2843
rect 530188 2787 530244 2843
rect 530268 2787 530324 2843
rect 530028 2707 530084 2763
rect 530108 2707 530164 2763
rect 530188 2707 530244 2763
rect 530268 2707 530324 2763
rect 530028 908 530084 964
rect 530108 908 530164 964
rect 530188 908 530244 964
rect 530268 908 530324 964
rect 530028 828 530084 884
rect 530108 828 530164 884
rect 530188 828 530244 884
rect 530268 828 530324 884
rect 530028 748 530084 804
rect 530108 748 530164 804
rect 530188 748 530244 804
rect 530268 748 530324 804
rect 530028 668 530084 724
rect 530108 668 530164 724
rect 530188 668 530244 724
rect 530268 668 530324 724
rect 530688 7684 530744 7740
rect 530768 7684 530824 7740
rect 530848 7684 530904 7740
rect 530928 7684 530984 7740
rect 530688 7604 530744 7660
rect 530768 7604 530824 7660
rect 530848 7604 530904 7660
rect 530928 7604 530984 7660
rect 530688 7524 530744 7580
rect 530768 7524 530824 7580
rect 530848 7524 530904 7580
rect 530928 7524 530984 7580
rect 530688 7444 530744 7500
rect 530768 7444 530824 7500
rect 530848 7444 530904 7500
rect 530928 7444 530984 7500
rect 530688 6325 530744 6381
rect 530768 6325 530824 6381
rect 530848 6325 530904 6381
rect 530928 6325 530984 6381
rect 530688 6245 530744 6301
rect 530768 6245 530824 6301
rect 530848 6245 530904 6301
rect 530928 6245 530984 6301
rect 530688 6165 530744 6221
rect 530768 6165 530824 6221
rect 530848 6165 530904 6221
rect 530928 6165 530984 6221
rect 530688 6085 530744 6141
rect 530768 6085 530824 6141
rect 530848 6085 530904 6141
rect 530928 6085 530984 6141
rect 530688 4966 530744 5022
rect 530768 4966 530824 5022
rect 530848 4966 530904 5022
rect 530928 4966 530984 5022
rect 530688 4886 530744 4942
rect 530768 4886 530824 4942
rect 530848 4886 530904 4942
rect 530928 4886 530984 4942
rect 530688 4806 530744 4862
rect 530768 4806 530824 4862
rect 530848 4806 530904 4862
rect 530928 4806 530984 4862
rect 530688 4726 530744 4782
rect 530768 4726 530824 4782
rect 530848 4726 530904 4782
rect 530928 4726 530984 4782
rect 530688 3607 530744 3663
rect 530768 3607 530824 3663
rect 530848 3607 530904 3663
rect 530928 3607 530984 3663
rect 530688 3527 530744 3583
rect 530768 3527 530824 3583
rect 530848 3527 530904 3583
rect 530928 3527 530984 3583
rect 530688 3447 530744 3503
rect 530768 3447 530824 3503
rect 530848 3447 530904 3503
rect 530928 3447 530984 3503
rect 530688 3367 530744 3423
rect 530768 3367 530824 3423
rect 530848 3367 530904 3423
rect 530928 3367 530984 3423
rect 479706 448 479762 504
rect 482650 448 482706 504
rect 530688 248 530744 304
rect 530768 248 530824 304
rect 530848 248 530904 304
rect 530928 248 530984 304
rect 530688 168 530744 224
rect 530768 168 530824 224
rect 530848 168 530904 224
rect 530928 168 530984 224
rect 530688 88 530744 144
rect 530768 88 530824 144
rect 530848 88 530904 144
rect 530928 88 530984 144
rect 463364 8 463420 64
rect 463444 8 463500 64
rect 463524 8 463580 64
rect 463604 8 463660 64
rect 530688 8 530744 64
rect 530768 8 530824 64
rect 530848 8 530904 64
rect 530928 8 530984 64
<< metal3 >>
rect -1076 9784 530996 9796
rect -1076 9728 -1064 9784
rect -1008 9728 -984 9784
rect -928 9728 -904 9784
rect -848 9728 -824 9784
rect -768 9728 67580 9784
rect 67636 9728 67660 9784
rect 67716 9728 67740 9784
rect 67796 9728 67820 9784
rect 67876 9728 199508 9784
rect 199564 9728 199588 9784
rect 199644 9728 199668 9784
rect 199724 9728 199748 9784
rect 199804 9728 331436 9784
rect 331492 9728 331516 9784
rect 331572 9728 331596 9784
rect 331652 9728 331676 9784
rect 331732 9728 463364 9784
rect 463420 9728 463444 9784
rect 463500 9728 463524 9784
rect 463580 9728 463604 9784
rect 463660 9728 530688 9784
rect 530744 9728 530768 9784
rect 530824 9728 530848 9784
rect 530904 9728 530928 9784
rect 530984 9728 530996 9784
rect -1076 9704 530996 9728
rect -1076 9648 -1064 9704
rect -1008 9648 -984 9704
rect -928 9648 -904 9704
rect -848 9648 -824 9704
rect -768 9648 67580 9704
rect 67636 9648 67660 9704
rect 67716 9648 67740 9704
rect 67796 9648 67820 9704
rect 67876 9648 199508 9704
rect 199564 9648 199588 9704
rect 199644 9648 199668 9704
rect 199724 9648 199748 9704
rect 199804 9648 331436 9704
rect 331492 9648 331516 9704
rect 331572 9648 331596 9704
rect 331652 9648 331676 9704
rect 331732 9648 463364 9704
rect 463420 9648 463444 9704
rect 463500 9648 463524 9704
rect 463580 9648 463604 9704
rect 463660 9648 530688 9704
rect 530744 9648 530768 9704
rect 530824 9648 530848 9704
rect 530904 9648 530928 9704
rect 530984 9648 530996 9704
rect -1076 9624 530996 9648
rect -1076 9568 -1064 9624
rect -1008 9568 -984 9624
rect -928 9568 -904 9624
rect -848 9568 -824 9624
rect -768 9568 67580 9624
rect 67636 9568 67660 9624
rect 67716 9568 67740 9624
rect 67796 9568 67820 9624
rect 67876 9568 199508 9624
rect 199564 9568 199588 9624
rect 199644 9568 199668 9624
rect 199724 9568 199748 9624
rect 199804 9568 331436 9624
rect 331492 9568 331516 9624
rect 331572 9568 331596 9624
rect 331652 9568 331676 9624
rect 331732 9568 463364 9624
rect 463420 9568 463444 9624
rect 463500 9568 463524 9624
rect 463580 9568 463604 9624
rect 463660 9568 530688 9624
rect 530744 9568 530768 9624
rect 530824 9568 530848 9624
rect 530904 9568 530928 9624
rect 530984 9568 530996 9624
rect -1076 9544 530996 9568
rect -1076 9488 -1064 9544
rect -1008 9488 -984 9544
rect -928 9488 -904 9544
rect -848 9488 -824 9544
rect -768 9488 67580 9544
rect 67636 9488 67660 9544
rect 67716 9488 67740 9544
rect 67796 9488 67820 9544
rect 67876 9488 199508 9544
rect 199564 9488 199588 9544
rect 199644 9488 199668 9544
rect 199724 9488 199748 9544
rect 199804 9488 331436 9544
rect 331492 9488 331516 9544
rect 331572 9488 331596 9544
rect 331652 9488 331676 9544
rect 331732 9488 463364 9544
rect 463420 9488 463444 9544
rect 463500 9488 463524 9544
rect 463580 9488 463604 9544
rect 463660 9488 530688 9544
rect 530744 9488 530768 9544
rect 530824 9488 530848 9544
rect 530904 9488 530928 9544
rect 530984 9488 530996 9544
rect -1076 9476 530996 9488
rect -416 9124 530336 9136
rect -416 9068 -404 9124
rect -348 9068 -324 9124
rect -268 9068 -244 9124
rect -188 9068 -164 9124
rect -108 9068 66920 9124
rect 66976 9068 67000 9124
rect 67056 9068 67080 9124
rect 67136 9068 67160 9124
rect 67216 9068 198848 9124
rect 198904 9068 198928 9124
rect 198984 9068 199008 9124
rect 199064 9068 199088 9124
rect 199144 9068 330776 9124
rect 330832 9068 330856 9124
rect 330912 9068 330936 9124
rect 330992 9068 331016 9124
rect 331072 9068 462704 9124
rect 462760 9068 462784 9124
rect 462840 9068 462864 9124
rect 462920 9068 462944 9124
rect 463000 9068 530028 9124
rect 530084 9068 530108 9124
rect 530164 9068 530188 9124
rect 530244 9068 530268 9124
rect 530324 9068 530336 9124
rect -416 9044 530336 9068
rect -416 8988 -404 9044
rect -348 8988 -324 9044
rect -268 8988 -244 9044
rect -188 8988 -164 9044
rect -108 8988 66920 9044
rect 66976 8988 67000 9044
rect 67056 8988 67080 9044
rect 67136 8988 67160 9044
rect 67216 8988 198848 9044
rect 198904 8988 198928 9044
rect 198984 8988 199008 9044
rect 199064 8988 199088 9044
rect 199144 8988 330776 9044
rect 330832 8988 330856 9044
rect 330912 8988 330936 9044
rect 330992 8988 331016 9044
rect 331072 8988 462704 9044
rect 462760 8988 462784 9044
rect 462840 8988 462864 9044
rect 462920 8988 462944 9044
rect 463000 8988 530028 9044
rect 530084 8988 530108 9044
rect 530164 8988 530188 9044
rect 530244 8988 530268 9044
rect 530324 8988 530336 9044
rect -416 8964 530336 8988
rect -416 8908 -404 8964
rect -348 8908 -324 8964
rect -268 8908 -244 8964
rect -188 8908 -164 8964
rect -108 8908 66920 8964
rect 66976 8908 67000 8964
rect 67056 8908 67080 8964
rect 67136 8908 67160 8964
rect 67216 8908 198848 8964
rect 198904 8908 198928 8964
rect 198984 8908 199008 8964
rect 199064 8908 199088 8964
rect 199144 8908 330776 8964
rect 330832 8908 330856 8964
rect 330912 8908 330936 8964
rect 330992 8908 331016 8964
rect 331072 8908 462704 8964
rect 462760 8908 462784 8964
rect 462840 8908 462864 8964
rect 462920 8908 462944 8964
rect 463000 8908 530028 8964
rect 530084 8908 530108 8964
rect 530164 8908 530188 8964
rect 530244 8908 530268 8964
rect 530324 8908 530336 8964
rect -416 8884 530336 8908
rect -416 8828 -404 8884
rect -348 8828 -324 8884
rect -268 8828 -244 8884
rect -188 8828 -164 8884
rect -108 8828 66920 8884
rect 66976 8828 67000 8884
rect 67056 8828 67080 8884
rect 67136 8828 67160 8884
rect 67216 8828 198848 8884
rect 198904 8828 198928 8884
rect 198984 8828 199008 8884
rect 199064 8828 199088 8884
rect 199144 8828 330776 8884
rect 330832 8828 330856 8884
rect 330912 8828 330936 8884
rect 330992 8828 331016 8884
rect 331072 8828 462704 8884
rect 462760 8828 462784 8884
rect 462840 8828 462864 8884
rect 462920 8828 462944 8884
rect 463000 8828 530028 8884
rect 530084 8828 530108 8884
rect 530164 8828 530188 8884
rect 530244 8828 530268 8884
rect 530324 8828 530336 8884
rect -416 8816 530336 8828
rect -1076 7740 530996 7752
rect -1076 7684 -1064 7740
rect -1008 7684 -984 7740
rect -928 7684 -904 7740
rect -848 7684 -824 7740
rect -768 7684 67580 7740
rect 67636 7684 67660 7740
rect 67716 7684 67740 7740
rect 67796 7684 67820 7740
rect 67876 7684 199508 7740
rect 199564 7684 199588 7740
rect 199644 7684 199668 7740
rect 199724 7684 199748 7740
rect 199804 7684 331436 7740
rect 331492 7684 331516 7740
rect 331572 7684 331596 7740
rect 331652 7684 331676 7740
rect 331732 7684 463364 7740
rect 463420 7684 463444 7740
rect 463500 7684 463524 7740
rect 463580 7684 463604 7740
rect 463660 7684 530688 7740
rect 530744 7684 530768 7740
rect 530824 7684 530848 7740
rect 530904 7684 530928 7740
rect 530984 7684 530996 7740
rect -1076 7660 530996 7684
rect -1076 7604 -1064 7660
rect -1008 7604 -984 7660
rect -928 7604 -904 7660
rect -848 7604 -824 7660
rect -768 7604 67580 7660
rect 67636 7604 67660 7660
rect 67716 7604 67740 7660
rect 67796 7604 67820 7660
rect 67876 7604 199508 7660
rect 199564 7604 199588 7660
rect 199644 7604 199668 7660
rect 199724 7604 199748 7660
rect 199804 7604 331436 7660
rect 331492 7604 331516 7660
rect 331572 7604 331596 7660
rect 331652 7604 331676 7660
rect 331732 7604 463364 7660
rect 463420 7604 463444 7660
rect 463500 7604 463524 7660
rect 463580 7604 463604 7660
rect 463660 7604 530688 7660
rect 530744 7604 530768 7660
rect 530824 7604 530848 7660
rect 530904 7604 530928 7660
rect 530984 7604 530996 7660
rect -1076 7580 530996 7604
rect -1076 7524 -1064 7580
rect -1008 7524 -984 7580
rect -928 7524 -904 7580
rect -848 7524 -824 7580
rect -768 7524 67580 7580
rect 67636 7524 67660 7580
rect 67716 7524 67740 7580
rect 67796 7524 67820 7580
rect 67876 7524 199508 7580
rect 199564 7524 199588 7580
rect 199644 7524 199668 7580
rect 199724 7524 199748 7580
rect 199804 7524 331436 7580
rect 331492 7524 331516 7580
rect 331572 7524 331596 7580
rect 331652 7524 331676 7580
rect 331732 7524 463364 7580
rect 463420 7524 463444 7580
rect 463500 7524 463524 7580
rect 463580 7524 463604 7580
rect 463660 7524 530688 7580
rect 530744 7524 530768 7580
rect 530824 7524 530848 7580
rect 530904 7524 530928 7580
rect 530984 7524 530996 7580
rect -1076 7500 530996 7524
rect -1076 7444 -1064 7500
rect -1008 7444 -984 7500
rect -928 7444 -904 7500
rect -848 7444 -824 7500
rect -768 7444 67580 7500
rect 67636 7444 67660 7500
rect 67716 7444 67740 7500
rect 67796 7444 67820 7500
rect 67876 7444 199508 7500
rect 199564 7444 199588 7500
rect 199644 7444 199668 7500
rect 199724 7444 199748 7500
rect 199804 7444 331436 7500
rect 331492 7444 331516 7500
rect 331572 7444 331596 7500
rect 331652 7444 331676 7500
rect 331732 7444 463364 7500
rect 463420 7444 463444 7500
rect 463500 7444 463524 7500
rect 463580 7444 463604 7500
rect 463660 7444 530688 7500
rect 530744 7444 530768 7500
rect 530824 7444 530848 7500
rect 530904 7444 530928 7500
rect 530984 7444 530996 7500
rect -1076 7432 530996 7444
rect -1076 7080 530996 7092
rect -1076 7024 -404 7080
rect -348 7024 -324 7080
rect -268 7024 -244 7080
rect -188 7024 -164 7080
rect -108 7024 66920 7080
rect 66976 7024 67000 7080
rect 67056 7024 67080 7080
rect 67136 7024 67160 7080
rect 67216 7024 198848 7080
rect 198904 7024 198928 7080
rect 198984 7024 199008 7080
rect 199064 7024 199088 7080
rect 199144 7024 330776 7080
rect 330832 7024 330856 7080
rect 330912 7024 330936 7080
rect 330992 7024 331016 7080
rect 331072 7024 462704 7080
rect 462760 7024 462784 7080
rect 462840 7024 462864 7080
rect 462920 7024 462944 7080
rect 463000 7024 530028 7080
rect 530084 7024 530108 7080
rect 530164 7024 530188 7080
rect 530244 7024 530268 7080
rect 530324 7024 530996 7080
rect -1076 7000 530996 7024
rect -1076 6944 -404 7000
rect -348 6944 -324 7000
rect -268 6944 -244 7000
rect -188 6944 -164 7000
rect -108 6944 66920 7000
rect 66976 6944 67000 7000
rect 67056 6944 67080 7000
rect 67136 6944 67160 7000
rect 67216 6944 198848 7000
rect 198904 6944 198928 7000
rect 198984 6944 199008 7000
rect 199064 6944 199088 7000
rect 199144 6944 330776 7000
rect 330832 6944 330856 7000
rect 330912 6944 330936 7000
rect 330992 6944 331016 7000
rect 331072 6944 462704 7000
rect 462760 6944 462784 7000
rect 462840 6944 462864 7000
rect 462920 6944 462944 7000
rect 463000 6944 530028 7000
rect 530084 6944 530108 7000
rect 530164 6944 530188 7000
rect 530244 6944 530268 7000
rect 530324 6944 530996 7000
rect -1076 6920 530996 6944
rect -1076 6864 -404 6920
rect -348 6864 -324 6920
rect -268 6864 -244 6920
rect -188 6864 -164 6920
rect -108 6864 66920 6920
rect 66976 6864 67000 6920
rect 67056 6864 67080 6920
rect 67136 6864 67160 6920
rect 67216 6864 198848 6920
rect 198904 6864 198928 6920
rect 198984 6864 199008 6920
rect 199064 6864 199088 6920
rect 199144 6864 330776 6920
rect 330832 6864 330856 6920
rect 330912 6864 330936 6920
rect 330992 6864 331016 6920
rect 331072 6864 462704 6920
rect 462760 6864 462784 6920
rect 462840 6864 462864 6920
rect 462920 6864 462944 6920
rect 463000 6864 530028 6920
rect 530084 6864 530108 6920
rect 530164 6864 530188 6920
rect 530244 6864 530268 6920
rect 530324 6864 530996 6920
rect -1076 6840 530996 6864
rect -1076 6784 -404 6840
rect -348 6784 -324 6840
rect -268 6784 -244 6840
rect -188 6784 -164 6840
rect -108 6784 66920 6840
rect 66976 6784 67000 6840
rect 67056 6784 67080 6840
rect 67136 6784 67160 6840
rect 67216 6784 198848 6840
rect 198904 6784 198928 6840
rect 198984 6784 199008 6840
rect 199064 6784 199088 6840
rect 199144 6784 330776 6840
rect 330832 6784 330856 6840
rect 330912 6784 330936 6840
rect 330992 6784 331016 6840
rect 331072 6784 462704 6840
rect 462760 6784 462784 6840
rect 462840 6784 462864 6840
rect 462920 6784 462944 6840
rect 463000 6784 530028 6840
rect 530084 6784 530108 6840
rect 530164 6784 530188 6840
rect 530244 6784 530268 6840
rect 530324 6784 530996 6840
rect -1076 6772 530996 6784
rect -1076 6381 530996 6393
rect -1076 6325 -1064 6381
rect -1008 6325 -984 6381
rect -928 6325 -904 6381
rect -848 6325 -824 6381
rect -768 6325 67580 6381
rect 67636 6325 67660 6381
rect 67716 6325 67740 6381
rect 67796 6325 67820 6381
rect 67876 6325 199508 6381
rect 199564 6325 199588 6381
rect 199644 6325 199668 6381
rect 199724 6325 199748 6381
rect 199804 6325 331436 6381
rect 331492 6325 331516 6381
rect 331572 6325 331596 6381
rect 331652 6325 331676 6381
rect 331732 6325 463364 6381
rect 463420 6325 463444 6381
rect 463500 6325 463524 6381
rect 463580 6325 463604 6381
rect 463660 6325 530688 6381
rect 530744 6325 530768 6381
rect 530824 6325 530848 6381
rect 530904 6325 530928 6381
rect 530984 6325 530996 6381
rect -1076 6301 530996 6325
rect -1076 6245 -1064 6301
rect -1008 6245 -984 6301
rect -928 6245 -904 6301
rect -848 6245 -824 6301
rect -768 6245 67580 6301
rect 67636 6245 67660 6301
rect 67716 6245 67740 6301
rect 67796 6245 67820 6301
rect 67876 6245 199508 6301
rect 199564 6245 199588 6301
rect 199644 6245 199668 6301
rect 199724 6245 199748 6301
rect 199804 6245 331436 6301
rect 331492 6245 331516 6301
rect 331572 6245 331596 6301
rect 331652 6245 331676 6301
rect 331732 6245 463364 6301
rect 463420 6245 463444 6301
rect 463500 6245 463524 6301
rect 463580 6245 463604 6301
rect 463660 6245 530688 6301
rect 530744 6245 530768 6301
rect 530824 6245 530848 6301
rect 530904 6245 530928 6301
rect 530984 6245 530996 6301
rect -1076 6221 530996 6245
rect -1076 6165 -1064 6221
rect -1008 6165 -984 6221
rect -928 6165 -904 6221
rect -848 6165 -824 6221
rect -768 6165 67580 6221
rect 67636 6165 67660 6221
rect 67716 6165 67740 6221
rect 67796 6165 67820 6221
rect 67876 6165 199508 6221
rect 199564 6165 199588 6221
rect 199644 6165 199668 6221
rect 199724 6165 199748 6221
rect 199804 6165 331436 6221
rect 331492 6165 331516 6221
rect 331572 6165 331596 6221
rect 331652 6165 331676 6221
rect 331732 6165 463364 6221
rect 463420 6165 463444 6221
rect 463500 6165 463524 6221
rect 463580 6165 463604 6221
rect 463660 6165 530688 6221
rect 530744 6165 530768 6221
rect 530824 6165 530848 6221
rect 530904 6165 530928 6221
rect 530984 6165 530996 6221
rect -1076 6141 530996 6165
rect -1076 6085 -1064 6141
rect -1008 6085 -984 6141
rect -928 6085 -904 6141
rect -848 6085 -824 6141
rect -768 6085 67580 6141
rect 67636 6085 67660 6141
rect 67716 6085 67740 6141
rect 67796 6085 67820 6141
rect 67876 6085 199508 6141
rect 199564 6085 199588 6141
rect 199644 6085 199668 6141
rect 199724 6085 199748 6141
rect 199804 6085 331436 6141
rect 331492 6085 331516 6141
rect 331572 6085 331596 6141
rect 331652 6085 331676 6141
rect 331732 6085 463364 6141
rect 463420 6085 463444 6141
rect 463500 6085 463524 6141
rect 463580 6085 463604 6141
rect 463660 6085 530688 6141
rect 530744 6085 530768 6141
rect 530824 6085 530848 6141
rect 530904 6085 530928 6141
rect 530984 6085 530996 6141
rect -1076 6073 530996 6085
rect -1076 5721 530996 5733
rect -1076 5665 -404 5721
rect -348 5665 -324 5721
rect -268 5665 -244 5721
rect -188 5665 -164 5721
rect -108 5665 66920 5721
rect 66976 5665 67000 5721
rect 67056 5665 67080 5721
rect 67136 5665 67160 5721
rect 67216 5665 198848 5721
rect 198904 5665 198928 5721
rect 198984 5665 199008 5721
rect 199064 5665 199088 5721
rect 199144 5665 330776 5721
rect 330832 5665 330856 5721
rect 330912 5665 330936 5721
rect 330992 5665 331016 5721
rect 331072 5665 462704 5721
rect 462760 5665 462784 5721
rect 462840 5665 462864 5721
rect 462920 5665 462944 5721
rect 463000 5665 530028 5721
rect 530084 5665 530108 5721
rect 530164 5665 530188 5721
rect 530244 5665 530268 5721
rect 530324 5665 530996 5721
rect -1076 5641 530996 5665
rect -1076 5585 -404 5641
rect -348 5585 -324 5641
rect -268 5585 -244 5641
rect -188 5585 -164 5641
rect -108 5585 66920 5641
rect 66976 5585 67000 5641
rect 67056 5585 67080 5641
rect 67136 5585 67160 5641
rect 67216 5585 198848 5641
rect 198904 5585 198928 5641
rect 198984 5585 199008 5641
rect 199064 5585 199088 5641
rect 199144 5585 330776 5641
rect 330832 5585 330856 5641
rect 330912 5585 330936 5641
rect 330992 5585 331016 5641
rect 331072 5585 462704 5641
rect 462760 5585 462784 5641
rect 462840 5585 462864 5641
rect 462920 5585 462944 5641
rect 463000 5585 530028 5641
rect 530084 5585 530108 5641
rect 530164 5585 530188 5641
rect 530244 5585 530268 5641
rect 530324 5585 530996 5641
rect -1076 5561 530996 5585
rect -1076 5505 -404 5561
rect -348 5505 -324 5561
rect -268 5505 -244 5561
rect -188 5505 -164 5561
rect -108 5505 66920 5561
rect 66976 5505 67000 5561
rect 67056 5505 67080 5561
rect 67136 5505 67160 5561
rect 67216 5505 198848 5561
rect 198904 5505 198928 5561
rect 198984 5505 199008 5561
rect 199064 5505 199088 5561
rect 199144 5505 330776 5561
rect 330832 5505 330856 5561
rect 330912 5505 330936 5561
rect 330992 5505 331016 5561
rect 331072 5505 462704 5561
rect 462760 5505 462784 5561
rect 462840 5505 462864 5561
rect 462920 5505 462944 5561
rect 463000 5505 530028 5561
rect 530084 5505 530108 5561
rect 530164 5505 530188 5561
rect 530244 5505 530268 5561
rect 530324 5505 530996 5561
rect -1076 5481 530996 5505
rect -1076 5425 -404 5481
rect -348 5425 -324 5481
rect -268 5425 -244 5481
rect -188 5425 -164 5481
rect -108 5425 66920 5481
rect 66976 5425 67000 5481
rect 67056 5425 67080 5481
rect 67136 5425 67160 5481
rect 67216 5425 198848 5481
rect 198904 5425 198928 5481
rect 198984 5425 199008 5481
rect 199064 5425 199088 5481
rect 199144 5425 330776 5481
rect 330832 5425 330856 5481
rect 330912 5425 330936 5481
rect 330992 5425 331016 5481
rect 331072 5425 462704 5481
rect 462760 5425 462784 5481
rect 462840 5425 462864 5481
rect 462920 5425 462944 5481
rect 463000 5425 530028 5481
rect 530084 5425 530108 5481
rect 530164 5425 530188 5481
rect 530244 5425 530268 5481
rect 530324 5425 530996 5481
rect -1076 5413 530996 5425
rect -1076 5022 530996 5034
rect -1076 4966 -1064 5022
rect -1008 4966 -984 5022
rect -928 4966 -904 5022
rect -848 4966 -824 5022
rect -768 4966 67580 5022
rect 67636 4966 67660 5022
rect 67716 4966 67740 5022
rect 67796 4966 67820 5022
rect 67876 4966 199508 5022
rect 199564 4966 199588 5022
rect 199644 4966 199668 5022
rect 199724 4966 199748 5022
rect 199804 4966 331436 5022
rect 331492 4966 331516 5022
rect 331572 4966 331596 5022
rect 331652 4966 331676 5022
rect 331732 4966 463364 5022
rect 463420 4966 463444 5022
rect 463500 4966 463524 5022
rect 463580 4966 463604 5022
rect 463660 4966 530688 5022
rect 530744 4966 530768 5022
rect 530824 4966 530848 5022
rect 530904 4966 530928 5022
rect 530984 4966 530996 5022
rect -1076 4942 530996 4966
rect -1076 4886 -1064 4942
rect -1008 4886 -984 4942
rect -928 4886 -904 4942
rect -848 4886 -824 4942
rect -768 4886 67580 4942
rect 67636 4886 67660 4942
rect 67716 4886 67740 4942
rect 67796 4886 67820 4942
rect 67876 4886 199508 4942
rect 199564 4886 199588 4942
rect 199644 4886 199668 4942
rect 199724 4886 199748 4942
rect 199804 4886 331436 4942
rect 331492 4886 331516 4942
rect 331572 4886 331596 4942
rect 331652 4886 331676 4942
rect 331732 4886 463364 4942
rect 463420 4886 463444 4942
rect 463500 4886 463524 4942
rect 463580 4886 463604 4942
rect 463660 4886 530688 4942
rect 530744 4886 530768 4942
rect 530824 4886 530848 4942
rect 530904 4886 530928 4942
rect 530984 4886 530996 4942
rect -1076 4862 530996 4886
rect -1076 4806 -1064 4862
rect -1008 4806 -984 4862
rect -928 4806 -904 4862
rect -848 4806 -824 4862
rect -768 4806 67580 4862
rect 67636 4806 67660 4862
rect 67716 4806 67740 4862
rect 67796 4806 67820 4862
rect 67876 4806 199508 4862
rect 199564 4806 199588 4862
rect 199644 4806 199668 4862
rect 199724 4806 199748 4862
rect 199804 4806 331436 4862
rect 331492 4806 331516 4862
rect 331572 4806 331596 4862
rect 331652 4806 331676 4862
rect 331732 4806 463364 4862
rect 463420 4806 463444 4862
rect 463500 4806 463524 4862
rect 463580 4806 463604 4862
rect 463660 4806 530688 4862
rect 530744 4806 530768 4862
rect 530824 4806 530848 4862
rect 530904 4806 530928 4862
rect 530984 4806 530996 4862
rect -1076 4782 530996 4806
rect -1076 4726 -1064 4782
rect -1008 4726 -984 4782
rect -928 4726 -904 4782
rect -848 4726 -824 4782
rect -768 4726 67580 4782
rect 67636 4726 67660 4782
rect 67716 4726 67740 4782
rect 67796 4726 67820 4782
rect 67876 4726 199508 4782
rect 199564 4726 199588 4782
rect 199644 4726 199668 4782
rect 199724 4726 199748 4782
rect 199804 4726 331436 4782
rect 331492 4726 331516 4782
rect 331572 4726 331596 4782
rect 331652 4726 331676 4782
rect 331732 4726 463364 4782
rect 463420 4726 463444 4782
rect 463500 4726 463524 4782
rect 463580 4726 463604 4782
rect 463660 4726 530688 4782
rect 530744 4726 530768 4782
rect 530824 4726 530848 4782
rect 530904 4726 530928 4782
rect 530984 4726 530996 4782
rect -1076 4714 530996 4726
rect -1076 4362 530996 4374
rect -1076 4306 -404 4362
rect -348 4306 -324 4362
rect -268 4306 -244 4362
rect -188 4306 -164 4362
rect -108 4306 66920 4362
rect 66976 4306 67000 4362
rect 67056 4306 67080 4362
rect 67136 4306 67160 4362
rect 67216 4306 198848 4362
rect 198904 4306 198928 4362
rect 198984 4306 199008 4362
rect 199064 4306 199088 4362
rect 199144 4306 330776 4362
rect 330832 4306 330856 4362
rect 330912 4306 330936 4362
rect 330992 4306 331016 4362
rect 331072 4306 462704 4362
rect 462760 4306 462784 4362
rect 462840 4306 462864 4362
rect 462920 4306 462944 4362
rect 463000 4306 530028 4362
rect 530084 4306 530108 4362
rect 530164 4306 530188 4362
rect 530244 4306 530268 4362
rect 530324 4306 530996 4362
rect -1076 4282 530996 4306
rect -1076 4226 -404 4282
rect -348 4226 -324 4282
rect -268 4226 -244 4282
rect -188 4226 -164 4282
rect -108 4226 66920 4282
rect 66976 4226 67000 4282
rect 67056 4226 67080 4282
rect 67136 4226 67160 4282
rect 67216 4226 198848 4282
rect 198904 4226 198928 4282
rect 198984 4226 199008 4282
rect 199064 4226 199088 4282
rect 199144 4226 330776 4282
rect 330832 4226 330856 4282
rect 330912 4226 330936 4282
rect 330992 4226 331016 4282
rect 331072 4226 462704 4282
rect 462760 4226 462784 4282
rect 462840 4226 462864 4282
rect 462920 4226 462944 4282
rect 463000 4226 530028 4282
rect 530084 4226 530108 4282
rect 530164 4226 530188 4282
rect 530244 4226 530268 4282
rect 530324 4226 530996 4282
rect -1076 4202 530996 4226
rect -1076 4146 -404 4202
rect -348 4146 -324 4202
rect -268 4146 -244 4202
rect -188 4146 -164 4202
rect -108 4146 66920 4202
rect 66976 4146 67000 4202
rect 67056 4146 67080 4202
rect 67136 4146 67160 4202
rect 67216 4146 198848 4202
rect 198904 4146 198928 4202
rect 198984 4146 199008 4202
rect 199064 4146 199088 4202
rect 199144 4146 330776 4202
rect 330832 4146 330856 4202
rect 330912 4146 330936 4202
rect 330992 4146 331016 4202
rect 331072 4146 462704 4202
rect 462760 4146 462784 4202
rect 462840 4146 462864 4202
rect 462920 4146 462944 4202
rect 463000 4146 530028 4202
rect 530084 4146 530108 4202
rect 530164 4146 530188 4202
rect 530244 4146 530268 4202
rect 530324 4146 530996 4202
rect -1076 4122 530996 4146
rect -1076 4066 -404 4122
rect -348 4066 -324 4122
rect -268 4066 -244 4122
rect -188 4066 -164 4122
rect -108 4066 66920 4122
rect 66976 4066 67000 4122
rect 67056 4066 67080 4122
rect 67136 4066 67160 4122
rect 67216 4066 198848 4122
rect 198904 4066 198928 4122
rect 198984 4066 199008 4122
rect 199064 4066 199088 4122
rect 199144 4066 330776 4122
rect 330832 4066 330856 4122
rect 330912 4066 330936 4122
rect 330992 4066 331016 4122
rect 331072 4066 462704 4122
rect 462760 4066 462784 4122
rect 462840 4066 462864 4122
rect 462920 4066 462944 4122
rect 463000 4066 530028 4122
rect 530084 4066 530108 4122
rect 530164 4066 530188 4122
rect 530244 4066 530268 4122
rect 530324 4066 530996 4122
rect -1076 4054 530996 4066
rect 214281 3906 214347 3909
rect 310881 3906 310947 3909
rect 214281 3904 310947 3906
rect 214281 3848 214286 3904
rect 214342 3848 310886 3904
rect 310942 3848 310947 3904
rect 214281 3846 310947 3848
rect 214281 3843 214347 3846
rect 310881 3843 310947 3846
rect -1076 3663 530996 3675
rect -1076 3607 -1064 3663
rect -1008 3607 -984 3663
rect -928 3607 -904 3663
rect -848 3607 -824 3663
rect -768 3607 67580 3663
rect 67636 3607 67660 3663
rect 67716 3607 67740 3663
rect 67796 3607 67820 3663
rect 67876 3607 199508 3663
rect 199564 3607 199588 3663
rect 199644 3607 199668 3663
rect 199724 3607 199748 3663
rect 199804 3607 331436 3663
rect 331492 3607 331516 3663
rect 331572 3607 331596 3663
rect 331652 3607 331676 3663
rect 331732 3607 463364 3663
rect 463420 3607 463444 3663
rect 463500 3607 463524 3663
rect 463580 3607 463604 3663
rect 463660 3607 530688 3663
rect 530744 3607 530768 3663
rect 530824 3607 530848 3663
rect 530904 3607 530928 3663
rect 530984 3607 530996 3663
rect -1076 3583 530996 3607
rect -1076 3527 -1064 3583
rect -1008 3527 -984 3583
rect -928 3527 -904 3583
rect -848 3527 -824 3583
rect -768 3527 67580 3583
rect 67636 3527 67660 3583
rect 67716 3527 67740 3583
rect 67796 3527 67820 3583
rect 67876 3527 199508 3583
rect 199564 3527 199588 3583
rect 199644 3527 199668 3583
rect 199724 3527 199748 3583
rect 199804 3527 331436 3583
rect 331492 3527 331516 3583
rect 331572 3527 331596 3583
rect 331652 3527 331676 3583
rect 331732 3527 463364 3583
rect 463420 3527 463444 3583
rect 463500 3527 463524 3583
rect 463580 3527 463604 3583
rect 463660 3527 530688 3583
rect 530744 3527 530768 3583
rect 530824 3527 530848 3583
rect 530904 3527 530928 3583
rect 530984 3527 530996 3583
rect -1076 3503 530996 3527
rect -1076 3447 -1064 3503
rect -1008 3447 -984 3503
rect -928 3447 -904 3503
rect -848 3447 -824 3503
rect -768 3447 67580 3503
rect 67636 3447 67660 3503
rect 67716 3447 67740 3503
rect 67796 3447 67820 3503
rect 67876 3447 199508 3503
rect 199564 3447 199588 3503
rect 199644 3447 199668 3503
rect 199724 3447 199748 3503
rect 199804 3447 331436 3503
rect 331492 3447 331516 3503
rect 331572 3447 331596 3503
rect 331652 3447 331676 3503
rect 331732 3447 463364 3503
rect 463420 3447 463444 3503
rect 463500 3447 463524 3503
rect 463580 3447 463604 3503
rect 463660 3447 530688 3503
rect 530744 3447 530768 3503
rect 530824 3447 530848 3503
rect 530904 3447 530928 3503
rect 530984 3447 530996 3503
rect -1076 3423 530996 3447
rect -1076 3367 -1064 3423
rect -1008 3367 -984 3423
rect -928 3367 -904 3423
rect -848 3367 -824 3423
rect -768 3367 67580 3423
rect 67636 3367 67660 3423
rect 67716 3367 67740 3423
rect 67796 3367 67820 3423
rect 67876 3367 199508 3423
rect 199564 3367 199588 3423
rect 199644 3367 199668 3423
rect 199724 3367 199748 3423
rect 199804 3367 331436 3423
rect 331492 3367 331516 3423
rect 331572 3367 331596 3423
rect 331652 3367 331676 3423
rect 331732 3367 463364 3423
rect 463420 3367 463444 3423
rect 463500 3367 463524 3423
rect 463580 3367 463604 3423
rect 463660 3367 530688 3423
rect 530744 3367 530768 3423
rect 530824 3367 530848 3423
rect 530904 3367 530928 3423
rect 530984 3367 530996 3423
rect -1076 3355 530996 3367
rect 122557 3226 122623 3229
rect 216673 3226 216739 3229
rect 122557 3224 216739 3226
rect 122557 3168 122562 3224
rect 122618 3168 216678 3224
rect 216734 3168 216739 3224
rect 122557 3166 216739 3168
rect 122557 3163 122623 3166
rect 216673 3163 216739 3166
rect -1076 3003 530996 3015
rect -1076 2947 -404 3003
rect -348 2947 -324 3003
rect -268 2947 -244 3003
rect -188 2947 -164 3003
rect -108 2947 66920 3003
rect 66976 2947 67000 3003
rect 67056 2947 67080 3003
rect 67136 2947 67160 3003
rect 67216 2947 198848 3003
rect 198904 2947 198928 3003
rect 198984 2947 199008 3003
rect 199064 2947 199088 3003
rect 199144 2947 330776 3003
rect 330832 2947 330856 3003
rect 330912 2947 330936 3003
rect 330992 2947 331016 3003
rect 331072 2947 462704 3003
rect 462760 2947 462784 3003
rect 462840 2947 462864 3003
rect 462920 2947 462944 3003
rect 463000 2947 530028 3003
rect 530084 2947 530108 3003
rect 530164 2947 530188 3003
rect 530244 2947 530268 3003
rect 530324 2947 530996 3003
rect -1076 2923 530996 2947
rect -1076 2867 -404 2923
rect -348 2867 -324 2923
rect -268 2867 -244 2923
rect -188 2867 -164 2923
rect -108 2867 66920 2923
rect 66976 2867 67000 2923
rect 67056 2867 67080 2923
rect 67136 2867 67160 2923
rect 67216 2867 198848 2923
rect 198904 2867 198928 2923
rect 198984 2867 199008 2923
rect 199064 2867 199088 2923
rect 199144 2867 330776 2923
rect 330832 2867 330856 2923
rect 330912 2867 330936 2923
rect 330992 2867 331016 2923
rect 331072 2867 462704 2923
rect 462760 2867 462784 2923
rect 462840 2867 462864 2923
rect 462920 2867 462944 2923
rect 463000 2867 530028 2923
rect 530084 2867 530108 2923
rect 530164 2867 530188 2923
rect 530244 2867 530268 2923
rect 530324 2867 530996 2923
rect -1076 2843 530996 2867
rect -1076 2787 -404 2843
rect -348 2787 -324 2843
rect -268 2787 -244 2843
rect -188 2787 -164 2843
rect -108 2787 66920 2843
rect 66976 2787 67000 2843
rect 67056 2787 67080 2843
rect 67136 2787 67160 2843
rect 67216 2787 198848 2843
rect 198904 2787 198928 2843
rect 198984 2787 199008 2843
rect 199064 2787 199088 2843
rect 199144 2787 330776 2843
rect 330832 2787 330856 2843
rect 330912 2787 330936 2843
rect 330992 2787 331016 2843
rect 331072 2787 462704 2843
rect 462760 2787 462784 2843
rect 462840 2787 462864 2843
rect 462920 2787 462944 2843
rect 463000 2787 530028 2843
rect 530084 2787 530108 2843
rect 530164 2787 530188 2843
rect 530244 2787 530268 2843
rect 530324 2787 530996 2843
rect -1076 2763 530996 2787
rect -1076 2707 -404 2763
rect -348 2707 -324 2763
rect -268 2707 -244 2763
rect -188 2707 -164 2763
rect -108 2707 66920 2763
rect 66976 2707 67000 2763
rect 67056 2707 67080 2763
rect 67136 2707 67160 2763
rect 67216 2707 198848 2763
rect 198904 2707 198928 2763
rect 198984 2707 199008 2763
rect 199064 2707 199088 2763
rect 199144 2707 330776 2763
rect 330832 2707 330856 2763
rect 330912 2707 330936 2763
rect 330992 2707 331016 2763
rect 331072 2707 462704 2763
rect 462760 2707 462784 2763
rect 462840 2707 462864 2763
rect 462920 2707 462944 2763
rect 463000 2707 530028 2763
rect 530084 2707 530108 2763
rect 530164 2707 530188 2763
rect 530244 2707 530268 2763
rect 530324 2707 530996 2763
rect -1076 2695 530996 2707
rect 54661 2546 54727 2549
rect 148225 2546 148291 2549
rect 54661 2544 148291 2546
rect 54661 2488 54666 2544
rect 54722 2488 148230 2544
rect 148286 2488 148291 2544
rect 54661 2486 148291 2488
rect 54661 2483 54727 2486
rect 148225 2483 148291 2486
rect 296989 2546 297055 2549
rect 391105 2546 391171 2549
rect 296989 2544 391171 2546
rect 296989 2488 296994 2544
rect 297050 2488 391110 2544
rect 391166 2488 391171 2544
rect 296989 2486 391171 2488
rect 296989 2483 297055 2486
rect 391105 2483 391171 2486
rect 396073 2546 396139 2549
rect 400765 2546 400831 2549
rect 396073 2544 400831 2546
rect 396073 2488 396078 2544
rect 396134 2488 400770 2544
rect 400826 2488 400831 2544
rect 396073 2486 400831 2488
rect 396073 2483 396139 2486
rect 400765 2483 400831 2486
rect 107653 2410 107719 2413
rect 201677 2410 201743 2413
rect 107653 2408 201743 2410
rect 107653 2352 107658 2408
rect 107714 2352 201682 2408
rect 201738 2352 201743 2408
rect 107653 2350 201743 2352
rect 107653 2347 107719 2350
rect 201677 2347 201743 2350
rect 213545 2410 213611 2413
rect 310697 2410 310763 2413
rect 213545 2408 310763 2410
rect 213545 2352 213550 2408
rect 213606 2352 310702 2408
rect 310758 2352 310763 2408
rect 213545 2350 310763 2352
rect 213545 2347 213611 2350
rect 310697 2347 310763 2350
rect 372429 2410 372495 2413
rect 465717 2410 465783 2413
rect 372429 2408 465783 2410
rect 372429 2352 372434 2408
rect 372490 2352 465722 2408
rect 465778 2352 465783 2408
rect 372429 2350 465783 2352
rect 372429 2347 372495 2350
rect 465717 2347 465783 2350
rect 122649 2274 122715 2277
rect 214005 2274 214071 2277
rect 122649 2272 214071 2274
rect 122649 2216 122654 2272
rect 122710 2216 214010 2272
rect 214066 2216 214071 2272
rect 122649 2214 214071 2216
rect 122649 2211 122715 2214
rect 214005 2211 214071 2214
rect 300761 2274 300827 2277
rect 394417 2274 394483 2277
rect 300761 2272 394483 2274
rect 300761 2216 300766 2272
rect 300822 2216 394422 2272
rect 394478 2216 394483 2272
rect 300761 2214 394483 2216
rect 300761 2211 300827 2214
rect 394417 2211 394483 2214
rect 123201 2138 123267 2141
rect 215385 2138 215451 2141
rect 123201 2136 215451 2138
rect 123201 2080 123206 2136
rect 123262 2080 215390 2136
rect 215446 2080 215451 2136
rect 123201 2078 215451 2080
rect 123201 2075 123267 2078
rect 215385 2075 215451 2078
rect 224217 2138 224283 2141
rect 317045 2138 317111 2141
rect 224217 2136 317111 2138
rect 224217 2080 224222 2136
rect 224278 2080 317050 2136
rect 317106 2080 317111 2136
rect 224217 2078 317111 2080
rect 224217 2075 224283 2078
rect 317045 2075 317111 2078
rect 355961 2138 356027 2141
rect 439405 2138 439471 2141
rect 355961 2136 439471 2138
rect 355961 2080 355966 2136
rect 356022 2080 439410 2136
rect 439466 2080 439471 2136
rect 355961 2078 439471 2080
rect 355961 2075 356027 2078
rect 439405 2075 439471 2078
rect 36721 2002 36787 2005
rect 130193 2002 130259 2005
rect 36721 2000 130259 2002
rect 36721 1944 36726 2000
rect 36782 1944 130198 2000
rect 130254 1944 130259 2000
rect 36721 1942 130259 1944
rect 36721 1939 36787 1942
rect 130193 1939 130259 1942
rect 260281 2002 260347 2005
rect 353293 2002 353359 2005
rect 260281 2000 353359 2002
rect 260281 1944 260286 2000
rect 260342 1944 353298 2000
rect 353354 1944 353359 2000
rect 260281 1942 353359 1944
rect 260281 1939 260347 1942
rect 353293 1939 353359 1942
rect 390553 2002 390619 2005
rect 435449 2002 435515 2005
rect 390553 2000 435515 2002
rect 390553 1944 390558 2000
rect 390614 1944 435454 2000
rect 435510 1944 435515 2000
rect 390553 1942 435515 1944
rect 390553 1939 390619 1942
rect 435449 1939 435515 1942
rect 29085 1866 29151 1869
rect 36537 1866 36603 1869
rect 29085 1864 36603 1866
rect 29085 1808 29090 1864
rect 29146 1808 36542 1864
rect 36598 1808 36603 1864
rect 29085 1806 36603 1808
rect 29085 1803 29151 1806
rect 36537 1803 36603 1806
rect 303981 1866 304047 1869
rect 396901 1866 396967 1869
rect 303981 1864 396967 1866
rect 303981 1808 303986 1864
rect 304042 1808 396906 1864
rect 396962 1808 396967 1864
rect 303981 1806 396967 1808
rect 303981 1803 304047 1806
rect 396901 1803 396967 1806
rect 31201 1730 31267 1733
rect 33777 1730 33843 1733
rect 31201 1728 33843 1730
rect 31201 1672 31206 1728
rect 31262 1672 33782 1728
rect 33838 1672 33843 1728
rect 31201 1670 33843 1672
rect 31201 1667 31267 1670
rect 33777 1667 33843 1670
rect 399477 1730 399543 1733
rect 408585 1730 408651 1733
rect 399477 1728 408651 1730
rect 399477 1672 399482 1728
rect 399538 1672 408590 1728
rect 408646 1672 408651 1728
rect 399477 1670 408651 1672
rect 399477 1667 399543 1670
rect 408585 1667 408651 1670
rect 26049 1594 26115 1597
rect 32857 1594 32923 1597
rect 26049 1592 32923 1594
rect 26049 1536 26054 1592
rect 26110 1536 32862 1592
rect 32918 1536 32923 1592
rect 26049 1534 32923 1536
rect 26049 1531 26115 1534
rect 32857 1531 32923 1534
rect 399293 1594 399359 1597
rect 402605 1594 402671 1597
rect 399293 1592 402671 1594
rect 399293 1536 399298 1592
rect 399354 1536 402610 1592
rect 402666 1536 402671 1592
rect 399293 1534 402671 1536
rect 399293 1531 399359 1534
rect 402605 1531 402671 1534
rect 26969 1458 27035 1461
rect 31845 1458 31911 1461
rect 26969 1456 31911 1458
rect 26969 1400 26974 1456
rect 27030 1400 31850 1456
rect 31906 1400 31911 1456
rect 26969 1398 31911 1400
rect 26969 1395 27035 1398
rect 31845 1395 31911 1398
rect 398005 1458 398071 1461
rect 399017 1458 399083 1461
rect 404813 1458 404879 1461
rect 398005 1456 399083 1458
rect 398005 1400 398010 1456
rect 398066 1400 399022 1456
rect 399078 1400 399083 1456
rect 398005 1398 399083 1400
rect 398005 1395 398071 1398
rect 399017 1395 399083 1398
rect 399158 1456 404879 1458
rect 399158 1400 404818 1456
rect 404874 1400 404879 1456
rect 399158 1398 404879 1400
rect 31201 1322 31267 1325
rect 31753 1322 31819 1325
rect 31201 1320 31819 1322
rect 31201 1264 31206 1320
rect 31262 1264 31758 1320
rect 31814 1264 31819 1320
rect 31201 1262 31819 1264
rect 31201 1259 31267 1262
rect 31753 1259 31819 1262
rect 398833 1322 398899 1325
rect 399158 1322 399218 1398
rect 404813 1395 404879 1398
rect 398833 1320 399218 1322
rect 398833 1264 398838 1320
rect 398894 1264 399218 1320
rect 398833 1262 399218 1264
rect 399661 1322 399727 1325
rect 404261 1322 404327 1325
rect 399661 1320 404327 1322
rect 399661 1264 399666 1320
rect 399722 1264 404266 1320
rect 404322 1264 404327 1320
rect 399661 1262 404327 1264
rect 398833 1259 398899 1262
rect 399661 1259 399727 1262
rect 404261 1259 404327 1262
rect 407481 1322 407547 1325
rect 410793 1322 410859 1325
rect 407481 1320 410859 1322
rect 407481 1264 407486 1320
rect 407542 1264 410798 1320
rect 410854 1264 410859 1320
rect 407481 1262 410859 1264
rect 407481 1259 407547 1262
rect 410793 1259 410859 1262
rect 28533 1186 28599 1189
rect 31569 1186 31635 1189
rect 28533 1184 31635 1186
rect 28533 1128 28538 1184
rect 28594 1128 31574 1184
rect 31630 1128 31635 1184
rect 28533 1126 31635 1128
rect 28533 1123 28599 1126
rect 31569 1123 31635 1126
rect 399845 1186 399911 1189
rect 407481 1186 407547 1189
rect 399845 1184 407547 1186
rect 399845 1128 399850 1184
rect 399906 1128 407486 1184
rect 407542 1128 407547 1184
rect 399845 1126 407547 1128
rect 399845 1123 399911 1126
rect 407481 1123 407547 1126
rect -416 964 530336 976
rect -416 908 -404 964
rect -348 908 -324 964
rect -268 908 -244 964
rect -188 908 -164 964
rect -108 908 66920 964
rect 66976 908 67000 964
rect 67056 908 67080 964
rect 67136 908 67160 964
rect 67216 908 198848 964
rect 198904 908 198928 964
rect 198984 908 199008 964
rect 199064 908 199088 964
rect 199144 908 330776 964
rect 330832 908 330856 964
rect 330912 908 330936 964
rect 330992 908 331016 964
rect 331072 908 462704 964
rect 462760 908 462784 964
rect 462840 908 462864 964
rect 462920 908 462944 964
rect 463000 908 530028 964
rect 530084 908 530108 964
rect 530164 908 530188 964
rect 530244 908 530268 964
rect 530324 908 530336 964
rect -416 884 530336 908
rect -416 828 -404 884
rect -348 828 -324 884
rect -268 828 -244 884
rect -188 828 -164 884
rect -108 828 66920 884
rect 66976 828 67000 884
rect 67056 828 67080 884
rect 67136 828 67160 884
rect 67216 828 198848 884
rect 198904 828 198928 884
rect 198984 828 199008 884
rect 199064 828 199088 884
rect 199144 828 330776 884
rect 330832 828 330856 884
rect 330912 828 330936 884
rect 330992 828 331016 884
rect 331072 828 462704 884
rect 462760 828 462784 884
rect 462840 828 462864 884
rect 462920 828 462944 884
rect 463000 828 530028 884
rect 530084 828 530108 884
rect 530164 828 530188 884
rect 530244 828 530268 884
rect 530324 828 530336 884
rect -416 804 530336 828
rect -416 748 -404 804
rect -348 748 -324 804
rect -268 748 -244 804
rect -188 748 -164 804
rect -108 748 66920 804
rect 66976 748 67000 804
rect 67056 748 67080 804
rect 67136 748 67160 804
rect 67216 748 198848 804
rect 198904 748 198928 804
rect 198984 748 199008 804
rect 199064 748 199088 804
rect 199144 748 330776 804
rect 330832 748 330856 804
rect 330912 748 330936 804
rect 330992 748 331016 804
rect 331072 748 462704 804
rect 462760 748 462784 804
rect 462840 748 462864 804
rect 462920 748 462944 804
rect 463000 748 530028 804
rect 530084 748 530108 804
rect 530164 748 530188 804
rect 530244 748 530268 804
rect 530324 748 530336 804
rect -416 724 530336 748
rect -416 668 -404 724
rect -348 668 -324 724
rect -268 668 -244 724
rect -188 668 -164 724
rect -108 668 66920 724
rect 66976 668 67000 724
rect 67056 668 67080 724
rect 67136 668 67160 724
rect 67216 668 198848 724
rect 198904 668 198928 724
rect 198984 668 199008 724
rect 199064 668 199088 724
rect 199144 668 330776 724
rect 330832 668 330856 724
rect 330912 668 330936 724
rect 330992 668 331016 724
rect 331072 668 462704 724
rect 462760 668 462784 724
rect 462840 668 462864 724
rect 462920 668 462944 724
rect 463000 668 530028 724
rect 530084 668 530108 724
rect 530164 668 530188 724
rect 530244 668 530268 724
rect 530324 668 530336 724
rect -416 656 530336 668
rect 28625 506 28691 509
rect 122925 506 122991 509
rect 28625 504 122991 506
rect 28625 448 28630 504
rect 28686 448 122930 504
rect 122986 448 122991 504
rect 28625 446 122991 448
rect 28625 443 28691 446
rect 122925 443 122991 446
rect 307661 506 307727 509
rect 400489 506 400555 509
rect 307661 504 400555 506
rect 307661 448 307666 504
rect 307722 448 400494 504
rect 400550 448 400555 504
rect 307661 446 400555 448
rect 307661 443 307727 446
rect 400489 443 400555 446
rect 400673 506 400739 509
rect 403433 506 403499 509
rect 400673 504 403499 506
rect 400673 448 400678 504
rect 400734 448 403438 504
rect 403494 448 403499 504
rect 400673 446 403499 448
rect 400673 443 400739 446
rect 403433 443 403499 446
rect 406377 506 406443 509
rect 409689 506 409755 509
rect 406377 504 409755 506
rect 406377 448 406382 504
rect 406438 448 409694 504
rect 409750 448 409755 504
rect 406377 446 409755 448
rect 406377 443 406443 446
rect 409689 443 409755 446
rect 479701 506 479767 509
rect 482645 506 482711 509
rect 479701 504 482711 506
rect 479701 448 479706 504
rect 479762 448 482650 504
rect 482706 448 482711 504
rect 479701 446 482711 448
rect 479701 443 479767 446
rect 482645 443 482711 446
rect -1076 304 530996 316
rect -1076 248 -1064 304
rect -1008 248 -984 304
rect -928 248 -904 304
rect -848 248 -824 304
rect -768 248 67580 304
rect 67636 248 67660 304
rect 67716 248 67740 304
rect 67796 248 67820 304
rect 67876 248 199508 304
rect 199564 248 199588 304
rect 199644 248 199668 304
rect 199724 248 199748 304
rect 199804 248 331436 304
rect 331492 248 331516 304
rect 331572 248 331596 304
rect 331652 248 331676 304
rect 331732 248 463364 304
rect 463420 248 463444 304
rect 463500 248 463524 304
rect 463580 248 463604 304
rect 463660 248 530688 304
rect 530744 248 530768 304
rect 530824 248 530848 304
rect 530904 248 530928 304
rect 530984 248 530996 304
rect -1076 224 530996 248
rect -1076 168 -1064 224
rect -1008 168 -984 224
rect -928 168 -904 224
rect -848 168 -824 224
rect -768 168 67580 224
rect 67636 168 67660 224
rect 67716 168 67740 224
rect 67796 168 67820 224
rect 67876 168 199508 224
rect 199564 168 199588 224
rect 199644 168 199668 224
rect 199724 168 199748 224
rect 199804 168 331436 224
rect 331492 168 331516 224
rect 331572 168 331596 224
rect 331652 168 331676 224
rect 331732 168 463364 224
rect 463420 168 463444 224
rect 463500 168 463524 224
rect 463580 168 463604 224
rect 463660 168 530688 224
rect 530744 168 530768 224
rect 530824 168 530848 224
rect 530904 168 530928 224
rect 530984 168 530996 224
rect -1076 144 530996 168
rect -1076 88 -1064 144
rect -1008 88 -984 144
rect -928 88 -904 144
rect -848 88 -824 144
rect -768 88 67580 144
rect 67636 88 67660 144
rect 67716 88 67740 144
rect 67796 88 67820 144
rect 67876 88 199508 144
rect 199564 88 199588 144
rect 199644 88 199668 144
rect 199724 88 199748 144
rect 199804 88 331436 144
rect 331492 88 331516 144
rect 331572 88 331596 144
rect 331652 88 331676 144
rect 331732 88 463364 144
rect 463420 88 463444 144
rect 463500 88 463524 144
rect 463580 88 463604 144
rect 463660 88 530688 144
rect 530744 88 530768 144
rect 530824 88 530848 144
rect 530904 88 530928 144
rect 530984 88 530996 144
rect -1076 64 530996 88
rect -1076 8 -1064 64
rect -1008 8 -984 64
rect -928 8 -904 64
rect -848 8 -824 64
rect -768 8 67580 64
rect 67636 8 67660 64
rect 67716 8 67740 64
rect 67796 8 67820 64
rect 67876 8 199508 64
rect 199564 8 199588 64
rect 199644 8 199668 64
rect 199724 8 199748 64
rect 199804 8 331436 64
rect 331492 8 331516 64
rect 331572 8 331596 64
rect 331652 8 331676 64
rect 331732 8 463364 64
rect 463420 8 463444 64
rect 463500 8 463524 64
rect 463580 8 463604 64
rect 463660 8 530688 64
rect 530744 8 530768 64
rect 530824 8 530848 64
rect 530904 8 530928 64
rect 530984 8 530996 64
rect -1076 -4 530996 8
use sky130_fd_sc_hd__diode_2  ANTENNA__00__A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 331936 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__01__A
timestamp 1676037725
transform -1 0 330096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__02__A
timestamp 1676037725
transform -1 0 325496 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__03__A
timestamp 1676037725
transform -1 0 324944 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__04__A
timestamp 1676037725
transform -1 0 323840 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__05__A
timestamp 1676037725
transform -1 0 319792 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__06__A
timestamp 1676037725
transform -1 0 319240 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__07__A
timestamp 1676037725
transform 1 0 317768 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__08__A
timestamp 1676037725
transform 1 0 313996 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__09__A
timestamp 1676037725
transform -1 0 315836 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__10__A
timestamp 1676037725
transform -1 0 313260 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__11__A
timestamp 1676037725
transform -1 0 310500 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__12__A
timestamp 1676037725
transform -1 0 313444 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__13__A
timestamp 1676037725
transform -1 0 311788 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__14__A
timestamp 1676037725
transform 1 0 304152 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__15__A
timestamp 1676037725
transform -1 0 307464 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__16__A
timestamp 1676037725
transform -1 0 303508 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__17__A
timestamp 1676037725
transform -1 0 301944 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__18__A
timestamp 1676037725
transform 1 0 302772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__19__A
timestamp 1676037725
transform -1 0 300932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__20__A
timestamp 1676037725
transform -1 0 298172 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__21__A
timestamp 1676037725
transform -1 0 298724 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__22__A
timestamp 1676037725
transform -1 0 296148 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__23__A
timestamp 1676037725
transform -1 0 357328 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__24__A
timestamp 1676037725
transform -1 0 358248 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__25__A
timestamp 1676037725
transform -1 0 356316 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__26__A
timestamp 1676037725
transform 1 0 353188 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__27__A
timestamp 1676037725
transform -1 0 355212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__28__A
timestamp 1676037725
transform -1 0 352728 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__29__A
timestamp 1676037725
transform -1 0 350612 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__30__A
timestamp 1676037725
transform -1 0 350060 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__31__A
timestamp 1676037725
transform -1 0 348772 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1676037725
transform -1 0 347484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1676037725
transform -1 0 346748 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1676037725
transform 1 0 344908 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1676037725
transform -1 0 343068 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1676037725
transform -1 0 342148 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1676037725
transform 1 0 340676 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1676037725
transform -1 0 338192 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1676037725
transform -1 0 337640 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1676037725
transform -1 0 336444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1676037725
transform -1 0 333224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[0\].u_buf_A
timestamp 1676037725
transform -1 0 2668 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[1\].u_buf_A
timestamp 1676037725
transform -1 0 20700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[2\].u_buf_A
timestamp 1676037725
transform 1 0 37628 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[3\].u_buf_A
timestamp 1676037725
transform -1 0 56764 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[4\].u_buf_A
timestamp 1676037725
transform -1 0 75164 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[5\].u_buf_A
timestamp 1676037725
transform -1 0 92828 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[6\].u_buf_A
timestamp 1676037725
transform 1 0 110676 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[7\].u_buf_A
timestamp 1676037725
transform -1 0 128892 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[8\].u_buf_A
timestamp 1676037725
transform 1 0 145820 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[9\].u_buf_A
timestamp 1676037725
transform -1 0 164404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[10\].u_buf_A
timestamp 1676037725
transform -1 0 182988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[11\].u_buf_A
timestamp 1676037725
transform -1 0 201020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[12\].u_buf_A
timestamp 1676037725
transform -1 0 218224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[13\].u_buf_A
timestamp 1676037725
transform -1 0 237084 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[14\].u_buf_A
timestamp 1676037725
transform 1 0 254012 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[15\].u_buf_A
timestamp 1676037725
transform -1 0 273148 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[16\].u_buf_A
timestamp 1676037725
transform -1 0 291180 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[17\].u_buf_A
timestamp 1676037725
transform -1 0 312524 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[18\].u_buf_A
timestamp 1676037725
transform -1 0 327244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[19\].u_buf_A
timestamp 1676037725
transform -1 0 345644 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[20\].u_buf_A
timestamp 1676037725
transform 1 0 362204 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[21\].u_buf_A
timestamp 1676037725
transform -1 0 380972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[22\].u_buf_A
timestamp 1676037725
transform -1 0 399004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[23\].u_buf_A
timestamp 1676037725
transform 1 0 416300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[24\].u_buf_A
timestamp 1676037725
transform -1 0 435068 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[25\].u_buf_A
timestamp 1676037725
transform -1 0 453468 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[26\].u_buf_A
timestamp 1676037725
transform 1 0 470396 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire1_A
timestamp 1676037725
transform -1 0 394312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire2_A
timestamp 1676037725
transform -1 0 300196 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire3_A
timestamp 1676037725
transform -1 0 205068 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire4_A
timestamp 1676037725
transform -1 0 391828 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire5_A
timestamp 1676037725
transform -1 0 296700 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire6_A
timestamp 1676037725
transform 1 0 201664 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire8_A
timestamp 1676037725
transform -1 0 387320 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire9_A
timestamp 1676037725
transform -1 0 292744 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire10_A
timestamp 1676037725
transform -1 0 198076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire11_A
timestamp 1676037725
transform -1 0 103960 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire12_A
timestamp 1676037725
transform -1 0 409492 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire13_A
timestamp 1676037725
transform 1 0 403972 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire14_A
timestamp 1676037725
transform -1 0 401028 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire15_A
timestamp 1676037725
transform -1 0 306912 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire16_A
timestamp 1676037725
transform -1 0 396796 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire17_A
timestamp 1676037725
transform -1 0 302956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire19_A
timestamp 1676037725
transform -1 0 118404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire20_A
timestamp 1676037725
transform -1 0 213624 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire21_A
timestamp 1676037725
transform -1 0 312340 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire22_A
timestamp 1676037725
transform 1 0 119232 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire23_A
timestamp 1676037725
transform -1 0 214176 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire24_A
timestamp 1676037725
transform -1 0 311420 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire25_A
timestamp 1676037725
transform -1 0 117944 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire26_A
timestamp 1676037725
transform -1 0 212888 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire27_A
timestamp 1676037725
transform -1 0 309212 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire28_A
timestamp 1676037725
transform -1 0 119048 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire29_A
timestamp 1676037725
transform -1 0 213072 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire30_A
timestamp 1676037725
transform -1 0 308844 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire31_A
timestamp 1676037725
transform -1 0 118496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire32_A
timestamp 1676037725
transform -1 0 212520 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire33_A
timestamp 1676037725
transform -1 0 307648 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire34_A
timestamp 1676037725
transform -1 0 117576 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire35_A
timestamp 1676037725
transform -1 0 211140 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire36_A
timestamp 1676037725
transform 1 0 306912 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire37_A
timestamp 1676037725
transform -1 0 117024 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire38_A
timestamp 1676037725
transform -1 0 211692 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire39_A
timestamp 1676037725
transform -1 0 308200 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire40_A
timestamp 1676037725
transform -1 0 115552 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire41_A
timestamp 1676037725
transform -1 0 207000 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire42_A
timestamp 1676037725
transform -1 0 306912 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire43_A
timestamp 1676037725
transform -1 0 113068 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire44_A
timestamp 1676037725
transform -1 0 208380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire45_A
timestamp 1676037725
transform -1 0 305808 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire46_A
timestamp 1676037725
transform -1 0 114448 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire47_A
timestamp 1676037725
transform -1 0 208564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire48_A
timestamp 1676037725
transform -1 0 306360 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire49_A
timestamp 1676037725
transform -1 0 116104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire50_A
timestamp 1676037725
transform -1 0 210496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire51_A
timestamp 1676037725
transform -1 0 304888 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire52_A
timestamp 1676037725
transform -1 0 113896 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire53_A
timestamp 1676037725
transform -1 0 209116 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire54_A
timestamp 1676037725
transform -1 0 305532 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire55_A
timestamp 1676037725
transform -1 0 126500 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire56_A
timestamp 1676037725
transform 1 0 220984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire57_A
timestamp 1676037725
transform 1 0 126132 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire58_A
timestamp 1676037725
transform -1 0 221720 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire60_A
timestamp 1676037725
transform -1 0 125948 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire61_A
timestamp 1676037725
transform -1 0 219604 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire62_A
timestamp 1676037725
transform -1 0 124568 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire63_A
timestamp 1676037725
transform -1 0 220524 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire65_A
timestamp 1676037725
transform 1 0 127236 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire66_A
timestamp 1676037725
transform -1 0 216844 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire67_A
timestamp 1676037725
transform -1 0 125212 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire68_A
timestamp 1676037725
transform -1 0 218592 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire69_A
timestamp 1676037725
transform -1 0 123556 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire70_A
timestamp 1676037725
transform -1 0 217948 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire71_A
timestamp 1676037725
transform -1 0 123280 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire72_A
timestamp 1676037725
transform -1 0 216844 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire73_A
timestamp 1676037725
transform -1 0 122636 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire74_A
timestamp 1676037725
transform -1 0 217396 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire75_A
timestamp 1676037725
transform 1 0 122452 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire76_A
timestamp 1676037725
transform 1 0 217764 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire77_A
timestamp 1676037725
transform -1 0 120336 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire78_A
timestamp 1676037725
transform -1 0 216292 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire80_A
timestamp 1676037725
transform 1 0 122452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire81_A
timestamp 1676037725
transform -1 0 214360 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire83_A
timestamp 1676037725
transform -1 0 121440 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire84_A
timestamp 1676037725
transform -1 0 215464 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire86_A
timestamp 1676037725
transform -1 0 116840 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire87_A
timestamp 1676037725
transform -1 0 215832 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire89_A
timestamp 1676037725
transform -1 0 120888 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire90_A
timestamp 1676037725
transform -1 0 213716 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire91_A
timestamp 1676037725
transform 1 0 309580 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire92_A
timestamp 1676037725
transform -1 0 119600 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire93_A
timestamp 1676037725
transform -1 0 214912 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire94_A
timestamp 1676037725
transform -1 0 309764 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire95_A
timestamp 1676037725
transform 1 0 260176 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire96_A
timestamp 1676037725
transform -1 0 354660 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire97_A
timestamp 1676037725
transform -1 0 448684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire98_A
timestamp 1676037725
transform -1 0 224296 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire99_A
timestamp 1676037725
transform -1 0 318412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire100_A
timestamp 1676037725
transform -1 0 413080 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire101_A
timestamp 1676037725
transform 1 0 205988 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire102_A
timestamp 1676037725
transform -1 0 299736 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire103_A
timestamp 1676037725
transform -1 0 394864 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire104_A
timestamp 1676037725
transform -1 0 170844 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire105_A
timestamp 1676037725
transform -1 0 265788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire106_A
timestamp 1676037725
transform 1 0 359444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire107_A
timestamp 1676037725
transform 1 0 453284 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire108_A
timestamp 1676037725
transform -1 0 152444 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire109_A
timestamp 1676037725
transform -1 0 247388 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire110_A
timestamp 1676037725
transform -1 0 341596 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire111_A
timestamp 1676037725
transform -1 0 435988 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire112_A
timestamp 1676037725
transform -1 0 493580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire113_A
timestamp 1676037725
transform -1 0 475548 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire114_A
timestamp 1676037725
transform -1 0 116380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire115_A
timestamp 1676037725
transform -1 0 211692 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire116_A
timestamp 1676037725
transform -1 0 306360 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire117_A
timestamp 1676037725
transform -1 0 400200 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire118_A
timestamp 1676037725
transform -1 0 440680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire119_A
timestamp 1676037725
transform -1 0 422648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire120_A
timestamp 1676037725
transform -1 0 386584 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire121_A
timestamp 1676037725
transform -1 0 479872 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire122_A
timestamp 1676037725
transform -1 0 368552 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire123_A
timestamp 1676037725
transform -1 0 461932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire124_A
timestamp 1676037725
transform -1 0 332672 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire125_A
timestamp 1676037725
transform -1 0 426604 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire126_A
timestamp 1676037725
transform -1 0 315836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire127_A
timestamp 1676037725
transform -1 0 408572 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire128_A
timestamp 1676037725
transform -1 0 278392 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire129_A
timestamp 1676037725
transform -1 0 372508 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire130_A
timestamp 1676037725
transform -1 0 466624 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire131_A
timestamp 1676037725
transform -1 0 98716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire132_A
timestamp 1676037725
transform -1 0 193660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire133_A
timestamp 1676037725
transform -1 0 287500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire134_A
timestamp 1676037725
transform -1 0 382812 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire135_A
timestamp 1676037725
transform -1 0 251620 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire136_A
timestamp 1676037725
transform -1 0 156860 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire137_A
timestamp 1676037725
transform -1 0 62744 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire138_A
timestamp 1676037725
transform -1 0 255944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire139_A
timestamp 1676037725
transform -1 0 160632 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire140_A
timestamp 1676037725
transform -1 0 66424 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire141_A
timestamp 1676037725
transform -1 0 390540 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire142_A
timestamp 1676037725
transform 1 0 391092 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire143_A
timestamp 1676037725
transform -1 0 258520 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire144_A
timestamp 1676037725
transform -1 0 164956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire145_A
timestamp 1676037725
transform -1 0 70472 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire146_A
timestamp 1676037725
transform -1 0 202860 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire147_A
timestamp 1676037725
transform -1 0 108284 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire148_A
timestamp 1676037725
transform -1 0 393668 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire149_A
timestamp 1676037725
transform -1 0 396244 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire150_A
timestamp 1676037725
transform 1 0 206816 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire151_A
timestamp 1676037725
transform -1 0 112240 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire152_A
timestamp 1676037725
transform 1 0 398084 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire153_A
timestamp 1676037725
transform -1 0 211140 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire154_A
timestamp 1676037725
transform -1 0 116748 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire155_A
timestamp 1676037725
transform -1 0 214728 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire156_A
timestamp 1676037725
transform -1 0 120888 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire157_A
timestamp 1676037725
transform -1 0 221720 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire158_A
timestamp 1676037725
transform -1 0 126868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire159_A
timestamp 1676037725
transform -1 0 225032 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire160_A
timestamp 1676037725
transform -1 0 130364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire161_A
timestamp 1676037725
transform -1 0 36064 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire162_A
timestamp 1676037725
transform -1 0 230920 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire163_A
timestamp 1676037725
transform -1 0 136252 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire164_A
timestamp 1676037725
transform -1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire165_A
timestamp 1676037725
transform -1 0 237912 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire166_A
timestamp 1676037725
transform -1 0 143244 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire167_A
timestamp 1676037725
transform -1 0 48484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire168_A
timestamp 1676037725
transform -1 0 243064 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire169_A
timestamp 1676037725
transform -1 0 148396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire170_A
timestamp 1676037725
transform -1 0 54004 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire171_A
timestamp 1676037725
transform -1 0 248216 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire172_A
timestamp 1676037725
transform -1 0 152904 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire173_A
timestamp 1676037725
transform -1 0 58328 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire174_A
timestamp 1676037725
transform 1 0 262292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire175_A
timestamp 1676037725
transform 1 0 167992 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire176_A
timestamp 1676037725
transform -1 0 74612 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11
timestamp 1676037725
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1676037725
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1676037725
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1676037725
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1676037725
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1676037725
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1676037725
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_197 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_207
timestamp 1676037725
transform 1 0 20148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_213
timestamp 1676037725
transform 1 0 20700 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1676037725
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1676037725
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1676037725
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1676037725
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1676037725
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1676037725
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1676037725
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1676037725
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1676037725
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_377 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_380
timestamp 1676037725
transform 1 0 36064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_403
timestamp 1676037725
transform 1 0 38180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_415
timestamp 1676037725
transform 1 0 39284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1676037725
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_433
timestamp 1676037725
transform 1 0 40940 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_441
timestamp 1676037725
transform 1 0 41676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1676037725
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_457
timestamp 1676037725
transform 1 0 43148 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_469
timestamp 1676037725
transform 1 0 44252 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1676037725
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1676037725
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1676037725
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_515
timestamp 1676037725
transform 1 0 48484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_525
timestamp 1676037725
transform 1 0 49404 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_531
timestamp 1676037725
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1676037725
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_545
timestamp 1676037725
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1676037725
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_561
timestamp 1676037725
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_575
timestamp 1676037725
transform 1 0 54004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1676037725
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_589
timestamp 1676037725
transform 1 0 55292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_599
timestamp 1676037725
transform 1 0 56212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_605
timestamp 1676037725
transform 1 0 56764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1676037725
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_617
timestamp 1676037725
transform 1 0 57868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_622
timestamp 1676037725
transform 1 0 58328 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_632
timestamp 1676037725
transform 1 0 59248 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_645
timestamp 1676037725
transform 1 0 60444 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_657
timestamp 1676037725
transform 1 0 61548 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_665
timestamp 1676037725
transform 1 0 62284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_670
timestamp 1676037725
transform 1 0 62744 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_673
timestamp 1676037725
transform 1 0 63020 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_681
timestamp 1676037725
transform 1 0 63756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_693
timestamp 1676037725
transform 1 0 64860 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_699
timestamp 1676037725
transform 1 0 65412 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_701
timestamp 1676037725
transform 1 0 65596 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_707
timestamp 1676037725
transform 1 0 66148 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_710
timestamp 1676037725
transform 1 0 66424 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_720
timestamp 1676037725
transform 1 0 67344 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_729
timestamp 1676037725
transform 1 0 68172 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_741
timestamp 1676037725
transform 1 0 69276 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_749
timestamp 1676037725
transform 1 0 70012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_754
timestamp 1676037725
transform 1 0 70472 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_757
timestamp 1676037725
transform 1 0 70748 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_768
timestamp 1676037725
transform 1 0 71760 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_780
timestamp 1676037725
transform 1 0 72864 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_785
timestamp 1676037725
transform 1 0 73324 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_795
timestamp 1676037725
transform 1 0 74244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_808
timestamp 1676037725
transform 1 0 75440 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_813
timestamp 1676037725
transform 1 0 75900 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_825
timestamp 1676037725
transform 1 0 77004 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_837
timestamp 1676037725
transform 1 0 78108 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_841
timestamp 1676037725
transform 1 0 78476 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_853
timestamp 1676037725
transform 1 0 79580 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_865
timestamp 1676037725
transform 1 0 80684 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_869
timestamp 1676037725
transform 1 0 81052 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_881
timestamp 1676037725
transform 1 0 82156 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_893
timestamp 1676037725
transform 1 0 83260 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_897
timestamp 1676037725
transform 1 0 83628 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_909
timestamp 1676037725
transform 1 0 84732 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_921
timestamp 1676037725
transform 1 0 85836 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_925
timestamp 1676037725
transform 1 0 86204 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_937
timestamp 1676037725
transform 1 0 87308 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_949
timestamp 1676037725
transform 1 0 88412 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_953
timestamp 1676037725
transform 1 0 88780 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_965
timestamp 1676037725
transform 1 0 89884 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_977
timestamp 1676037725
transform 1 0 90988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_981
timestamp 1676037725
transform 1 0 91356 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_987
timestamp 1676037725
transform 1 0 91908 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_991
timestamp 1676037725
transform 1 0 92276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_997
timestamp 1676037725
transform 1 0 92828 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1005
timestamp 1676037725
transform 1 0 93564 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1009
timestamp 1676037725
transform 1 0 93932 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1021
timestamp 1676037725
transform 1 0 95036 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1033
timestamp 1676037725
transform 1 0 96140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1037
timestamp 1676037725
transform 1 0 96508 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1055
timestamp 1676037725
transform 1 0 98164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1061
timestamp 1676037725
transform 1 0 98716 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1065
timestamp 1676037725
transform 1 0 99084 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1077
timestamp 1676037725
transform 1 0 100188 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1089
timestamp 1676037725
transform 1 0 101292 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1093
timestamp 1676037725
transform 1 0 101660 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1105
timestamp 1676037725
transform 1 0 102764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1113
timestamp 1676037725
transform 1 0 103500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1118
timestamp 1676037725
transform 1 0 103960 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1121
timestamp 1676037725
transform 1 0 104236 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1132
timestamp 1676037725
transform 1 0 105248 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1144
timestamp 1676037725
transform 1 0 106352 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1149
timestamp 1676037725
transform 1 0 106812 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1161
timestamp 1676037725
transform 1 0 107916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1174
timestamp 1676037725
transform 1 0 109112 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1177
timestamp 1676037725
transform 1 0 109388 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1187
timestamp 1676037725
transform 1 0 110308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1193
timestamp 1676037725
transform 1 0 110860 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1201
timestamp 1676037725
transform 1 0 111596 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1205
timestamp 1676037725
transform 1 0 111964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1217
timestamp 1676037725
transform 1 0 113068 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1230
timestamp 1676037725
transform 1 0 114264 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1233
timestamp 1676037725
transform 1 0 114540 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1251
timestamp 1676037725
transform 1 0 116196 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1255
timestamp 1676037725
transform 1 0 116564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1258
timestamp 1676037725
transform 1 0 116840 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1261
timestamp 1676037725
transform 1 0 117116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1273
timestamp 1676037725
transform 1 0 118220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1286
timestamp 1676037725
transform 1 0 119416 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1289
timestamp 1676037725
transform 1 0 119692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1301
timestamp 1676037725
transform 1 0 120796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1314
timestamp 1676037725
transform 1 0 121992 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1317
timestamp 1676037725
transform 1 0 122268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1329
timestamp 1676037725
transform 1 0 123372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1342
timestamp 1676037725
transform 1 0 124568 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1345
timestamp 1676037725
transform 1 0 124844 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1353
timestamp 1676037725
transform 1 0 125580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1366
timestamp 1676037725
transform 1 0 126776 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1373
timestamp 1676037725
transform 1 0 127420 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1383
timestamp 1676037725
transform 1 0 128340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1389
timestamp 1676037725
transform 1 0 128892 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1397
timestamp 1676037725
transform 1 0 129628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1401
timestamp 1676037725
transform 1 0 129996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1405
timestamp 1676037725
transform 1 0 130364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1418
timestamp 1676037725
transform 1 0 131560 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1426
timestamp 1676037725
transform 1 0 132296 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1429
timestamp 1676037725
transform 1 0 132572 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1441
timestamp 1676037725
transform 1 0 133676 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1453
timestamp 1676037725
transform 1 0 134780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1457
timestamp 1676037725
transform 1 0 135148 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1465
timestamp 1676037725
transform 1 0 135884 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1469
timestamp 1676037725
transform 1 0 136252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1482
timestamp 1676037725
transform 1 0 137448 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1485
timestamp 1676037725
transform 1 0 137724 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1497
timestamp 1676037725
transform 1 0 138828 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1509
timestamp 1676037725
transform 1 0 139932 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1513
timestamp 1676037725
transform 1 0 140300 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1525
timestamp 1676037725
transform 1 0 141404 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1537
timestamp 1676037725
transform 1 0 142508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1541
timestamp 1676037725
transform 1 0 142876 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1554
timestamp 1676037725
transform 1 0 144072 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1566
timestamp 1676037725
transform 1 0 145176 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1569
timestamp 1676037725
transform 1 0 145452 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1579
timestamp 1676037725
transform 1 0 146372 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1591
timestamp 1676037725
transform 1 0 147476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1595
timestamp 1676037725
transform 1 0 147844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1597
timestamp 1676037725
transform 1 0 148028 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1601
timestamp 1676037725
transform 1 0 148396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1614
timestamp 1676037725
transform 1 0 149592 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1622
timestamp 1676037725
transform 1 0 150328 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1625
timestamp 1676037725
transform 1 0 150604 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1643
timestamp 1676037725
transform 1 0 152260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1647
timestamp 1676037725
transform 1 0 152628 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1650
timestamp 1676037725
transform 1 0 152904 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1653
timestamp 1676037725
transform 1 0 153180 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1664
timestamp 1676037725
transform 1 0 154192 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1676
timestamp 1676037725
transform 1 0 155296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1681
timestamp 1676037725
transform 1 0 155756 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1689
timestamp 1676037725
transform 1 0 156492 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1693
timestamp 1676037725
transform 1 0 156860 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1706
timestamp 1676037725
transform 1 0 158056 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1709
timestamp 1676037725
transform 1 0 158332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1721
timestamp 1676037725
transform 1 0 159436 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1729
timestamp 1676037725
transform 1 0 160172 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1734
timestamp 1676037725
transform 1 0 160632 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1737
timestamp 1676037725
transform 1 0 160908 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1749
timestamp 1676037725
transform 1 0 162012 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1761
timestamp 1676037725
transform 1 0 163116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1765
timestamp 1676037725
transform 1 0 163484 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1775
timestamp 1676037725
transform 1 0 164404 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1790
timestamp 1676037725
transform 1 0 165784 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1793
timestamp 1676037725
transform 1 0 166060 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1805
timestamp 1676037725
transform 1 0 167164 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1817
timestamp 1676037725
transform 1 0 168268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1821
timestamp 1676037725
transform 1 0 168636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1839
timestamp 1676037725
transform 1 0 170292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1845
timestamp 1676037725
transform 1 0 170844 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1849
timestamp 1676037725
transform 1 0 171212 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1861
timestamp 1676037725
transform 1 0 172316 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1873
timestamp 1676037725
transform 1 0 173420 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1877
timestamp 1676037725
transform 1 0 173788 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1889
timestamp 1676037725
transform 1 0 174892 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1901
timestamp 1676037725
transform 1 0 175996 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1905
timestamp 1676037725
transform 1 0 176364 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1917
timestamp 1676037725
transform 1 0 177468 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1929
timestamp 1676037725
transform 1 0 178572 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1933
timestamp 1676037725
transform 1 0 178940 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1945
timestamp 1676037725
transform 1 0 180044 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1957
timestamp 1676037725
transform 1 0 181148 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1961
timestamp 1676037725
transform 1 0 181516 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1971
timestamp 1676037725
transform 1 0 182436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1977
timestamp 1676037725
transform 1 0 182988 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1985
timestamp 1676037725
transform 1 0 183724 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1989
timestamp 1676037725
transform 1 0 184092 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2001
timestamp 1676037725
transform 1 0 185196 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2013
timestamp 1676037725
transform 1 0 186300 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2017
timestamp 1676037725
transform 1 0 186668 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2029
timestamp 1676037725
transform 1 0 187772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2041
timestamp 1676037725
transform 1 0 188876 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2045
timestamp 1676037725
transform 1 0 189244 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2057
timestamp 1676037725
transform 1 0 190348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2069
timestamp 1676037725
transform 1 0 191452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2073
timestamp 1676037725
transform 1 0 191820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2087
timestamp 1676037725
transform 1 0 193108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2093
timestamp 1676037725
transform 1 0 193660 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2099
timestamp 1676037725
transform 1 0 194212 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2101
timestamp 1676037725
transform 1 0 194396 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2113
timestamp 1676037725
transform 1 0 195500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2125
timestamp 1676037725
transform 1 0 196604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2129
timestamp 1676037725
transform 1 0 196972 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2137
timestamp 1676037725
transform 1 0 197708 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2141
timestamp 1676037725
transform 1 0 198076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2154
timestamp 1676037725
transform 1 0 199272 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2157
timestamp 1676037725
transform 1 0 199548 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2163
timestamp 1676037725
transform 1 0 200100 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2167
timestamp 1676037725
transform 1 0 200468 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2173
timestamp 1676037725
transform 1 0 201020 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2181
timestamp 1676037725
transform 1 0 201756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2185
timestamp 1676037725
transform 1 0 202124 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2193
timestamp 1676037725
transform 1 0 202860 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2206
timestamp 1676037725
transform 1 0 204056 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2213
timestamp 1676037725
transform 1 0 204700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2217
timestamp 1676037725
transform 1 0 205068 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2230
timestamp 1676037725
transform 1 0 206264 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2238
timestamp 1676037725
transform 1 0 207000 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2241
timestamp 1676037725
transform 1 0 207276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2253
timestamp 1676037725
transform 1 0 208380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2266
timestamp 1676037725
transform 1 0 209576 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2269
timestamp 1676037725
transform 1 0 209852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2283
timestamp 1676037725
transform 1 0 211140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2293
timestamp 1676037725
transform 1 0 212060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2297
timestamp 1676037725
transform 1 0 212428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2309
timestamp 1676037725
transform 1 0 213532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2322
timestamp 1676037725
transform 1 0 214728 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2325
timestamp 1676037725
transform 1 0 215004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2337
timestamp 1676037725
transform 1 0 216108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2350
timestamp 1676037725
transform 1 0 217304 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2353
timestamp 1676037725
transform 1 0 217580 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2363
timestamp 1676037725
transform 1 0 218500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2378
timestamp 1676037725
transform 1 0 219880 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2381
timestamp 1676037725
transform 1 0 220156 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2392
timestamp 1676037725
transform 1 0 221168 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2398
timestamp 1676037725
transform 1 0 221720 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2406
timestamp 1676037725
transform 1 0 222456 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2409
timestamp 1676037725
transform 1 0 222732 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2420
timestamp 1676037725
transform 1 0 223744 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2426
timestamp 1676037725
transform 1 0 224296 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2434
timestamp 1676037725
transform 1 0 225032 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2437
timestamp 1676037725
transform 1 0 225308 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2448
timestamp 1676037725
transform 1 0 226320 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2460
timestamp 1676037725
transform 1 0 227424 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2465
timestamp 1676037725
transform 1 0 227884 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2477
timestamp 1676037725
transform 1 0 228988 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2489
timestamp 1676037725
transform 1 0 230092 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2493
timestamp 1676037725
transform 1 0 230460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2498
timestamp 1676037725
transform 1 0 230920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2511
timestamp 1676037725
transform 1 0 232116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2519
timestamp 1676037725
transform 1 0 232852 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2521
timestamp 1676037725
transform 1 0 233036 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2533
timestamp 1676037725
transform 1 0 234140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2545
timestamp 1676037725
transform 1 0 235244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2549
timestamp 1676037725
transform 1 0 235612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2559
timestamp 1676037725
transform 1 0 236532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2565
timestamp 1676037725
transform 1 0 237084 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2571
timestamp 1676037725
transform 1 0 237636 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2574
timestamp 1676037725
transform 1 0 237912 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2577
timestamp 1676037725
transform 1 0 238188 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2588
timestamp 1676037725
transform 1 0 239200 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2600
timestamp 1676037725
transform 1 0 240304 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2605
timestamp 1676037725
transform 1 0 240764 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2617
timestamp 1676037725
transform 1 0 241868 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2625
timestamp 1676037725
transform 1 0 242604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2630
timestamp 1676037725
transform 1 0 243064 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2633
timestamp 1676037725
transform 1 0 243340 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2644
timestamp 1676037725
transform 1 0 244352 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2656
timestamp 1676037725
transform 1 0 245456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2661
timestamp 1676037725
transform 1 0 245916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2675
timestamp 1676037725
transform 1 0 247204 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2683
timestamp 1676037725
transform 1 0 247940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2686
timestamp 1676037725
transform 1 0 248216 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2689
timestamp 1676037725
transform 1 0 248492 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2700
timestamp 1676037725
transform 1 0 249504 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2712
timestamp 1676037725
transform 1 0 250608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2717
timestamp 1676037725
transform 1 0 251068 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2732
timestamp 1676037725
transform 1 0 252448 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2745
timestamp 1676037725
transform 1 0 253644 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2755
timestamp 1676037725
transform 1 0 254564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2767
timestamp 1676037725
transform 1 0 255668 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2770
timestamp 1676037725
transform 1 0 255944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2773
timestamp 1676037725
transform 1 0 256220 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2784
timestamp 1676037725
transform 1 0 257232 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2798
timestamp 1676037725
transform 1 0 258520 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2801
timestamp 1676037725
transform 1 0 258796 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2816
timestamp 1676037725
transform 1 0 260176 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2829
timestamp 1676037725
transform 1 0 261372 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2837
timestamp 1676037725
transform 1 0 262108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2841
timestamp 1676037725
transform 1 0 262476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2854
timestamp 1676037725
transform 1 0 263672 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2857
timestamp 1676037725
transform 1 0 263948 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2871
timestamp 1676037725
transform 1 0 265236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2877
timestamp 1676037725
transform 1 0 265788 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2883
timestamp 1676037725
transform 1 0 266340 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2885
timestamp 1676037725
transform 1 0 266524 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2897
timestamp 1676037725
transform 1 0 267628 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2909
timestamp 1676037725
transform 1 0 268732 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2913
timestamp 1676037725
transform 1 0 269100 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2925
timestamp 1676037725
transform 1 0 270204 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2937
timestamp 1676037725
transform 1 0 271308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2941
timestamp 1676037725
transform 1 0 271676 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2951
timestamp 1676037725
transform 1 0 272596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2957
timestamp 1676037725
transform 1 0 273148 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2965
timestamp 1676037725
transform 1 0 273884 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2969
timestamp 1676037725
transform 1 0 274252 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2981
timestamp 1676037725
transform 1 0 275356 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2993
timestamp 1676037725
transform 1 0 276460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2997
timestamp 1676037725
transform 1 0 276828 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3008
timestamp 1676037725
transform 1 0 277840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3014
timestamp 1676037725
transform 1 0 278392 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3022
timestamp 1676037725
transform 1 0 279128 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3025
timestamp 1676037725
transform 1 0 279404 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3037
timestamp 1676037725
transform 1 0 280508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3049
timestamp 1676037725
transform 1 0 281612 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3053
timestamp 1676037725
transform 1 0 281980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3065
timestamp 1676037725
transform 1 0 283084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3077
timestamp 1676037725
transform 1 0 284188 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3081
timestamp 1676037725
transform 1 0 284556 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3093
timestamp 1676037725
transform 1 0 285660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3104
timestamp 1676037725
transform 1 0 286672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3109
timestamp 1676037725
transform 1 0 287132 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3113
timestamp 1676037725
transform 1 0 287500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3125
timestamp 1676037725
transform 1 0 288604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3133
timestamp 1676037725
transform 1 0 289340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3137
timestamp 1676037725
transform 1 0 289708 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3147
timestamp 1676037725
transform 1 0 290628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3153
timestamp 1676037725
transform 1 0 291180 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3161
timestamp 1676037725
transform 1 0 291916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3165
timestamp 1676037725
transform 1 0 292284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3170
timestamp 1676037725
transform 1 0 292744 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3183
timestamp 1676037725
transform 1 0 293940 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3191
timestamp 1676037725
transform 1 0 294676 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3193
timestamp 1676037725
transform 1 0 294860 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3205
timestamp 1676037725
transform 1 0 295964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3218
timestamp 1676037725
transform 1 0 297160 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3221
timestamp 1676037725
transform 1 0 297436 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3229
timestamp 1676037725
transform 1 0 298172 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3246
timestamp 1676037725
transform 1 0 299736 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3249
timestamp 1676037725
transform 1 0 300012 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3260
timestamp 1676037725
transform 1 0 301024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3270
timestamp 1676037725
transform 1 0 301944 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3277
timestamp 1676037725
transform 1 0 302588 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3281
timestamp 1676037725
transform 1 0 302956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3294
timestamp 1676037725
transform 1 0 304152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3302
timestamp 1676037725
transform 1 0 304888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3305
timestamp 1676037725
transform 1 0 305164 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3316
timestamp 1676037725
transform 1 0 306176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3320
timestamp 1676037725
transform 1 0 306544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3330
timestamp 1676037725
transform 1 0 307464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3333
timestamp 1676037725
transform 1 0 307740 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3343
timestamp 1676037725
transform 1 0 308660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3353
timestamp 1676037725
transform 1 0 309580 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3359
timestamp 1676037725
transform 1 0 310132 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3361
timestamp 1676037725
transform 1 0 310316 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3369
timestamp 1676037725
transform 1 0 311052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3379
timestamp 1676037725
transform 1 0 311972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3385
timestamp 1676037725
transform 1 0 312524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3389
timestamp 1676037725
transform 1 0 312892 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3400
timestamp 1676037725
transform 1 0 313904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3410
timestamp 1676037725
transform 1 0 314824 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3417
timestamp 1676037725
transform 1 0 315468 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3421
timestamp 1676037725
transform 1 0 315836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3442
timestamp 1676037725
transform 1 0 317768 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3445
timestamp 1676037725
transform 1 0 318044 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3449
timestamp 1676037725
transform 1 0 318412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3456
timestamp 1676037725
transform 1 0 319056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3464
timestamp 1676037725
transform 1 0 319792 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3473
timestamp 1676037725
transform 1 0 320620 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3485
timestamp 1676037725
transform 1 0 321724 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3497
timestamp 1676037725
transform 1 0 322828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3501
timestamp 1676037725
transform 1 0 323196 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3506
timestamp 1676037725
transform 1 0 323656 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3514
timestamp 1676037725
transform 1 0 324392 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3518
timestamp 1676037725
transform 1 0 324760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3526
timestamp 1676037725
transform 1 0 325496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3529
timestamp 1676037725
transform 1 0 325772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3539
timestamp 1676037725
transform 1 0 326692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3545
timestamp 1676037725
transform 1 0 327244 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3553
timestamp 1676037725
transform 1 0 327980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3557
timestamp 1676037725
transform 1 0 328348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3565
timestamp 1676037725
transform 1 0 329084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3570
timestamp 1676037725
transform 1 0 329544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3576
timestamp 1676037725
transform 1 0 330096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3585
timestamp 1676037725
transform 1 0 330924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3596
timestamp 1676037725
transform 1 0 331936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3604
timestamp 1676037725
transform 1 0 332672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3610
timestamp 1676037725
transform 1 0 333224 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3613
timestamp 1676037725
transform 1 0 333500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3625
timestamp 1676037725
transform 1 0 334604 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3631
timestamp 1676037725
transform 1 0 335156 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3636
timestamp 1676037725
transform 1 0 335616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3641
timestamp 1676037725
transform 1 0 336076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3645
timestamp 1676037725
transform 1 0 336444 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3651
timestamp 1676037725
transform 1 0 336996 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3656
timestamp 1676037725
transform 1 0 337456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3664
timestamp 1676037725
transform 1 0 338192 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3669
timestamp 1676037725
transform 1 0 338652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3681
timestamp 1676037725
transform 1 0 339756 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3691
timestamp 1676037725
transform 1 0 340676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3695
timestamp 1676037725
transform 1 0 341044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3697
timestamp 1676037725
transform 1 0 341228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3703
timestamp 1676037725
transform 1 0 341780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3711
timestamp 1676037725
transform 1 0 342516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3717
timestamp 1676037725
transform 1 0 343068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3723
timestamp 1676037725
transform 1 0 343620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3725
timestamp 1676037725
transform 1 0 343804 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3735
timestamp 1676037725
transform 1 0 344724 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3743
timestamp 1676037725
transform 1 0 345460 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3748
timestamp 1676037725
transform 1 0 345920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3753
timestamp 1676037725
transform 1 0 346380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3759
timestamp 1676037725
transform 1 0 346932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3765
timestamp 1676037725
transform 1 0 347484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3777
timestamp 1676037725
transform 1 0 348588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3781
timestamp 1676037725
transform 1 0 348956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3791
timestamp 1676037725
transform 1 0 349876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3799
timestamp 1676037725
transform 1 0 350612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3807
timestamp 1676037725
transform 1 0 351348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3809
timestamp 1676037725
transform 1 0 351532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3815
timestamp 1676037725
transform 1 0 352084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3820
timestamp 1676037725
transform 1 0 352544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3824
timestamp 1676037725
transform 1 0 352912 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3834
timestamp 1676037725
transform 1 0 353832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3837
timestamp 1676037725
transform 1 0 354108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3843
timestamp 1676037725
transform 1 0 354660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3849
timestamp 1676037725
transform 1 0 355212 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3859
timestamp 1676037725
transform 1 0 356132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3863
timestamp 1676037725
transform 1 0 356500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3865
timestamp 1676037725
transform 1 0 356684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3872
timestamp 1676037725
transform 1 0 357328 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3876
timestamp 1676037725
transform 1 0 357696 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3886
timestamp 1676037725
transform 1 0 358616 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3893
timestamp 1676037725
transform 1 0 359260 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3897
timestamp 1676037725
transform 1 0 359628 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3909
timestamp 1676037725
transform 1 0 360732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3917
timestamp 1676037725
transform 1 0 361468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3921
timestamp 1676037725
transform 1 0 361836 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3931
timestamp 1676037725
transform 1 0 362756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3943
timestamp 1676037725
transform 1 0 363860 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3947
timestamp 1676037725
transform 1 0 364228 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3949
timestamp 1676037725
transform 1 0 364412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3961
timestamp 1676037725
transform 1 0 365516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3973
timestamp 1676037725
transform 1 0 366620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3977
timestamp 1676037725
transform 1 0 366988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3988
timestamp 1676037725
transform 1 0 368000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3994
timestamp 1676037725
transform 1 0 368552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4002
timestamp 1676037725
transform 1 0 369288 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4005
timestamp 1676037725
transform 1 0 369564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4017
timestamp 1676037725
transform 1 0 370668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4030
timestamp 1676037725
transform 1 0 371864 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4033
timestamp 1676037725
transform 1 0 372140 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4037
timestamp 1676037725
transform 1 0 372508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4049
timestamp 1676037725
transform 1 0 373612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4057
timestamp 1676037725
transform 1 0 374348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4061
timestamp 1676037725
transform 1 0 374716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4073
timestamp 1676037725
transform 1 0 375820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4085
timestamp 1676037725
transform 1 0 376924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4089
timestamp 1676037725
transform 1 0 377292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4101
timestamp 1676037725
transform 1 0 378396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4113
timestamp 1676037725
transform 1 0 379500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4117
timestamp 1676037725
transform 1 0 379868 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4127
timestamp 1676037725
transform 1 0 380788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4140
timestamp 1676037725
transform 1 0 381984 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4145
timestamp 1676037725
transform 1 0 382444 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4149
timestamp 1676037725
transform 1 0 382812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4161
timestamp 1676037725
transform 1 0 383916 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4169
timestamp 1676037725
transform 1 0 384652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4173
timestamp 1676037725
transform 1 0 385020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4184
timestamp 1676037725
transform 1 0 386032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4190
timestamp 1676037725
transform 1 0 386584 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4198
timestamp 1676037725
transform 1 0 387320 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4201
timestamp 1676037725
transform 1 0 387596 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4212
timestamp 1676037725
transform 1 0 388608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4216
timestamp 1676037725
transform 1 0 388976 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4223
timestamp 1676037725
transform 1 0 389620 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4227
timestamp 1676037725
transform 1 0 389988 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4229
timestamp 1676037725
transform 1 0 390172 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4233
timestamp 1676037725
transform 1 0 390540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4237
timestamp 1676037725
transform 1 0 390908 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4247
timestamp 1676037725
transform 1 0 391828 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4255
timestamp 1676037725
transform 1 0 392564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4257
timestamp 1676037725
transform 1 0 392748 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4265
timestamp 1676037725
transform 1 0 393484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4277
timestamp 1676037725
transform 1 0 394588 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4283
timestamp 1676037725
transform 1 0 395140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4285
timestamp 1676037725
transform 1 0 395324 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4293
timestamp 1676037725
transform 1 0 396060 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4310
timestamp 1676037725
transform 1 0 397624 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4313
timestamp 1676037725
transform 1 0 397900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4323
timestamp 1676037725
transform 1 0 398820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4336
timestamp 1676037725
transform 1 0 400016 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4341
timestamp 1676037725
transform 1 0 400476 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4356
timestamp 1676037725
transform 1 0 401856 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4369
timestamp 1676037725
transform 1 0 403052 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4377
timestamp 1676037725
transform 1 0 403788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4381
timestamp 1676037725
transform 1 0 404156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4394
timestamp 1676037725
transform 1 0 405352 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4397
timestamp 1676037725
transform 1 0 405628 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4409
timestamp 1676037725
transform 1 0 406732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4422
timestamp 1676037725
transform 1 0 407928 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4425
timestamp 1676037725
transform 1 0 408204 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4433
timestamp 1676037725
transform 1 0 408940 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4439
timestamp 1676037725
transform 1 0 409492 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4451
timestamp 1676037725
transform 1 0 410596 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4453
timestamp 1676037725
transform 1 0 410780 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4461
timestamp 1676037725
transform 1 0 411516 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4472
timestamp 1676037725
transform 1 0 412528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4478
timestamp 1676037725
transform 1 0 413080 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4481
timestamp 1676037725
transform 1 0 413356 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4493
timestamp 1676037725
transform 1 0 414460 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4505
timestamp 1676037725
transform 1 0 415564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4509
timestamp 1676037725
transform 1 0 415932 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4519
timestamp 1676037725
transform 1 0 416852 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4531
timestamp 1676037725
transform 1 0 417956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4535
timestamp 1676037725
transform 1 0 418324 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4537
timestamp 1676037725
transform 1 0 418508 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4549
timestamp 1676037725
transform 1 0 419612 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4561
timestamp 1676037725
transform 1 0 420716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4565
timestamp 1676037725
transform 1 0 421084 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4576
timestamp 1676037725
transform 1 0 422096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4582
timestamp 1676037725
transform 1 0 422648 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4590
timestamp 1676037725
transform 1 0 423384 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4593
timestamp 1676037725
transform 1 0 423660 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4605
timestamp 1676037725
transform 1 0 424764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4617
timestamp 1676037725
transform 1 0 425868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4621
timestamp 1676037725
transform 1 0 426236 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4625
timestamp 1676037725
transform 1 0 426604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4637
timestamp 1676037725
transform 1 0 427708 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4645
timestamp 1676037725
transform 1 0 428444 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4649
timestamp 1676037725
transform 1 0 428812 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4661
timestamp 1676037725
transform 1 0 429916 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4673
timestamp 1676037725
transform 1 0 431020 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4677
timestamp 1676037725
transform 1 0 431388 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4689
timestamp 1676037725
transform 1 0 432492 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4701
timestamp 1676037725
transform 1 0 433596 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4705
timestamp 1676037725
transform 1 0 433964 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4715
timestamp 1676037725
transform 1 0 434884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4725
timestamp 1676037725
transform 1 0 435804 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4731
timestamp 1676037725
transform 1 0 436356 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4733
timestamp 1676037725
transform 1 0 436540 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4745
timestamp 1676037725
transform 1 0 437644 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4757
timestamp 1676037725
transform 1 0 438748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4761
timestamp 1676037725
transform 1 0 439116 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4772
timestamp 1676037725
transform 1 0 440128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4778
timestamp 1676037725
transform 1 0 440680 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4786
timestamp 1676037725
transform 1 0 441416 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4789
timestamp 1676037725
transform 1 0 441692 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4801
timestamp 1676037725
transform 1 0 442796 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4813
timestamp 1676037725
transform 1 0 443900 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4817
timestamp 1676037725
transform 1 0 444268 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4829
timestamp 1676037725
transform 1 0 445372 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4841
timestamp 1676037725
transform 1 0 446476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4845
timestamp 1676037725
transform 1 0 446844 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4859
timestamp 1676037725
transform 1 0 448132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4865
timestamp 1676037725
transform 1 0 448684 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4871
timestamp 1676037725
transform 1 0 449236 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4873
timestamp 1676037725
transform 1 0 449420 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4885
timestamp 1676037725
transform 1 0 450524 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4897
timestamp 1676037725
transform 1 0 451628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4901
timestamp 1676037725
transform 1 0 451996 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4911
timestamp 1676037725
transform 1 0 452916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4917
timestamp 1676037725
transform 1 0 453468 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4925
timestamp 1676037725
transform 1 0 454204 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4929
timestamp 1676037725
transform 1 0 454572 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4941
timestamp 1676037725
transform 1 0 455676 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4953
timestamp 1676037725
transform 1 0 456780 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4957
timestamp 1676037725
transform 1 0 457148 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4969
timestamp 1676037725
transform 1 0 458252 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4981
timestamp 1676037725
transform 1 0 459356 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4985
timestamp 1676037725
transform 1 0 459724 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5003
timestamp 1676037725
transform 1 0 461380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5009
timestamp 1676037725
transform 1 0 461932 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5013
timestamp 1676037725
transform 1 0 462300 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5025
timestamp 1676037725
transform 1 0 463404 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5037
timestamp 1676037725
transform 1 0 464508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5041
timestamp 1676037725
transform 1 0 464876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5047
timestamp 1676037725
transform 1 0 465428 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5054
timestamp 1676037725
transform 1 0 466072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5060
timestamp 1676037725
transform 1 0 466624 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5069
timestamp 1676037725
transform 1 0 467452 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5081
timestamp 1676037725
transform 1 0 468556 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5093
timestamp 1676037725
transform 1 0 469660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5097
timestamp 1676037725
transform 1 0 470028 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5107
timestamp 1676037725
transform 1 0 470948 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5119
timestamp 1676037725
transform 1 0 472052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5123
timestamp 1676037725
transform 1 0 472420 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5125
timestamp 1676037725
transform 1 0 472604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5137
timestamp 1676037725
transform 1 0 473708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5141
timestamp 1676037725
transform 1 0 474076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5148
timestamp 1676037725
transform 1 0 474720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5153
timestamp 1676037725
transform 1 0 475180 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5157
timestamp 1676037725
transform 1 0 475548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5169
timestamp 1676037725
transform 1 0 476652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5177
timestamp 1676037725
transform 1 0 477388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5181
timestamp 1676037725
transform 1 0 477756 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5189
timestamp 1676037725
transform 1 0 478492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5198
timestamp 1676037725
transform 1 0 479320 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5204
timestamp 1676037725
transform 1 0 479872 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5209
timestamp 1676037725
transform 1 0 480332 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5221
timestamp 1676037725
transform 1 0 481436 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5233
timestamp 1676037725
transform 1 0 482540 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5237
timestamp 1676037725
transform 1 0 482908 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5249
timestamp 1676037725
transform 1 0 484012 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5261
timestamp 1676037725
transform 1 0 485116 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5265
timestamp 1676037725
transform 1 0 485484 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5277
timestamp 1676037725
transform 1 0 486588 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5289
timestamp 1676037725
transform 1 0 487692 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5293
timestamp 1676037725
transform 1 0 488060 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5305
timestamp 1676037725
transform 1 0 489164 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5317
timestamp 1676037725
transform 1 0 490268 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5321
timestamp 1676037725
transform 1 0 490636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5333
timestamp 1676037725
transform 1 0 491740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5342
timestamp 1676037725
transform 1 0 492568 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5349
timestamp 1676037725
transform 1 0 493212 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5353
timestamp 1676037725
transform 1 0 493580 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5365
timestamp 1676037725
transform 1 0 494684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5373
timestamp 1676037725
transform 1 0 495420 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5377
timestamp 1676037725
transform 1 0 495788 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5389
timestamp 1676037725
transform 1 0 496892 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5401
timestamp 1676037725
transform 1 0 497996 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5405
timestamp 1676037725
transform 1 0 498364 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5417
timestamp 1676037725
transform 1 0 499468 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5429
timestamp 1676037725
transform 1 0 500572 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5433
timestamp 1676037725
transform 1 0 500940 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5445
timestamp 1676037725
transform 1 0 502044 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5457
timestamp 1676037725
transform 1 0 503148 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5461
timestamp 1676037725
transform 1 0 503516 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5473
timestamp 1676037725
transform 1 0 504620 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5485
timestamp 1676037725
transform 1 0 505724 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5489
timestamp 1676037725
transform 1 0 506092 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5501
timestamp 1676037725
transform 1 0 507196 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5513
timestamp 1676037725
transform 1 0 508300 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5517
timestamp 1676037725
transform 1 0 508668 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5529
timestamp 1676037725
transform 1 0 509772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5541
timestamp 1676037725
transform 1 0 510876 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5545
timestamp 1676037725
transform 1 0 511244 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5557
timestamp 1676037725
transform 1 0 512348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5569
timestamp 1676037725
transform 1 0 513452 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5573
timestamp 1676037725
transform 1 0 513820 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5585
timestamp 1676037725
transform 1 0 514924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5597
timestamp 1676037725
transform 1 0 516028 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5601
timestamp 1676037725
transform 1 0 516396 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5613
timestamp 1676037725
transform 1 0 517500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5625
timestamp 1676037725
transform 1 0 518604 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5629
timestamp 1676037725
transform 1 0 518972 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5641
timestamp 1676037725
transform 1 0 520076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5653
timestamp 1676037725
transform 1 0 521180 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5657
timestamp 1676037725
transform 1 0 521548 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5669
timestamp 1676037725
transform 1 0 522652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5681
timestamp 1676037725
transform 1 0 523756 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5685
timestamp 1676037725
transform 1 0 524124 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5697
timestamp 1676037725
transform 1 0 525228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5709
timestamp 1676037725
transform 1 0 526332 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5713
timestamp 1676037725
transform 1 0 526700 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5725
timestamp 1676037725
transform 1 0 527804 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1676037725
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1676037725
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1676037725
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1676037725
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1676037725
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1676037725
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1676037725
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_399
timestamp 1676037725
transform 1 0 37812 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_411
timestamp 1676037725
transform 1 0 38916 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_423
timestamp 1676037725
transform 1 0 40020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_435
timestamp 1676037725
transform 1 0 41124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1676037725
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1676037725
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1676037725
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1676037725
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1676037725
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1676037725
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1676037725
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1676037725
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1676037725
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1676037725
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1676037725
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1676037725
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1676037725
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1676037725
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1676037725
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1676037725
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_617
timestamp 1676037725
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_629
timestamp 1676037725
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_641
timestamp 1676037725
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_653
timestamp 1676037725
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 1676037725
transform 1 0 62284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1676037725
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1676037725
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_685
timestamp 1676037725
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_697
timestamp 1676037725
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_709
timestamp 1676037725
transform 1 0 66332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 1676037725
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1676037725
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_729
timestamp 1676037725
transform 1 0 68172 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_741
timestamp 1676037725
transform 1 0 69276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_753
timestamp 1676037725
transform 1 0 70380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_765
timestamp 1676037725
transform 1 0 71484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_777
timestamp 1676037725
transform 1 0 72588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 1676037725
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_785
timestamp 1676037725
transform 1 0 73324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_799
timestamp 1676037725
transform 1 0 74612 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_805
timestamp 1676037725
transform 1 0 75164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_817
timestamp 1676037725
transform 1 0 76268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_829
timestamp 1676037725
transform 1 0 77372 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_837
timestamp 1676037725
transform 1 0 78108 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_841
timestamp 1676037725
transform 1 0 78476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_853
timestamp 1676037725
transform 1 0 79580 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_865
timestamp 1676037725
transform 1 0 80684 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_877
timestamp 1676037725
transform 1 0 81788 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_889
timestamp 1676037725
transform 1 0 82892 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_895
timestamp 1676037725
transform 1 0 83444 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_897
timestamp 1676037725
transform 1 0 83628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_909
timestamp 1676037725
transform 1 0 84732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_921
timestamp 1676037725
transform 1 0 85836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_933
timestamp 1676037725
transform 1 0 86940 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_945
timestamp 1676037725
transform 1 0 88044 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_951
timestamp 1676037725
transform 1 0 88596 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_953
timestamp 1676037725
transform 1 0 88780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_965
timestamp 1676037725
transform 1 0 89884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_977
timestamp 1676037725
transform 1 0 90988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_989
timestamp 1676037725
transform 1 0 92092 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1001
timestamp 1676037725
transform 1 0 93196 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1007
timestamp 1676037725
transform 1 0 93748 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1009
timestamp 1676037725
transform 1 0 93932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1021
timestamp 1676037725
transform 1 0 95036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1033
timestamp 1676037725
transform 1 0 96140 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1045
timestamp 1676037725
transform 1 0 97244 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1057
timestamp 1676037725
transform 1 0 98348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1063
timestamp 1676037725
transform 1 0 98900 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1065
timestamp 1676037725
transform 1 0 99084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1077
timestamp 1676037725
transform 1 0 100188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1089
timestamp 1676037725
transform 1 0 101292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1101
timestamp 1676037725
transform 1 0 102396 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1113
timestamp 1676037725
transform 1 0 103500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1119
timestamp 1676037725
transform 1 0 104052 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1121
timestamp 1676037725
transform 1 0 104236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1133
timestamp 1676037725
transform 1 0 105340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1145
timestamp 1676037725
transform 1 0 106444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1157
timestamp 1676037725
transform 1 0 107548 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1165
timestamp 1676037725
transform 1 0 108284 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1173
timestamp 1676037725
transform 1 0 109020 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1177
timestamp 1676037725
transform 1 0 109388 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1189
timestamp 1676037725
transform 1 0 110492 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1201
timestamp 1676037725
transform 1 0 111596 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1205
timestamp 1676037725
transform 1 0 111964 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1208
timestamp 1676037725
transform 1 0 112240 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1214
timestamp 1676037725
transform 1 0 112792 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1217
timestamp 1676037725
transform 1 0 113068 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1230
timestamp 1676037725
transform 1 0 114264 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1233
timestamp 1676037725
transform 1 0 114540 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1237
timestamp 1676037725
transform 1 0 114908 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1247
timestamp 1676037725
transform 1 0 115828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1260
timestamp 1676037725
transform 1 0 117024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1273
timestamp 1676037725
transform 1 0 118220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1286
timestamp 1676037725
transform 1 0 119416 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1289
timestamp 1676037725
transform 1 0 119692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1293
timestamp 1676037725
transform 1 0 120060 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1303
timestamp 1676037725
transform 1 0 120980 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1316
timestamp 1676037725
transform 1 0 122176 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1329
timestamp 1676037725
transform 1 0 123372 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1342
timestamp 1676037725
transform 1 0 124568 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1345
timestamp 1676037725
transform 1 0 124844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1355
timestamp 1676037725
transform 1 0 125764 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1361
timestamp 1676037725
transform 1 0 126316 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1367
timestamp 1676037725
transform 1 0 126868 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1373
timestamp 1676037725
transform 1 0 127420 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1385
timestamp 1676037725
transform 1 0 128524 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1397
timestamp 1676037725
transform 1 0 129628 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1401
timestamp 1676037725
transform 1 0 129996 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1413
timestamp 1676037725
transform 1 0 131100 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1425
timestamp 1676037725
transform 1 0 132204 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1437
timestamp 1676037725
transform 1 0 133308 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1449
timestamp 1676037725
transform 1 0 134412 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1455
timestamp 1676037725
transform 1 0 134964 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1457
timestamp 1676037725
transform 1 0 135148 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1469
timestamp 1676037725
transform 1 0 136252 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1481
timestamp 1676037725
transform 1 0 137356 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1493
timestamp 1676037725
transform 1 0 138460 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1505
timestamp 1676037725
transform 1 0 139564 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1511
timestamp 1676037725
transform 1 0 140116 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1513
timestamp 1676037725
transform 1 0 140300 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1525
timestamp 1676037725
transform 1 0 141404 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1537
timestamp 1676037725
transform 1 0 142508 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1545
timestamp 1676037725
transform 1 0 143244 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1557
timestamp 1676037725
transform 1 0 144348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1565
timestamp 1676037725
transform 1 0 145084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1569
timestamp 1676037725
transform 1 0 145452 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1575
timestamp 1676037725
transform 1 0 146004 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1587
timestamp 1676037725
transform 1 0 147108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1599
timestamp 1676037725
transform 1 0 148212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1611
timestamp 1676037725
transform 1 0 149316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1623
timestamp 1676037725
transform 1 0 150420 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1625
timestamp 1676037725
transform 1 0 150604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1637
timestamp 1676037725
transform 1 0 151708 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1645
timestamp 1676037725
transform 1 0 152444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1657
timestamp 1676037725
transform 1 0 153548 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1669
timestamp 1676037725
transform 1 0 154652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1677
timestamp 1676037725
transform 1 0 155388 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1681
timestamp 1676037725
transform 1 0 155756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1693
timestamp 1676037725
transform 1 0 156860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1705
timestamp 1676037725
transform 1 0 157964 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1717
timestamp 1676037725
transform 1 0 159068 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1729
timestamp 1676037725
transform 1 0 160172 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1735
timestamp 1676037725
transform 1 0 160724 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1737
timestamp 1676037725
transform 1 0 160908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1749
timestamp 1676037725
transform 1 0 162012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1761
timestamp 1676037725
transform 1 0 163116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1775
timestamp 1676037725
transform 1 0 164404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1781
timestamp 1676037725
transform 1 0 164956 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1789
timestamp 1676037725
transform 1 0 165692 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1793
timestamp 1676037725
transform 1 0 166060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1805
timestamp 1676037725
transform 1 0 167164 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1813
timestamp 1676037725
transform 1 0 167900 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1816
timestamp 1676037725
transform 1 0 168176 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1829
timestamp 1676037725
transform 1 0 169372 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1841
timestamp 1676037725
transform 1 0 170476 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1847
timestamp 1676037725
transform 1 0 171028 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1849
timestamp 1676037725
transform 1 0 171212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1861
timestamp 1676037725
transform 1 0 172316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1873
timestamp 1676037725
transform 1 0 173420 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1885
timestamp 1676037725
transform 1 0 174524 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1897
timestamp 1676037725
transform 1 0 175628 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1903
timestamp 1676037725
transform 1 0 176180 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1905
timestamp 1676037725
transform 1 0 176364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1917
timestamp 1676037725
transform 1 0 177468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1929
timestamp 1676037725
transform 1 0 178572 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1941
timestamp 1676037725
transform 1 0 179676 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1953
timestamp 1676037725
transform 1 0 180780 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1959
timestamp 1676037725
transform 1 0 181332 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1961
timestamp 1676037725
transform 1 0 181516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1973
timestamp 1676037725
transform 1 0 182620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1985
timestamp 1676037725
transform 1 0 183724 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1997
timestamp 1676037725
transform 1 0 184828 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2009
timestamp 1676037725
transform 1 0 185932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2015
timestamp 1676037725
transform 1 0 186484 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2017
timestamp 1676037725
transform 1 0 186668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2029
timestamp 1676037725
transform 1 0 187772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2041
timestamp 1676037725
transform 1 0 188876 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2053
timestamp 1676037725
transform 1 0 189980 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2065
timestamp 1676037725
transform 1 0 191084 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2071
timestamp 1676037725
transform 1 0 191636 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2073
timestamp 1676037725
transform 1 0 191820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2085
timestamp 1676037725
transform 1 0 192924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2097
timestamp 1676037725
transform 1 0 194028 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2109
timestamp 1676037725
transform 1 0 195132 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2121
timestamp 1676037725
transform 1 0 196236 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2127
timestamp 1676037725
transform 1 0 196788 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2129
timestamp 1676037725
transform 1 0 196972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2141
timestamp 1676037725
transform 1 0 198076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2153
timestamp 1676037725
transform 1 0 199180 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2165
timestamp 1676037725
transform 1 0 200284 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_2177
timestamp 1676037725
transform 1 0 201388 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_2182
timestamp 1676037725
transform 1 0 201848 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_2185
timestamp 1676037725
transform 1 0 202124 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2196
timestamp 1676037725
transform 1 0 203136 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2208
timestamp 1676037725
transform 1 0 204240 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2223
timestamp 1676037725
transform 1 0 205620 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2229
timestamp 1676037725
transform 1 0 206172 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2235
timestamp 1676037725
transform 1 0 206724 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_2238
timestamp 1676037725
transform 1 0 207000 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_2241
timestamp 1676037725
transform 1 0 207276 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2252
timestamp 1676037725
transform 1 0 208288 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2258
timestamp 1676037725
transform 1 0 208840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2268
timestamp 1676037725
transform 1 0 209760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2281
timestamp 1676037725
transform 1 0 210956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_2294
timestamp 1676037725
transform 1 0 212152 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2297
timestamp 1676037725
transform 1 0 212428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2301
timestamp 1676037725
transform 1 0 212796 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2311
timestamp 1676037725
transform 1 0 213716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2324
timestamp 1676037725
transform 1 0 214912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2337
timestamp 1676037725
transform 1 0 216108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_2350
timestamp 1676037725
transform 1 0 217304 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2353
timestamp 1676037725
transform 1 0 217580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2357
timestamp 1676037725
transform 1 0 217948 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2360
timestamp 1676037725
transform 1 0 218224 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2373
timestamp 1676037725
transform 1 0 219420 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2386
timestamp 1676037725
transform 1 0 220616 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2392
timestamp 1676037725
transform 1 0 221168 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2398
timestamp 1676037725
transform 1 0 221720 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_2406
timestamp 1676037725
transform 1 0 222456 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2409
timestamp 1676037725
transform 1 0 222732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2421
timestamp 1676037725
transform 1 0 223836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2433
timestamp 1676037725
transform 1 0 224940 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2445
timestamp 1676037725
transform 1 0 226044 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2457
timestamp 1676037725
transform 1 0 227148 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2463
timestamp 1676037725
transform 1 0 227700 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2465
timestamp 1676037725
transform 1 0 227884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2477
timestamp 1676037725
transform 1 0 228988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2489
timestamp 1676037725
transform 1 0 230092 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2501
timestamp 1676037725
transform 1 0 231196 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2513
timestamp 1676037725
transform 1 0 232300 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2519
timestamp 1676037725
transform 1 0 232852 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2521
timestamp 1676037725
transform 1 0 233036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2533
timestamp 1676037725
transform 1 0 234140 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2545
timestamp 1676037725
transform 1 0 235244 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2557
timestamp 1676037725
transform 1 0 236348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2569
timestamp 1676037725
transform 1 0 237452 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2575
timestamp 1676037725
transform 1 0 238004 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2577
timestamp 1676037725
transform 1 0 238188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2589
timestamp 1676037725
transform 1 0 239292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2601
timestamp 1676037725
transform 1 0 240396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2613
timestamp 1676037725
transform 1 0 241500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2625
timestamp 1676037725
transform 1 0 242604 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2631
timestamp 1676037725
transform 1 0 243156 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2633
timestamp 1676037725
transform 1 0 243340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2645
timestamp 1676037725
transform 1 0 244444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2657
timestamp 1676037725
transform 1 0 245548 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2669
timestamp 1676037725
transform 1 0 246652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2677
timestamp 1676037725
transform 1 0 247388 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_2685
timestamp 1676037725
transform 1 0 248124 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2689
timestamp 1676037725
transform 1 0 248492 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2701
timestamp 1676037725
transform 1 0 249596 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2713
timestamp 1676037725
transform 1 0 250700 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2723
timestamp 1676037725
transform 1 0 251620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2735
timestamp 1676037725
transform 1 0 252724 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2743
timestamp 1676037725
transform 1 0 253460 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2745
timestamp 1676037725
transform 1 0 253644 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2751
timestamp 1676037725
transform 1 0 254196 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2763
timestamp 1676037725
transform 1 0 255300 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2775
timestamp 1676037725
transform 1 0 256404 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2787
timestamp 1676037725
transform 1 0 257508 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2799
timestamp 1676037725
transform 1 0 258612 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_2801
timestamp 1676037725
transform 1 0 258796 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2812
timestamp 1676037725
transform 1 0 259808 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2818
timestamp 1676037725
transform 1 0 260360 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2830
timestamp 1676037725
transform 1 0 261464 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2842
timestamp 1676037725
transform 1 0 262568 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_2854
timestamp 1676037725
transform 1 0 263672 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2857
timestamp 1676037725
transform 1 0 263948 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2869
timestamp 1676037725
transform 1 0 265052 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2881
timestamp 1676037725
transform 1 0 266156 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2893
timestamp 1676037725
transform 1 0 267260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2905
timestamp 1676037725
transform 1 0 268364 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2911
timestamp 1676037725
transform 1 0 268916 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2913
timestamp 1676037725
transform 1 0 269100 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2925
timestamp 1676037725
transform 1 0 270204 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2937
timestamp 1676037725
transform 1 0 271308 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2949
timestamp 1676037725
transform 1 0 272412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2961
timestamp 1676037725
transform 1 0 273516 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2967
timestamp 1676037725
transform 1 0 274068 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2969
timestamp 1676037725
transform 1 0 274252 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2981
timestamp 1676037725
transform 1 0 275356 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2993
timestamp 1676037725
transform 1 0 276460 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3005
timestamp 1676037725
transform 1 0 277564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3017
timestamp 1676037725
transform 1 0 278668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3023
timestamp 1676037725
transform 1 0 279220 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3025
timestamp 1676037725
transform 1 0 279404 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3037
timestamp 1676037725
transform 1 0 280508 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3049
timestamp 1676037725
transform 1 0 281612 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3061
timestamp 1676037725
transform 1 0 282716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3073
timestamp 1676037725
transform 1 0 283820 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3079
timestamp 1676037725
transform 1 0 284372 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3081
timestamp 1676037725
transform 1 0 284556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3093
timestamp 1676037725
transform 1 0 285660 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3105
timestamp 1676037725
transform 1 0 286764 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3117
timestamp 1676037725
transform 1 0 287868 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3129
timestamp 1676037725
transform 1 0 288972 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3135
timestamp 1676037725
transform 1 0 289524 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3137
timestamp 1676037725
transform 1 0 289708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3149
timestamp 1676037725
transform 1 0 290812 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3161
timestamp 1676037725
transform 1 0 291916 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3173
timestamp 1676037725
transform 1 0 293020 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3185
timestamp 1676037725
transform 1 0 294124 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3191
timestamp 1676037725
transform 1 0 294676 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3193
timestamp 1676037725
transform 1 0 294860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3207
timestamp 1676037725
transform 1 0 296148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3213
timestamp 1676037725
transform 1 0 296700 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3219
timestamp 1676037725
transform 1 0 297252 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3223
timestamp 1676037725
transform 1 0 297620 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3229
timestamp 1676037725
transform 1 0 298172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3235
timestamp 1676037725
transform 1 0 298724 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3243
timestamp 1676037725
transform 1 0 299460 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3246
timestamp 1676037725
transform 1 0 299736 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3249
timestamp 1676037725
transform 1 0 300012 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3257
timestamp 1676037725
transform 1 0 300748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3264
timestamp 1676037725
transform 1 0 301392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3270
timestamp 1676037725
transform 1 0 301944 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3278
timestamp 1676037725
transform 1 0 302680 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3285
timestamp 1676037725
transform 1 0 303324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3298
timestamp 1676037725
transform 1 0 304520 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3305
timestamp 1676037725
transform 1 0 305164 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3313
timestamp 1676037725
transform 1 0 305900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3323
timestamp 1676037725
transform 1 0 306820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3333
timestamp 1676037725
transform 1 0 307740 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3343
timestamp 1676037725
transform 1 0 308660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3353
timestamp 1676037725
transform 1 0 309580 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3359
timestamp 1676037725
transform 1 0 310132 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3361
timestamp 1676037725
transform 1 0 310316 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3369
timestamp 1676037725
transform 1 0 311052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3379
timestamp 1676037725
transform 1 0 311972 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3389
timestamp 1676037725
transform 1 0 312892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3395
timestamp 1676037725
transform 1 0 313444 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3403
timestamp 1676037725
transform 1 0 314180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3411
timestamp 1676037725
transform 1 0 314916 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3415
timestamp 1676037725
transform 1 0 315284 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3417
timestamp 1676037725
transform 1 0 315468 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3421
timestamp 1676037725
transform 1 0 315836 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3433
timestamp 1676037725
transform 1 0 316940 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3438
timestamp 1676037725
transform 1 0 317400 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3444
timestamp 1676037725
transform 1 0 317952 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3458
timestamp 1676037725
transform 1 0 319240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3464
timestamp 1676037725
transform 1 0 319792 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3473
timestamp 1676037725
transform 1 0 320620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3485
timestamp 1676037725
transform 1 0 321724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3497
timestamp 1676037725
transform 1 0 322828 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3505
timestamp 1676037725
transform 1 0 323564 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3508
timestamp 1676037725
transform 1 0 323840 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3516
timestamp 1676037725
transform 1 0 324576 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3520
timestamp 1676037725
transform 1 0 324944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3526
timestamp 1676037725
transform 1 0 325496 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3529
timestamp 1676037725
transform 1 0 325772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3541
timestamp 1676037725
transform 1 0 326876 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3553
timestamp 1676037725
transform 1 0 327980 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3565
timestamp 1676037725
transform 1 0 329084 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3577
timestamp 1676037725
transform 1 0 330188 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3583
timestamp 1676037725
transform 1 0 330740 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3585
timestamp 1676037725
transform 1 0 330924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3592
timestamp 1676037725
transform 1 0 331568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3598
timestamp 1676037725
transform 1 0 332120 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3604
timestamp 1676037725
transform 1 0 332672 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3616
timestamp 1676037725
transform 1 0 333776 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3628
timestamp 1676037725
transform 1 0 334880 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3641
timestamp 1676037725
transform 1 0 336076 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3653
timestamp 1676037725
transform 1 0 337180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3658
timestamp 1676037725
transform 1 0 337640 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3664
timestamp 1676037725
transform 1 0 338192 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3676
timestamp 1676037725
transform 1 0 339296 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3682
timestamp 1676037725
transform 1 0 339848 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3687
timestamp 1676037725
transform 1 0 340308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3693
timestamp 1676037725
transform 1 0 340860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3697
timestamp 1676037725
transform 1 0 341228 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3701
timestamp 1676037725
transform 1 0 341596 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3707
timestamp 1676037725
transform 1 0 342148 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3719
timestamp 1676037725
transform 1 0 343252 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3727
timestamp 1676037725
transform 1 0 343988 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3733
timestamp 1676037725
transform 1 0 344540 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3739
timestamp 1676037725
transform 1 0 345092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3745
timestamp 1676037725
transform 1 0 345644 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3751
timestamp 1676037725
transform 1 0 346196 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3753
timestamp 1676037725
transform 1 0 346380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3757
timestamp 1676037725
transform 1 0 346748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3769
timestamp 1676037725
transform 1 0 347852 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3779
timestamp 1676037725
transform 1 0 348772 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3793
timestamp 1676037725
transform 1 0 350060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3799
timestamp 1676037725
transform 1 0 350612 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3807
timestamp 1676037725
transform 1 0 351348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3809
timestamp 1676037725
transform 1 0 351532 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3817
timestamp 1676037725
transform 1 0 352268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3822
timestamp 1676037725
transform 1 0 352728 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3826
timestamp 1676037725
transform 1 0 353096 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3829
timestamp 1676037725
transform 1 0 353372 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3837
timestamp 1676037725
transform 1 0 354108 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3843
timestamp 1676037725
transform 1 0 354660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3855
timestamp 1676037725
transform 1 0 355764 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3861
timestamp 1676037725
transform 1 0 356316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3865
timestamp 1676037725
transform 1 0 356684 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3871
timestamp 1676037725
transform 1 0 357236 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3876
timestamp 1676037725
transform 1 0 357696 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3882
timestamp 1676037725
transform 1 0 358248 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3894
timestamp 1676037725
transform 1 0 359352 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3906
timestamp 1676037725
transform 1 0 360456 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3918
timestamp 1676037725
transform 1 0 361560 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3921
timestamp 1676037725
transform 1 0 361836 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3927
timestamp 1676037725
transform 1 0 362388 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3939
timestamp 1676037725
transform 1 0 363492 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3951
timestamp 1676037725
transform 1 0 364596 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3963
timestamp 1676037725
transform 1 0 365700 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3975
timestamp 1676037725
transform 1 0 366804 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3977
timestamp 1676037725
transform 1 0 366988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3989
timestamp 1676037725
transform 1 0 368092 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4001
timestamp 1676037725
transform 1 0 369196 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4013
timestamp 1676037725
transform 1 0 370300 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4025
timestamp 1676037725
transform 1 0 371404 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4031
timestamp 1676037725
transform 1 0 371956 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4033
timestamp 1676037725
transform 1 0 372140 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4045
timestamp 1676037725
transform 1 0 373244 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4057
timestamp 1676037725
transform 1 0 374348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4069
timestamp 1676037725
transform 1 0 375452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4081
timestamp 1676037725
transform 1 0 376556 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4087
timestamp 1676037725
transform 1 0 377108 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4089
timestamp 1676037725
transform 1 0 377292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4101
timestamp 1676037725
transform 1 0 378396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4113
timestamp 1676037725
transform 1 0 379500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_4125
timestamp 1676037725
transform 1 0 380604 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4129
timestamp 1676037725
transform 1 0 380972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_4141
timestamp 1676037725
transform 1 0 382076 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4145
timestamp 1676037725
transform 1 0 382444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4157
timestamp 1676037725
transform 1 0 383548 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4169
timestamp 1676037725
transform 1 0 384652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4181
timestamp 1676037725
transform 1 0 385756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4193
timestamp 1676037725
transform 1 0 386860 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4199
timestamp 1676037725
transform 1 0 387412 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4201
timestamp 1676037725
transform 1 0 387596 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4213
timestamp 1676037725
transform 1 0 388700 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_4225
timestamp 1676037725
transform 1 0 389804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_4235
timestamp 1676037725
transform 1 0 390724 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_4241
timestamp 1676037725
transform 1 0 391276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_4247
timestamp 1676037725
transform 1 0 391828 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4255
timestamp 1676037725
transform 1 0 392564 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_4257
timestamp 1676037725
transform 1 0 392748 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_4265
timestamp 1676037725
transform 1 0 393484 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4273
timestamp 1676037725
transform 1 0 394220 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_4283
timestamp 1676037725
transform 1 0 395140 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_4291
timestamp 1676037725
transform 1 0 395876 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_4295
timestamp 1676037725
transform 1 0 396244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4299
timestamp 1676037725
transform 1 0 396612 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4306
timestamp 1676037725
transform 1 0 397256 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_4313
timestamp 1676037725
transform 1 0 397900 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4317
timestamp 1676037725
transform 1 0 398268 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_4325
timestamp 1676037725
transform 1 0 399004 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_4333
timestamp 1676037725
transform 1 0 399740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4338
timestamp 1676037725
transform 1 0 400200 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4344
timestamp 1676037725
transform 1 0 400752 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4347
timestamp 1676037725
transform 1 0 401028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_4359
timestamp 1676037725
transform 1 0 402132 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4367
timestamp 1676037725
transform 1 0 402868 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4369
timestamp 1676037725
transform 1 0 403052 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4381
timestamp 1676037725
transform 1 0 404156 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4393
timestamp 1676037725
transform 1 0 405260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4405
timestamp 1676037725
transform 1 0 406364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4417
timestamp 1676037725
transform 1 0 407468 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4423
timestamp 1676037725
transform 1 0 408020 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_4425
timestamp 1676037725
transform 1 0 408204 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4429
timestamp 1676037725
transform 1 0 408572 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4441
timestamp 1676037725
transform 1 0 409676 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4453
timestamp 1676037725
transform 1 0 410780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4465
timestamp 1676037725
transform 1 0 411884 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_4477
timestamp 1676037725
transform 1 0 412988 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4481
timestamp 1676037725
transform 1 0 413356 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4493
timestamp 1676037725
transform 1 0 414460 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_4505
timestamp 1676037725
transform 1 0 415564 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4515
timestamp 1676037725
transform 1 0 416484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_4527
timestamp 1676037725
transform 1 0 417588 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4535
timestamp 1676037725
transform 1 0 418324 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4537
timestamp 1676037725
transform 1 0 418508 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4549
timestamp 1676037725
transform 1 0 419612 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4561
timestamp 1676037725
transform 1 0 420716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4573
timestamp 1676037725
transform 1 0 421820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4585
timestamp 1676037725
transform 1 0 422924 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4591
timestamp 1676037725
transform 1 0 423476 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4593
timestamp 1676037725
transform 1 0 423660 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4605
timestamp 1676037725
transform 1 0 424764 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4617
timestamp 1676037725
transform 1 0 425868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4629
timestamp 1676037725
transform 1 0 426972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4641
timestamp 1676037725
transform 1 0 428076 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4647
timestamp 1676037725
transform 1 0 428628 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4649
timestamp 1676037725
transform 1 0 428812 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4661
timestamp 1676037725
transform 1 0 429916 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4673
timestamp 1676037725
transform 1 0 431020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4685
timestamp 1676037725
transform 1 0 432124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4697
timestamp 1676037725
transform 1 0 433228 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4703
timestamp 1676037725
transform 1 0 433780 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_4705
timestamp 1676037725
transform 1 0 433964 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_4713
timestamp 1676037725
transform 1 0 434700 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_4717
timestamp 1676037725
transform 1 0 435068 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4727
timestamp 1676037725
transform 1 0 435988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4739
timestamp 1676037725
transform 1 0 437092 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_4751
timestamp 1676037725
transform 1 0 438196 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4759
timestamp 1676037725
transform 1 0 438932 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4761
timestamp 1676037725
transform 1 0 439116 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4773
timestamp 1676037725
transform 1 0 440220 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4785
timestamp 1676037725
transform 1 0 441324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4797
timestamp 1676037725
transform 1 0 442428 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4809
timestamp 1676037725
transform 1 0 443532 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4815
timestamp 1676037725
transform 1 0 444084 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4817
timestamp 1676037725
transform 1 0 444268 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4829
timestamp 1676037725
transform 1 0 445372 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4841
timestamp 1676037725
transform 1 0 446476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4853
timestamp 1676037725
transform 1 0 447580 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4865
timestamp 1676037725
transform 1 0 448684 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4871
timestamp 1676037725
transform 1 0 449236 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4873
timestamp 1676037725
transform 1 0 449420 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4885
timestamp 1676037725
transform 1 0 450524 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_4897
timestamp 1676037725
transform 1 0 451628 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_4911
timestamp 1676037725
transform 1 0 452916 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_4917
timestamp 1676037725
transform 1 0 453468 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_4925
timestamp 1676037725
transform 1 0 454204 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4929
timestamp 1676037725
transform 1 0 454572 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4941
timestamp 1676037725
transform 1 0 455676 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4953
timestamp 1676037725
transform 1 0 456780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4965
timestamp 1676037725
transform 1 0 457884 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4977
timestamp 1676037725
transform 1 0 458988 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4983
timestamp 1676037725
transform 1 0 459540 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4985
timestamp 1676037725
transform 1 0 459724 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4997
timestamp 1676037725
transform 1 0 460828 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5009
timestamp 1676037725
transform 1 0 461932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5021
timestamp 1676037725
transform 1 0 463036 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5033
timestamp 1676037725
transform 1 0 464140 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5039
timestamp 1676037725
transform 1 0 464692 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5041
timestamp 1676037725
transform 1 0 464876 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5053
timestamp 1676037725
transform 1 0 465980 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5065
timestamp 1676037725
transform 1 0 467084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5077
timestamp 1676037725
transform 1 0 468188 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5089
timestamp 1676037725
transform 1 0 469292 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5095
timestamp 1676037725
transform 1 0 469844 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5097
timestamp 1676037725
transform 1 0 470028 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5103
timestamp 1676037725
transform 1 0 470580 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5115
timestamp 1676037725
transform 1 0 471684 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5127
timestamp 1676037725
transform 1 0 472788 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5139
timestamp 1676037725
transform 1 0 473892 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5151
timestamp 1676037725
transform 1 0 474996 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5153
timestamp 1676037725
transform 1 0 475180 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5165
timestamp 1676037725
transform 1 0 476284 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5177
timestamp 1676037725
transform 1 0 477388 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5189
timestamp 1676037725
transform 1 0 478492 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5201
timestamp 1676037725
transform 1 0 479596 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5207
timestamp 1676037725
transform 1 0 480148 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5209
timestamp 1676037725
transform 1 0 480332 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5221
timestamp 1676037725
transform 1 0 481436 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5233
timestamp 1676037725
transform 1 0 482540 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5245
timestamp 1676037725
transform 1 0 483644 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5257
timestamp 1676037725
transform 1 0 484748 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5263
timestamp 1676037725
transform 1 0 485300 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5265
timestamp 1676037725
transform 1 0 485484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5277
timestamp 1676037725
transform 1 0 486588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5289
timestamp 1676037725
transform 1 0 487692 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5301
timestamp 1676037725
transform 1 0 488796 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5313
timestamp 1676037725
transform 1 0 489900 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5319
timestamp 1676037725
transform 1 0 490452 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5321
timestamp 1676037725
transform 1 0 490636 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5333
timestamp 1676037725
transform 1 0 491740 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5345
timestamp 1676037725
transform 1 0 492844 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5357
timestamp 1676037725
transform 1 0 493948 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5369
timestamp 1676037725
transform 1 0 495052 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5375
timestamp 1676037725
transform 1 0 495604 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5377
timestamp 1676037725
transform 1 0 495788 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5389
timestamp 1676037725
transform 1 0 496892 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5401
timestamp 1676037725
transform 1 0 497996 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5413
timestamp 1676037725
transform 1 0 499100 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5425
timestamp 1676037725
transform 1 0 500204 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5431
timestamp 1676037725
transform 1 0 500756 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5433
timestamp 1676037725
transform 1 0 500940 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5445
timestamp 1676037725
transform 1 0 502044 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5457
timestamp 1676037725
transform 1 0 503148 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5469
timestamp 1676037725
transform 1 0 504252 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5481
timestamp 1676037725
transform 1 0 505356 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5487
timestamp 1676037725
transform 1 0 505908 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5489
timestamp 1676037725
transform 1 0 506092 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5501
timestamp 1676037725
transform 1 0 507196 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5513
timestamp 1676037725
transform 1 0 508300 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5525
timestamp 1676037725
transform 1 0 509404 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5537
timestamp 1676037725
transform 1 0 510508 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5543
timestamp 1676037725
transform 1 0 511060 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5545
timestamp 1676037725
transform 1 0 511244 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5557
timestamp 1676037725
transform 1 0 512348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5569
timestamp 1676037725
transform 1 0 513452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5581
timestamp 1676037725
transform 1 0 514556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5593
timestamp 1676037725
transform 1 0 515660 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5599
timestamp 1676037725
transform 1 0 516212 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5601
timestamp 1676037725
transform 1 0 516396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5613
timestamp 1676037725
transform 1 0 517500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5625
timestamp 1676037725
transform 1 0 518604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5637
timestamp 1676037725
transform 1 0 519708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5649
timestamp 1676037725
transform 1 0 520812 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5655
timestamp 1676037725
transform 1 0 521364 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5657
timestamp 1676037725
transform 1 0 521548 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5669
timestamp 1676037725
transform 1 0 522652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5681
timestamp 1676037725
transform 1 0 523756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5693
timestamp 1676037725
transform 1 0 524860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5705
timestamp 1676037725
transform 1 0 525964 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5711
timestamp 1676037725
transform 1 0 526516 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5713
timestamp 1676037725
transform 1 0 526700 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_5725
timestamp 1676037725
transform 1 0 527804 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1676037725
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1676037725
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1676037725
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1676037725
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1676037725
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1676037725
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1676037725
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1676037725
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1676037725
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1676037725
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1676037725
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1676037725
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1676037725
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1676037725
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1676037725
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1676037725
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1676037725
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1676037725
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1676037725
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1676037725
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1676037725
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1676037725
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1676037725
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_625
timestamp 1676037725
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1676037725
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1676037725
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1676037725
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1676037725
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1676037725
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1676037725
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 1676037725
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1676037725
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1676037725
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1676037725
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1676037725
transform 1 0 67804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_737
timestamp 1676037725
transform 1 0 68908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 1676037725
transform 1 0 70012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1676037725
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_757
timestamp 1676037725
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_769
timestamp 1676037725
transform 1 0 71852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_781
timestamp 1676037725
transform 1 0 72956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_793
timestamp 1676037725
transform 1 0 74060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 1676037725
transform 1 0 75164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 1676037725
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_813
timestamp 1676037725
transform 1 0 75900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_825
timestamp 1676037725
transform 1 0 77004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_837
timestamp 1676037725
transform 1 0 78108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_849
timestamp 1676037725
transform 1 0 79212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_861
timestamp 1676037725
transform 1 0 80316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_867
timestamp 1676037725
transform 1 0 80868 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_869
timestamp 1676037725
transform 1 0 81052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_881
timestamp 1676037725
transform 1 0 82156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_893
timestamp 1676037725
transform 1 0 83260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_905
timestamp 1676037725
transform 1 0 84364 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_917
timestamp 1676037725
transform 1 0 85468 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_923
timestamp 1676037725
transform 1 0 86020 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_925
timestamp 1676037725
transform 1 0 86204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_937
timestamp 1676037725
transform 1 0 87308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_949
timestamp 1676037725
transform 1 0 88412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_961
timestamp 1676037725
transform 1 0 89516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_973
timestamp 1676037725
transform 1 0 90620 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_979
timestamp 1676037725
transform 1 0 91172 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_981
timestamp 1676037725
transform 1 0 91356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_993
timestamp 1676037725
transform 1 0 92460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1005
timestamp 1676037725
transform 1 0 93564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1017
timestamp 1676037725
transform 1 0 94668 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1029
timestamp 1676037725
transform 1 0 95772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1035
timestamp 1676037725
transform 1 0 96324 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1037
timestamp 1676037725
transform 1 0 96508 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1049
timestamp 1676037725
transform 1 0 97612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1061
timestamp 1676037725
transform 1 0 98716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1073
timestamp 1676037725
transform 1 0 99820 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1085
timestamp 1676037725
transform 1 0 100924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1091
timestamp 1676037725
transform 1 0 101476 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1093
timestamp 1676037725
transform 1 0 101660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1105
timestamp 1676037725
transform 1 0 102764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1117
timestamp 1676037725
transform 1 0 103868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1129
timestamp 1676037725
transform 1 0 104972 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1141
timestamp 1676037725
transform 1 0 106076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1147
timestamp 1676037725
transform 1 0 106628 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1149
timestamp 1676037725
transform 1 0 106812 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1161
timestamp 1676037725
transform 1 0 107916 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1173
timestamp 1676037725
transform 1 0 109020 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1185
timestamp 1676037725
transform 1 0 110124 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1197
timestamp 1676037725
transform 1 0 111228 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1203
timestamp 1676037725
transform 1 0 111780 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1205
timestamp 1676037725
transform 1 0 111964 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1217
timestamp 1676037725
transform 1 0 113068 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1223
timestamp 1676037725
transform 1 0 113620 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1226
timestamp 1676037725
transform 1 0 113896 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1232
timestamp 1676037725
transform 1 0 114448 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1245
timestamp 1676037725
transform 1 0 115644 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1258
timestamp 1676037725
transform 1 0 116840 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1261
timestamp 1676037725
transform 1 0 117116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1274
timestamp 1676037725
transform 1 0 118312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1287
timestamp 1676037725
transform 1 0 119508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1300
timestamp 1676037725
transform 1 0 120704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1304
timestamp 1676037725
transform 1 0 121072 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1314
timestamp 1676037725
transform 1 0 121992 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1317
timestamp 1676037725
transform 1 0 122268 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1321
timestamp 1676037725
transform 1 0 122636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1325
timestamp 1676037725
transform 1 0 123004 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1328
timestamp 1676037725
transform 1 0 123280 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1341
timestamp 1676037725
transform 1 0 124476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1351
timestamp 1676037725
transform 1 0 125396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1357
timestamp 1676037725
transform 1 0 125948 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1363
timestamp 1676037725
transform 1 0 126500 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1371
timestamp 1676037725
transform 1 0 127236 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1373
timestamp 1676037725
transform 1 0 127420 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1385
timestamp 1676037725
transform 1 0 128524 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1397
timestamp 1676037725
transform 1 0 129628 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1409
timestamp 1676037725
transform 1 0 130732 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1421
timestamp 1676037725
transform 1 0 131836 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1427
timestamp 1676037725
transform 1 0 132388 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1429
timestamp 1676037725
transform 1 0 132572 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1441
timestamp 1676037725
transform 1 0 133676 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1453
timestamp 1676037725
transform 1 0 134780 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1465
timestamp 1676037725
transform 1 0 135884 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1477
timestamp 1676037725
transform 1 0 136988 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1483
timestamp 1676037725
transform 1 0 137540 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1485
timestamp 1676037725
transform 1 0 137724 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1497
timestamp 1676037725
transform 1 0 138828 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1509
timestamp 1676037725
transform 1 0 139932 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1521
timestamp 1676037725
transform 1 0 141036 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1533
timestamp 1676037725
transform 1 0 142140 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1539
timestamp 1676037725
transform 1 0 142692 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1541
timestamp 1676037725
transform 1 0 142876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1553
timestamp 1676037725
transform 1 0 143980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1565
timestamp 1676037725
transform 1 0 145084 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1577
timestamp 1676037725
transform 1 0 146188 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1589
timestamp 1676037725
transform 1 0 147292 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1595
timestamp 1676037725
transform 1 0 147844 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1597
timestamp 1676037725
transform 1 0 148028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1609
timestamp 1676037725
transform 1 0 149132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1621
timestamp 1676037725
transform 1 0 150236 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1633
timestamp 1676037725
transform 1 0 151340 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1645
timestamp 1676037725
transform 1 0 152444 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1651
timestamp 1676037725
transform 1 0 152996 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1653
timestamp 1676037725
transform 1 0 153180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1665
timestamp 1676037725
transform 1 0 154284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1677
timestamp 1676037725
transform 1 0 155388 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1689
timestamp 1676037725
transform 1 0 156492 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1701
timestamp 1676037725
transform 1 0 157596 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1707
timestamp 1676037725
transform 1 0 158148 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1709
timestamp 1676037725
transform 1 0 158332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1721
timestamp 1676037725
transform 1 0 159436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1733
timestamp 1676037725
transform 1 0 160540 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1745
timestamp 1676037725
transform 1 0 161644 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1757
timestamp 1676037725
transform 1 0 162748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1763
timestamp 1676037725
transform 1 0 163300 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1765
timestamp 1676037725
transform 1 0 163484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1777
timestamp 1676037725
transform 1 0 164588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1789
timestamp 1676037725
transform 1 0 165692 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1801
timestamp 1676037725
transform 1 0 166796 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1813
timestamp 1676037725
transform 1 0 167900 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1819
timestamp 1676037725
transform 1 0 168452 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1821
timestamp 1676037725
transform 1 0 168636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1833
timestamp 1676037725
transform 1 0 169740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1845
timestamp 1676037725
transform 1 0 170844 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1857
timestamp 1676037725
transform 1 0 171948 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1869
timestamp 1676037725
transform 1 0 173052 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1875
timestamp 1676037725
transform 1 0 173604 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1877
timestamp 1676037725
transform 1 0 173788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1889
timestamp 1676037725
transform 1 0 174892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1901
timestamp 1676037725
transform 1 0 175996 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1913
timestamp 1676037725
transform 1 0 177100 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1925
timestamp 1676037725
transform 1 0 178204 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1931
timestamp 1676037725
transform 1 0 178756 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1933
timestamp 1676037725
transform 1 0 178940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1945
timestamp 1676037725
transform 1 0 180044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1957
timestamp 1676037725
transform 1 0 181148 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1969
timestamp 1676037725
transform 1 0 182252 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1981
timestamp 1676037725
transform 1 0 183356 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1987
timestamp 1676037725
transform 1 0 183908 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1989
timestamp 1676037725
transform 1 0 184092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2001
timestamp 1676037725
transform 1 0 185196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2013
timestamp 1676037725
transform 1 0 186300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2025
timestamp 1676037725
transform 1 0 187404 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2037
timestamp 1676037725
transform 1 0 188508 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2043
timestamp 1676037725
transform 1 0 189060 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2045
timestamp 1676037725
transform 1 0 189244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2057
timestamp 1676037725
transform 1 0 190348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2069
timestamp 1676037725
transform 1 0 191452 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2081
timestamp 1676037725
transform 1 0 192556 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2093
timestamp 1676037725
transform 1 0 193660 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2099
timestamp 1676037725
transform 1 0 194212 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2101
timestamp 1676037725
transform 1 0 194396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2113
timestamp 1676037725
transform 1 0 195500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2125
timestamp 1676037725
transform 1 0 196604 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2137
timestamp 1676037725
transform 1 0 197708 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2149
timestamp 1676037725
transform 1 0 198812 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2155
timestamp 1676037725
transform 1 0 199364 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2157
timestamp 1676037725
transform 1 0 199548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2169
timestamp 1676037725
transform 1 0 200652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2181
timestamp 1676037725
transform 1 0 201756 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2193
timestamp 1676037725
transform 1 0 202860 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2205
timestamp 1676037725
transform 1 0 203964 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2211
timestamp 1676037725
transform 1 0 204516 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2213
timestamp 1676037725
transform 1 0 204700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2225
timestamp 1676037725
transform 1 0 205804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2237
timestamp 1676037725
transform 1 0 206908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_2249
timestamp 1676037725
transform 1 0 208012 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_2253
timestamp 1676037725
transform 1 0 208380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_2266
timestamp 1676037725
transform 1 0 209576 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_2269
timestamp 1676037725
transform 1 0 209852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2273
timestamp 1676037725
transform 1 0 210220 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_2283
timestamp 1676037725
transform 1 0 211140 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_2296
timestamp 1676037725
transform 1 0 212336 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_2309
timestamp 1676037725
transform 1 0 213532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_2322
timestamp 1676037725
transform 1 0 214728 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_2325
timestamp 1676037725
transform 1 0 215004 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_2336
timestamp 1676037725
transform 1 0 216016 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_2349
timestamp 1676037725
transform 1 0 217212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_2362
timestamp 1676037725
transform 1 0 218408 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_2375
timestamp 1676037725
transform 1 0 219604 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2379
timestamp 1676037725
transform 1 0 219972 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_2381
timestamp 1676037725
transform 1 0 220156 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2385
timestamp 1676037725
transform 1 0 220524 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2397
timestamp 1676037725
transform 1 0 221628 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2409
timestamp 1676037725
transform 1 0 222732 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2421
timestamp 1676037725
transform 1 0 223836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_2433
timestamp 1676037725
transform 1 0 224940 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2437
timestamp 1676037725
transform 1 0 225308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2449
timestamp 1676037725
transform 1 0 226412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2461
timestamp 1676037725
transform 1 0 227516 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2473
timestamp 1676037725
transform 1 0 228620 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2485
timestamp 1676037725
transform 1 0 229724 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2491
timestamp 1676037725
transform 1 0 230276 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2493
timestamp 1676037725
transform 1 0 230460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2505
timestamp 1676037725
transform 1 0 231564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2517
timestamp 1676037725
transform 1 0 232668 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2529
timestamp 1676037725
transform 1 0 233772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2541
timestamp 1676037725
transform 1 0 234876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2547
timestamp 1676037725
transform 1 0 235428 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2549
timestamp 1676037725
transform 1 0 235612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2561
timestamp 1676037725
transform 1 0 236716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2573
timestamp 1676037725
transform 1 0 237820 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2585
timestamp 1676037725
transform 1 0 238924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2597
timestamp 1676037725
transform 1 0 240028 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2603
timestamp 1676037725
transform 1 0 240580 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2605
timestamp 1676037725
transform 1 0 240764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2617
timestamp 1676037725
transform 1 0 241868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2629
timestamp 1676037725
transform 1 0 242972 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2641
timestamp 1676037725
transform 1 0 244076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2653
timestamp 1676037725
transform 1 0 245180 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2659
timestamp 1676037725
transform 1 0 245732 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2661
timestamp 1676037725
transform 1 0 245916 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2673
timestamp 1676037725
transform 1 0 247020 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2685
timestamp 1676037725
transform 1 0 248124 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2697
timestamp 1676037725
transform 1 0 249228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2709
timestamp 1676037725
transform 1 0 250332 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2715
timestamp 1676037725
transform 1 0 250884 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2717
timestamp 1676037725
transform 1 0 251068 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2729
timestamp 1676037725
transform 1 0 252172 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2741
timestamp 1676037725
transform 1 0 253276 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2753
timestamp 1676037725
transform 1 0 254380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2765
timestamp 1676037725
transform 1 0 255484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2771
timestamp 1676037725
transform 1 0 256036 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2773
timestamp 1676037725
transform 1 0 256220 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2785
timestamp 1676037725
transform 1 0 257324 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2797
timestamp 1676037725
transform 1 0 258428 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2809
timestamp 1676037725
transform 1 0 259532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2821
timestamp 1676037725
transform 1 0 260636 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2827
timestamp 1676037725
transform 1 0 261188 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2829
timestamp 1676037725
transform 1 0 261372 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2841
timestamp 1676037725
transform 1 0 262476 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2853
timestamp 1676037725
transform 1 0 263580 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2865
timestamp 1676037725
transform 1 0 264684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2877
timestamp 1676037725
transform 1 0 265788 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2883
timestamp 1676037725
transform 1 0 266340 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2885
timestamp 1676037725
transform 1 0 266524 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2897
timestamp 1676037725
transform 1 0 267628 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2909
timestamp 1676037725
transform 1 0 268732 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2921
timestamp 1676037725
transform 1 0 269836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2933
timestamp 1676037725
transform 1 0 270940 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2939
timestamp 1676037725
transform 1 0 271492 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2941
timestamp 1676037725
transform 1 0 271676 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2953
timestamp 1676037725
transform 1 0 272780 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2965
timestamp 1676037725
transform 1 0 273884 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2977
timestamp 1676037725
transform 1 0 274988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2989
timestamp 1676037725
transform 1 0 276092 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2995
timestamp 1676037725
transform 1 0 276644 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2997
timestamp 1676037725
transform 1 0 276828 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3009
timestamp 1676037725
transform 1 0 277932 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3021
timestamp 1676037725
transform 1 0 279036 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3033
timestamp 1676037725
transform 1 0 280140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3045
timestamp 1676037725
transform 1 0 281244 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3051
timestamp 1676037725
transform 1 0 281796 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3053
timestamp 1676037725
transform 1 0 281980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3065
timestamp 1676037725
transform 1 0 283084 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3077
timestamp 1676037725
transform 1 0 284188 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3089
timestamp 1676037725
transform 1 0 285292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3101
timestamp 1676037725
transform 1 0 286396 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3107
timestamp 1676037725
transform 1 0 286948 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3109
timestamp 1676037725
transform 1 0 287132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3121
timestamp 1676037725
transform 1 0 288236 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3133
timestamp 1676037725
transform 1 0 289340 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3145
timestamp 1676037725
transform 1 0 290444 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3157
timestamp 1676037725
transform 1 0 291548 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3163
timestamp 1676037725
transform 1 0 292100 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3165
timestamp 1676037725
transform 1 0 292284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3177
timestamp 1676037725
transform 1 0 293388 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3189
timestamp 1676037725
transform 1 0 294492 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3201
timestamp 1676037725
transform 1 0 295596 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3213
timestamp 1676037725
transform 1 0 296700 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3219
timestamp 1676037725
transform 1 0 297252 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3221
timestamp 1676037725
transform 1 0 297436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3233
timestamp 1676037725
transform 1 0 298540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3245
timestamp 1676037725
transform 1 0 299644 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3251
timestamp 1676037725
transform 1 0 300196 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3259
timestamp 1676037725
transform 1 0 300932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3271
timestamp 1676037725
transform 1 0 302036 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3275
timestamp 1676037725
transform 1 0 302404 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3277
timestamp 1676037725
transform 1 0 302588 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3281
timestamp 1676037725
transform 1 0 302956 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3287
timestamp 1676037725
transform 1 0 303508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3300
timestamp 1676037725
transform 1 0 304704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3310
timestamp 1676037725
transform 1 0 305624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3320
timestamp 1676037725
transform 1 0 306544 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3330
timestamp 1676037725
transform 1 0 307464 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3333
timestamp 1676037725
transform 1 0 307740 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3341
timestamp 1676037725
transform 1 0 308476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3351
timestamp 1676037725
transform 1 0 309396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3361
timestamp 1676037725
transform 1 0 310316 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3371
timestamp 1676037725
transform 1 0 311236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3377
timestamp 1676037725
transform 1 0 311788 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3383
timestamp 1676037725
transform 1 0 312340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3387
timestamp 1676037725
transform 1 0 312708 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3389
timestamp 1676037725
transform 1 0 312892 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3393
timestamp 1676037725
transform 1 0 313260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3405
timestamp 1676037725
transform 1 0 314364 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3417
timestamp 1676037725
transform 1 0 315468 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3429
timestamp 1676037725
transform 1 0 316572 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3441
timestamp 1676037725
transform 1 0 317676 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3445
timestamp 1676037725
transform 1 0 318044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3457
timestamp 1676037725
transform 1 0 319148 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3469
timestamp 1676037725
transform 1 0 320252 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3481
timestamp 1676037725
transform 1 0 321356 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3493
timestamp 1676037725
transform 1 0 322460 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3499
timestamp 1676037725
transform 1 0 323012 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3501
timestamp 1676037725
transform 1 0 323196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3513
timestamp 1676037725
transform 1 0 324300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3525
timestamp 1676037725
transform 1 0 325404 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3537
timestamp 1676037725
transform 1 0 326508 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3549
timestamp 1676037725
transform 1 0 327612 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3555
timestamp 1676037725
transform 1 0 328164 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3557
timestamp 1676037725
transform 1 0 328348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3569
timestamp 1676037725
transform 1 0 329452 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3581
timestamp 1676037725
transform 1 0 330556 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3593
timestamp 1676037725
transform 1 0 331660 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3605
timestamp 1676037725
transform 1 0 332764 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3611
timestamp 1676037725
transform 1 0 333316 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3613
timestamp 1676037725
transform 1 0 333500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3625
timestamp 1676037725
transform 1 0 334604 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3637
timestamp 1676037725
transform 1 0 335708 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3649
timestamp 1676037725
transform 1 0 336812 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3661
timestamp 1676037725
transform 1 0 337916 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3667
timestamp 1676037725
transform 1 0 338468 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3669
timestamp 1676037725
transform 1 0 338652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3681
timestamp 1676037725
transform 1 0 339756 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3693
timestamp 1676037725
transform 1 0 340860 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3705
timestamp 1676037725
transform 1 0 341964 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3717
timestamp 1676037725
transform 1 0 343068 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3723
timestamp 1676037725
transform 1 0 343620 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3725
timestamp 1676037725
transform 1 0 343804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3737
timestamp 1676037725
transform 1 0 344908 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3749
timestamp 1676037725
transform 1 0 346012 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3761
timestamp 1676037725
transform 1 0 347116 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3773
timestamp 1676037725
transform 1 0 348220 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3779
timestamp 1676037725
transform 1 0 348772 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3781
timestamp 1676037725
transform 1 0 348956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3793
timestamp 1676037725
transform 1 0 350060 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3805
timestamp 1676037725
transform 1 0 351164 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3817
timestamp 1676037725
transform 1 0 352268 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3829
timestamp 1676037725
transform 1 0 353372 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3835
timestamp 1676037725
transform 1 0 353924 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3837
timestamp 1676037725
transform 1 0 354108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3849
timestamp 1676037725
transform 1 0 355212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3861
timestamp 1676037725
transform 1 0 356316 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3869
timestamp 1676037725
transform 1 0 357052 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3872
timestamp 1676037725
transform 1 0 357328 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3884
timestamp 1676037725
transform 1 0 358432 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3893
timestamp 1676037725
transform 1 0 359260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3905
timestamp 1676037725
transform 1 0 360364 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3917
timestamp 1676037725
transform 1 0 361468 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3929
timestamp 1676037725
transform 1 0 362572 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3941
timestamp 1676037725
transform 1 0 363676 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3947
timestamp 1676037725
transform 1 0 364228 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3949
timestamp 1676037725
transform 1 0 364412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3961
timestamp 1676037725
transform 1 0 365516 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3973
timestamp 1676037725
transform 1 0 366620 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3985
timestamp 1676037725
transform 1 0 367724 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3997
timestamp 1676037725
transform 1 0 368828 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4003
timestamp 1676037725
transform 1 0 369380 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4005
timestamp 1676037725
transform 1 0 369564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4017
timestamp 1676037725
transform 1 0 370668 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4029
timestamp 1676037725
transform 1 0 371772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4041
timestamp 1676037725
transform 1 0 372876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4053
timestamp 1676037725
transform 1 0 373980 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4059
timestamp 1676037725
transform 1 0 374532 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4061
timestamp 1676037725
transform 1 0 374716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4073
timestamp 1676037725
transform 1 0 375820 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4085
timestamp 1676037725
transform 1 0 376924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4097
timestamp 1676037725
transform 1 0 378028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4109
timestamp 1676037725
transform 1 0 379132 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4115
timestamp 1676037725
transform 1 0 379684 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4117
timestamp 1676037725
transform 1 0 379868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4129
timestamp 1676037725
transform 1 0 380972 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4141
timestamp 1676037725
transform 1 0 382076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4153
timestamp 1676037725
transform 1 0 383180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4165
timestamp 1676037725
transform 1 0 384284 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4171
timestamp 1676037725
transform 1 0 384836 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4173
timestamp 1676037725
transform 1 0 385020 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4185
timestamp 1676037725
transform 1 0 386124 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4197
timestamp 1676037725
transform 1 0 387228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4209
timestamp 1676037725
transform 1 0 388332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4221
timestamp 1676037725
transform 1 0 389436 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4227
timestamp 1676037725
transform 1 0 389988 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4229
timestamp 1676037725
transform 1 0 390172 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4241
timestamp 1676037725
transform 1 0 391276 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4253
timestamp 1676037725
transform 1 0 392380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_4267
timestamp 1676037725
transform 1 0 393668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4271
timestamp 1676037725
transform 1 0 394036 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_4274
timestamp 1676037725
transform 1 0 394312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_4280
timestamp 1676037725
transform 1 0 394864 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4285
timestamp 1676037725
transform 1 0 395324 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_4297
timestamp 1676037725
transform 1 0 396428 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4301
timestamp 1676037725
transform 1 0 396796 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4313
timestamp 1676037725
transform 1 0 397900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4325
timestamp 1676037725
transform 1 0 399004 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_4337
timestamp 1676037725
transform 1 0 400108 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4341
timestamp 1676037725
transform 1 0 400476 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4353
timestamp 1676037725
transform 1 0 401580 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4365
timestamp 1676037725
transform 1 0 402684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4377
timestamp 1676037725
transform 1 0 403788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4389
timestamp 1676037725
transform 1 0 404892 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4395
timestamp 1676037725
transform 1 0 405444 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4397
timestamp 1676037725
transform 1 0 405628 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4409
timestamp 1676037725
transform 1 0 406732 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4421
timestamp 1676037725
transform 1 0 407836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4433
timestamp 1676037725
transform 1 0 408940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4445
timestamp 1676037725
transform 1 0 410044 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4451
timestamp 1676037725
transform 1 0 410596 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4453
timestamp 1676037725
transform 1 0 410780 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4465
timestamp 1676037725
transform 1 0 411884 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4477
timestamp 1676037725
transform 1 0 412988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4489
timestamp 1676037725
transform 1 0 414092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4501
timestamp 1676037725
transform 1 0 415196 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4507
timestamp 1676037725
transform 1 0 415748 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4509
timestamp 1676037725
transform 1 0 415932 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4521
timestamp 1676037725
transform 1 0 417036 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4533
timestamp 1676037725
transform 1 0 418140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4545
timestamp 1676037725
transform 1 0 419244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4557
timestamp 1676037725
transform 1 0 420348 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4563
timestamp 1676037725
transform 1 0 420900 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4565
timestamp 1676037725
transform 1 0 421084 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4577
timestamp 1676037725
transform 1 0 422188 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4589
timestamp 1676037725
transform 1 0 423292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4601
timestamp 1676037725
transform 1 0 424396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4613
timestamp 1676037725
transform 1 0 425500 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4619
timestamp 1676037725
transform 1 0 426052 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4621
timestamp 1676037725
transform 1 0 426236 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4633
timestamp 1676037725
transform 1 0 427340 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4645
timestamp 1676037725
transform 1 0 428444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4657
timestamp 1676037725
transform 1 0 429548 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4669
timestamp 1676037725
transform 1 0 430652 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4675
timestamp 1676037725
transform 1 0 431204 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4677
timestamp 1676037725
transform 1 0 431388 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4689
timestamp 1676037725
transform 1 0 432492 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4701
timestamp 1676037725
transform 1 0 433596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4713
timestamp 1676037725
transform 1 0 434700 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4725
timestamp 1676037725
transform 1 0 435804 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4731
timestamp 1676037725
transform 1 0 436356 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4733
timestamp 1676037725
transform 1 0 436540 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4745
timestamp 1676037725
transform 1 0 437644 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4757
timestamp 1676037725
transform 1 0 438748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4769
timestamp 1676037725
transform 1 0 439852 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4781
timestamp 1676037725
transform 1 0 440956 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4787
timestamp 1676037725
transform 1 0 441508 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4789
timestamp 1676037725
transform 1 0 441692 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4801
timestamp 1676037725
transform 1 0 442796 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4813
timestamp 1676037725
transform 1 0 443900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4825
timestamp 1676037725
transform 1 0 445004 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4837
timestamp 1676037725
transform 1 0 446108 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4843
timestamp 1676037725
transform 1 0 446660 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4845
timestamp 1676037725
transform 1 0 446844 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4857
timestamp 1676037725
transform 1 0 447948 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4869
timestamp 1676037725
transform 1 0 449052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4881
timestamp 1676037725
transform 1 0 450156 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4893
timestamp 1676037725
transform 1 0 451260 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4899
timestamp 1676037725
transform 1 0 451812 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4901
timestamp 1676037725
transform 1 0 451996 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4913
timestamp 1676037725
transform 1 0 453100 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4925
timestamp 1676037725
transform 1 0 454204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4937
timestamp 1676037725
transform 1 0 455308 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4949
timestamp 1676037725
transform 1 0 456412 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4955
timestamp 1676037725
transform 1 0 456964 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4957
timestamp 1676037725
transform 1 0 457148 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4969
timestamp 1676037725
transform 1 0 458252 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4981
timestamp 1676037725
transform 1 0 459356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4993
timestamp 1676037725
transform 1 0 460460 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5005
timestamp 1676037725
transform 1 0 461564 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5011
timestamp 1676037725
transform 1 0 462116 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5013
timestamp 1676037725
transform 1 0 462300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5025
timestamp 1676037725
transform 1 0 463404 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5037
timestamp 1676037725
transform 1 0 464508 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5049
timestamp 1676037725
transform 1 0 465612 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5061
timestamp 1676037725
transform 1 0 466716 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5067
timestamp 1676037725
transform 1 0 467268 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5069
timestamp 1676037725
transform 1 0 467452 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5081
timestamp 1676037725
transform 1 0 468556 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5093
timestamp 1676037725
transform 1 0 469660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5105
timestamp 1676037725
transform 1 0 470764 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5117
timestamp 1676037725
transform 1 0 471868 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5123
timestamp 1676037725
transform 1 0 472420 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5125
timestamp 1676037725
transform 1 0 472604 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5137
timestamp 1676037725
transform 1 0 473708 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5149
timestamp 1676037725
transform 1 0 474812 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5161
timestamp 1676037725
transform 1 0 475916 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5173
timestamp 1676037725
transform 1 0 477020 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5179
timestamp 1676037725
transform 1 0 477572 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5181
timestamp 1676037725
transform 1 0 477756 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5193
timestamp 1676037725
transform 1 0 478860 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5205
timestamp 1676037725
transform 1 0 479964 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5217
timestamp 1676037725
transform 1 0 481068 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5229
timestamp 1676037725
transform 1 0 482172 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5235
timestamp 1676037725
transform 1 0 482724 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5237
timestamp 1676037725
transform 1 0 482908 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5249
timestamp 1676037725
transform 1 0 484012 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5261
timestamp 1676037725
transform 1 0 485116 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5273
timestamp 1676037725
transform 1 0 486220 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5285
timestamp 1676037725
transform 1 0 487324 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5291
timestamp 1676037725
transform 1 0 487876 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5293
timestamp 1676037725
transform 1 0 488060 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5305
timestamp 1676037725
transform 1 0 489164 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5317
timestamp 1676037725
transform 1 0 490268 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5329
timestamp 1676037725
transform 1 0 491372 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5341
timestamp 1676037725
transform 1 0 492476 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5347
timestamp 1676037725
transform 1 0 493028 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5349
timestamp 1676037725
transform 1 0 493212 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5361
timestamp 1676037725
transform 1 0 494316 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5373
timestamp 1676037725
transform 1 0 495420 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5385
timestamp 1676037725
transform 1 0 496524 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5397
timestamp 1676037725
transform 1 0 497628 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5403
timestamp 1676037725
transform 1 0 498180 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5405
timestamp 1676037725
transform 1 0 498364 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5417
timestamp 1676037725
transform 1 0 499468 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5429
timestamp 1676037725
transform 1 0 500572 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5441
timestamp 1676037725
transform 1 0 501676 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5453
timestamp 1676037725
transform 1 0 502780 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5459
timestamp 1676037725
transform 1 0 503332 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5461
timestamp 1676037725
transform 1 0 503516 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5473
timestamp 1676037725
transform 1 0 504620 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5485
timestamp 1676037725
transform 1 0 505724 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5497
timestamp 1676037725
transform 1 0 506828 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5509
timestamp 1676037725
transform 1 0 507932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5515
timestamp 1676037725
transform 1 0 508484 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5517
timestamp 1676037725
transform 1 0 508668 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5529
timestamp 1676037725
transform 1 0 509772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5541
timestamp 1676037725
transform 1 0 510876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5553
timestamp 1676037725
transform 1 0 511980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5565
timestamp 1676037725
transform 1 0 513084 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5571
timestamp 1676037725
transform 1 0 513636 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5573
timestamp 1676037725
transform 1 0 513820 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5585
timestamp 1676037725
transform 1 0 514924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5597
timestamp 1676037725
transform 1 0 516028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5609
timestamp 1676037725
transform 1 0 517132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5621
timestamp 1676037725
transform 1 0 518236 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5627
timestamp 1676037725
transform 1 0 518788 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5629
timestamp 1676037725
transform 1 0 518972 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5641
timestamp 1676037725
transform 1 0 520076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5653
timestamp 1676037725
transform 1 0 521180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5665
timestamp 1676037725
transform 1 0 522284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5677
timestamp 1676037725
transform 1 0 523388 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5683
timestamp 1676037725
transform 1 0 523940 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5685
timestamp 1676037725
transform 1 0 524124 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5697
timestamp 1676037725
transform 1 0 525228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5709
timestamp 1676037725
transform 1 0 526332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5721
timestamp 1676037725
transform 1 0 527436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1676037725
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1676037725
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1676037725
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1676037725
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1676037725
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1676037725
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1676037725
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1676037725
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1676037725
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1676037725
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1676037725
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1676037725
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1676037725
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1676037725
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1676037725
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1676037725
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1676037725
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1676037725
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1676037725
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1676037725
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1676037725
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1676037725
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1676037725
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1676037725
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1676037725
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1676037725
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1676037725
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1676037725
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1676037725
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1676037725
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1676037725
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1676037725
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 1676037725
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 1676037725
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1676037725
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1676037725
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1676037725
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_821
timestamp 1676037725
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 1676037725
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 1676037725
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_841
timestamp 1676037725
transform 1 0 78476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_853
timestamp 1676037725
transform 1 0 79580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_865
timestamp 1676037725
transform 1 0 80684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_877
timestamp 1676037725
transform 1 0 81788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_889
timestamp 1676037725
transform 1 0 82892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_895
timestamp 1676037725
transform 1 0 83444 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_897
timestamp 1676037725
transform 1 0 83628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_909
timestamp 1676037725
transform 1 0 84732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_921
timestamp 1676037725
transform 1 0 85836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_933
timestamp 1676037725
transform 1 0 86940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_945
timestamp 1676037725
transform 1 0 88044 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_951
timestamp 1676037725
transform 1 0 88596 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_953
timestamp 1676037725
transform 1 0 88780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_965
timestamp 1676037725
transform 1 0 89884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_977
timestamp 1676037725
transform 1 0 90988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_989
timestamp 1676037725
transform 1 0 92092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1001
timestamp 1676037725
transform 1 0 93196 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1007
timestamp 1676037725
transform 1 0 93748 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1009
timestamp 1676037725
transform 1 0 93932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1021
timestamp 1676037725
transform 1 0 95036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1033
timestamp 1676037725
transform 1 0 96140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1045
timestamp 1676037725
transform 1 0 97244 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1057
timestamp 1676037725
transform 1 0 98348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1063
timestamp 1676037725
transform 1 0 98900 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1065
timestamp 1676037725
transform 1 0 99084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1077
timestamp 1676037725
transform 1 0 100188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1089
timestamp 1676037725
transform 1 0 101292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1101
timestamp 1676037725
transform 1 0 102396 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1113
timestamp 1676037725
transform 1 0 103500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1119
timestamp 1676037725
transform 1 0 104052 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1121
timestamp 1676037725
transform 1 0 104236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1133
timestamp 1676037725
transform 1 0 105340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1145
timestamp 1676037725
transform 1 0 106444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1157
timestamp 1676037725
transform 1 0 107548 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1169
timestamp 1676037725
transform 1 0 108652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1175
timestamp 1676037725
transform 1 0 109204 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1177
timestamp 1676037725
transform 1 0 109388 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1189
timestamp 1676037725
transform 1 0 110492 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1201
timestamp 1676037725
transform 1 0 111596 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1213
timestamp 1676037725
transform 1 0 112700 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1225
timestamp 1676037725
transform 1 0 113804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1231
timestamp 1676037725
transform 1 0 114356 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1233
timestamp 1676037725
transform 1 0 114540 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1248
timestamp 1676037725
transform 1 0 115920 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1256
timestamp 1676037725
transform 1 0 116656 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1266
timestamp 1676037725
transform 1 0 117576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1270
timestamp 1676037725
transform 1 0 117944 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1280
timestamp 1676037725
transform 1 0 118864 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1286
timestamp 1676037725
transform 1 0 119416 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1289
timestamp 1676037725
transform 1 0 119692 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1293
timestamp 1676037725
transform 1 0 120060 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1296
timestamp 1676037725
transform 1 0 120336 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1302
timestamp 1676037725
transform 1 0 120888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1315
timestamp 1676037725
transform 1 0 122084 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1321
timestamp 1676037725
transform 1 0 122636 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1331
timestamp 1676037725
transform 1 0 123556 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1339
timestamp 1676037725
transform 1 0 124292 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1342
timestamp 1676037725
transform 1 0 124568 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1345
timestamp 1676037725
transform 1 0 124844 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1349
timestamp 1676037725
transform 1 0 125212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1361
timestamp 1676037725
transform 1 0 126316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1373
timestamp 1676037725
transform 1 0 127420 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1385
timestamp 1676037725
transform 1 0 128524 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1397
timestamp 1676037725
transform 1 0 129628 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1401
timestamp 1676037725
transform 1 0 129996 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1413
timestamp 1676037725
transform 1 0 131100 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1425
timestamp 1676037725
transform 1 0 132204 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1437
timestamp 1676037725
transform 1 0 133308 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1449
timestamp 1676037725
transform 1 0 134412 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1455
timestamp 1676037725
transform 1 0 134964 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1457
timestamp 1676037725
transform 1 0 135148 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1469
timestamp 1676037725
transform 1 0 136252 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1481
timestamp 1676037725
transform 1 0 137356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1493
timestamp 1676037725
transform 1 0 138460 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1505
timestamp 1676037725
transform 1 0 139564 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1511
timestamp 1676037725
transform 1 0 140116 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1513
timestamp 1676037725
transform 1 0 140300 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1525
timestamp 1676037725
transform 1 0 141404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1537
timestamp 1676037725
transform 1 0 142508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1549
timestamp 1676037725
transform 1 0 143612 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1561
timestamp 1676037725
transform 1 0 144716 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1567
timestamp 1676037725
transform 1 0 145268 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1569
timestamp 1676037725
transform 1 0 145452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1581
timestamp 1676037725
transform 1 0 146556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1593
timestamp 1676037725
transform 1 0 147660 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1605
timestamp 1676037725
transform 1 0 148764 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1617
timestamp 1676037725
transform 1 0 149868 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1623
timestamp 1676037725
transform 1 0 150420 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1625
timestamp 1676037725
transform 1 0 150604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1637
timestamp 1676037725
transform 1 0 151708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1649
timestamp 1676037725
transform 1 0 152812 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1661
timestamp 1676037725
transform 1 0 153916 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1673
timestamp 1676037725
transform 1 0 155020 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1679
timestamp 1676037725
transform 1 0 155572 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1681
timestamp 1676037725
transform 1 0 155756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1693
timestamp 1676037725
transform 1 0 156860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1705
timestamp 1676037725
transform 1 0 157964 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1717
timestamp 1676037725
transform 1 0 159068 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1729
timestamp 1676037725
transform 1 0 160172 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1735
timestamp 1676037725
transform 1 0 160724 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1737
timestamp 1676037725
transform 1 0 160908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1749
timestamp 1676037725
transform 1 0 162012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1761
timestamp 1676037725
transform 1 0 163116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1773
timestamp 1676037725
transform 1 0 164220 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1785
timestamp 1676037725
transform 1 0 165324 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1791
timestamp 1676037725
transform 1 0 165876 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1793
timestamp 1676037725
transform 1 0 166060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1805
timestamp 1676037725
transform 1 0 167164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1817
timestamp 1676037725
transform 1 0 168268 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1829
timestamp 1676037725
transform 1 0 169372 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1841
timestamp 1676037725
transform 1 0 170476 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1847
timestamp 1676037725
transform 1 0 171028 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1849
timestamp 1676037725
transform 1 0 171212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1861
timestamp 1676037725
transform 1 0 172316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1873
timestamp 1676037725
transform 1 0 173420 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1885
timestamp 1676037725
transform 1 0 174524 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1897
timestamp 1676037725
transform 1 0 175628 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1903
timestamp 1676037725
transform 1 0 176180 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1905
timestamp 1676037725
transform 1 0 176364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1917
timestamp 1676037725
transform 1 0 177468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1929
timestamp 1676037725
transform 1 0 178572 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1941
timestamp 1676037725
transform 1 0 179676 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1953
timestamp 1676037725
transform 1 0 180780 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1959
timestamp 1676037725
transform 1 0 181332 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1961
timestamp 1676037725
transform 1 0 181516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1973
timestamp 1676037725
transform 1 0 182620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1985
timestamp 1676037725
transform 1 0 183724 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1997
timestamp 1676037725
transform 1 0 184828 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2009
timestamp 1676037725
transform 1 0 185932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2015
timestamp 1676037725
transform 1 0 186484 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2017
timestamp 1676037725
transform 1 0 186668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2029
timestamp 1676037725
transform 1 0 187772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2041
timestamp 1676037725
transform 1 0 188876 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2053
timestamp 1676037725
transform 1 0 189980 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2065
timestamp 1676037725
transform 1 0 191084 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2071
timestamp 1676037725
transform 1 0 191636 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2073
timestamp 1676037725
transform 1 0 191820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2085
timestamp 1676037725
transform 1 0 192924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2097
timestamp 1676037725
transform 1 0 194028 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2109
timestamp 1676037725
transform 1 0 195132 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2121
timestamp 1676037725
transform 1 0 196236 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2127
timestamp 1676037725
transform 1 0 196788 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2129
timestamp 1676037725
transform 1 0 196972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2141
timestamp 1676037725
transform 1 0 198076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2153
timestamp 1676037725
transform 1 0 199180 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2165
timestamp 1676037725
transform 1 0 200284 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2177
timestamp 1676037725
transform 1 0 201388 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2183
timestamp 1676037725
transform 1 0 201940 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2185
timestamp 1676037725
transform 1 0 202124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2197
timestamp 1676037725
transform 1 0 203228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2209
timestamp 1676037725
transform 1 0 204332 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2221
timestamp 1676037725
transform 1 0 205436 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2233
timestamp 1676037725
transform 1 0 206540 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2239
timestamp 1676037725
transform 1 0 207092 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2241
timestamp 1676037725
transform 1 0 207276 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_2255
timestamp 1676037725
transform 1 0 208564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_2261
timestamp 1676037725
transform 1 0 209116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_2274
timestamp 1676037725
transform 1 0 210312 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2282
timestamp 1676037725
transform 1 0 211048 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_2292
timestamp 1676037725
transform 1 0 211968 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_2297
timestamp 1676037725
transform 1 0 212428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_2302
timestamp 1676037725
transform 1 0 212888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_2315
timestamp 1676037725
transform 1 0 214084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_2332
timestamp 1676037725
transform 1 0 215648 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_2349
timestamp 1676037725
transform 1 0 217212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_2353
timestamp 1676037725
transform 1 0 217580 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_2357
timestamp 1676037725
transform 1 0 217948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2361
timestamp 1676037725
transform 1 0 218316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_2364
timestamp 1676037725
transform 1 0 218592 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2372
timestamp 1676037725
transform 1 0 219328 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2375
timestamp 1676037725
transform 1 0 219604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2387
timestamp 1676037725
transform 1 0 220708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_2399
timestamp 1676037725
transform 1 0 221812 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2407
timestamp 1676037725
transform 1 0 222548 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2409
timestamp 1676037725
transform 1 0 222732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2421
timestamp 1676037725
transform 1 0 223836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2433
timestamp 1676037725
transform 1 0 224940 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2445
timestamp 1676037725
transform 1 0 226044 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2457
timestamp 1676037725
transform 1 0 227148 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2463
timestamp 1676037725
transform 1 0 227700 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2465
timestamp 1676037725
transform 1 0 227884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2477
timestamp 1676037725
transform 1 0 228988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2489
timestamp 1676037725
transform 1 0 230092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2501
timestamp 1676037725
transform 1 0 231196 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2513
timestamp 1676037725
transform 1 0 232300 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2519
timestamp 1676037725
transform 1 0 232852 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2521
timestamp 1676037725
transform 1 0 233036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2533
timestamp 1676037725
transform 1 0 234140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2545
timestamp 1676037725
transform 1 0 235244 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2557
timestamp 1676037725
transform 1 0 236348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2569
timestamp 1676037725
transform 1 0 237452 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2575
timestamp 1676037725
transform 1 0 238004 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2577
timestamp 1676037725
transform 1 0 238188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2589
timestamp 1676037725
transform 1 0 239292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2601
timestamp 1676037725
transform 1 0 240396 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2613
timestamp 1676037725
transform 1 0 241500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2625
timestamp 1676037725
transform 1 0 242604 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2631
timestamp 1676037725
transform 1 0 243156 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2633
timestamp 1676037725
transform 1 0 243340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2645
timestamp 1676037725
transform 1 0 244444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2657
timestamp 1676037725
transform 1 0 245548 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2669
timestamp 1676037725
transform 1 0 246652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2681
timestamp 1676037725
transform 1 0 247756 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2687
timestamp 1676037725
transform 1 0 248308 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2689
timestamp 1676037725
transform 1 0 248492 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2701
timestamp 1676037725
transform 1 0 249596 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2713
timestamp 1676037725
transform 1 0 250700 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2725
timestamp 1676037725
transform 1 0 251804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2737
timestamp 1676037725
transform 1 0 252908 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2743
timestamp 1676037725
transform 1 0 253460 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2745
timestamp 1676037725
transform 1 0 253644 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2757
timestamp 1676037725
transform 1 0 254748 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2769
timestamp 1676037725
transform 1 0 255852 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2781
timestamp 1676037725
transform 1 0 256956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2793
timestamp 1676037725
transform 1 0 258060 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2799
timestamp 1676037725
transform 1 0 258612 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2801
timestamp 1676037725
transform 1 0 258796 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2813
timestamp 1676037725
transform 1 0 259900 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2825
timestamp 1676037725
transform 1 0 261004 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2837
timestamp 1676037725
transform 1 0 262108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2849
timestamp 1676037725
transform 1 0 263212 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2855
timestamp 1676037725
transform 1 0 263764 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2857
timestamp 1676037725
transform 1 0 263948 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2869
timestamp 1676037725
transform 1 0 265052 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2881
timestamp 1676037725
transform 1 0 266156 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2893
timestamp 1676037725
transform 1 0 267260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2905
timestamp 1676037725
transform 1 0 268364 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2911
timestamp 1676037725
transform 1 0 268916 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2913
timestamp 1676037725
transform 1 0 269100 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2925
timestamp 1676037725
transform 1 0 270204 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2937
timestamp 1676037725
transform 1 0 271308 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2949
timestamp 1676037725
transform 1 0 272412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2961
timestamp 1676037725
transform 1 0 273516 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2967
timestamp 1676037725
transform 1 0 274068 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2969
timestamp 1676037725
transform 1 0 274252 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2981
timestamp 1676037725
transform 1 0 275356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2993
timestamp 1676037725
transform 1 0 276460 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3005
timestamp 1676037725
transform 1 0 277564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3017
timestamp 1676037725
transform 1 0 278668 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3023
timestamp 1676037725
transform 1 0 279220 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3025
timestamp 1676037725
transform 1 0 279404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3037
timestamp 1676037725
transform 1 0 280508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3049
timestamp 1676037725
transform 1 0 281612 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3061
timestamp 1676037725
transform 1 0 282716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3073
timestamp 1676037725
transform 1 0 283820 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3079
timestamp 1676037725
transform 1 0 284372 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3081
timestamp 1676037725
transform 1 0 284556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3093
timestamp 1676037725
transform 1 0 285660 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3105
timestamp 1676037725
transform 1 0 286764 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3117
timestamp 1676037725
transform 1 0 287868 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3129
timestamp 1676037725
transform 1 0 288972 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3135
timestamp 1676037725
transform 1 0 289524 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3137
timestamp 1676037725
transform 1 0 289708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3149
timestamp 1676037725
transform 1 0 290812 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3161
timestamp 1676037725
transform 1 0 291916 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3173
timestamp 1676037725
transform 1 0 293020 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3185
timestamp 1676037725
transform 1 0 294124 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3191
timestamp 1676037725
transform 1 0 294676 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3193
timestamp 1676037725
transform 1 0 294860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3205
timestamp 1676037725
transform 1 0 295964 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3217
timestamp 1676037725
transform 1 0 297068 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3229
timestamp 1676037725
transform 1 0 298172 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3241
timestamp 1676037725
transform 1 0 299276 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3247
timestamp 1676037725
transform 1 0 299828 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3249
timestamp 1676037725
transform 1 0 300012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3261
timestamp 1676037725
transform 1 0 301116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3273
timestamp 1676037725
transform 1 0 302220 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3285
timestamp 1676037725
transform 1 0 303324 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3293
timestamp 1676037725
transform 1 0 304060 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3296
timestamp 1676037725
transform 1 0 304336 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3302
timestamp 1676037725
transform 1 0 304888 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3305
timestamp 1676037725
transform 1 0 305164 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3309
timestamp 1676037725
transform 1 0 305532 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3313
timestamp 1676037725
transform 1 0 305900 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3320
timestamp 1676037725
transform 1 0 306544 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3326
timestamp 1676037725
transform 1 0 307096 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3334
timestamp 1676037725
transform 1 0 307832 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3342
timestamp 1676037725
transform 1 0 308568 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3349
timestamp 1676037725
transform 1 0 309212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3355
timestamp 1676037725
transform 1 0 309764 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3359
timestamp 1676037725
transform 1 0 310132 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3361
timestamp 1676037725
transform 1 0 310316 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3367
timestamp 1676037725
transform 1 0 310868 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3373
timestamp 1676037725
transform 1 0 311420 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3385
timestamp 1676037725
transform 1 0 312524 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3397
timestamp 1676037725
transform 1 0 313628 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3409
timestamp 1676037725
transform 1 0 314732 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3415
timestamp 1676037725
transform 1 0 315284 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3417
timestamp 1676037725
transform 1 0 315468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3429
timestamp 1676037725
transform 1 0 316572 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3441
timestamp 1676037725
transform 1 0 317676 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3453
timestamp 1676037725
transform 1 0 318780 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3465
timestamp 1676037725
transform 1 0 319884 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3471
timestamp 1676037725
transform 1 0 320436 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3473
timestamp 1676037725
transform 1 0 320620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3485
timestamp 1676037725
transform 1 0 321724 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3497
timestamp 1676037725
transform 1 0 322828 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3509
timestamp 1676037725
transform 1 0 323932 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3521
timestamp 1676037725
transform 1 0 325036 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3527
timestamp 1676037725
transform 1 0 325588 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3529
timestamp 1676037725
transform 1 0 325772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3541
timestamp 1676037725
transform 1 0 326876 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3553
timestamp 1676037725
transform 1 0 327980 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3565
timestamp 1676037725
transform 1 0 329084 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3577
timestamp 1676037725
transform 1 0 330188 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3583
timestamp 1676037725
transform 1 0 330740 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3585
timestamp 1676037725
transform 1 0 330924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3597
timestamp 1676037725
transform 1 0 332028 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3609
timestamp 1676037725
transform 1 0 333132 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3621
timestamp 1676037725
transform 1 0 334236 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3633
timestamp 1676037725
transform 1 0 335340 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3639
timestamp 1676037725
transform 1 0 335892 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3641
timestamp 1676037725
transform 1 0 336076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3653
timestamp 1676037725
transform 1 0 337180 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3665
timestamp 1676037725
transform 1 0 338284 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3677
timestamp 1676037725
transform 1 0 339388 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3689
timestamp 1676037725
transform 1 0 340492 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3695
timestamp 1676037725
transform 1 0 341044 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3697
timestamp 1676037725
transform 1 0 341228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3709
timestamp 1676037725
transform 1 0 342332 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3721
timestamp 1676037725
transform 1 0 343436 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3733
timestamp 1676037725
transform 1 0 344540 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3745
timestamp 1676037725
transform 1 0 345644 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3751
timestamp 1676037725
transform 1 0 346196 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3753
timestamp 1676037725
transform 1 0 346380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3765
timestamp 1676037725
transform 1 0 347484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3777
timestamp 1676037725
transform 1 0 348588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3789
timestamp 1676037725
transform 1 0 349692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3801
timestamp 1676037725
transform 1 0 350796 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3807
timestamp 1676037725
transform 1 0 351348 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3809
timestamp 1676037725
transform 1 0 351532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3821
timestamp 1676037725
transform 1 0 352636 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3833
timestamp 1676037725
transform 1 0 353740 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3845
timestamp 1676037725
transform 1 0 354844 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3857
timestamp 1676037725
transform 1 0 355948 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3863
timestamp 1676037725
transform 1 0 356500 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3865
timestamp 1676037725
transform 1 0 356684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3877
timestamp 1676037725
transform 1 0 357788 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3889
timestamp 1676037725
transform 1 0 358892 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3901
timestamp 1676037725
transform 1 0 359996 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3913
timestamp 1676037725
transform 1 0 361100 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3919
timestamp 1676037725
transform 1 0 361652 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3921
timestamp 1676037725
transform 1 0 361836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3933
timestamp 1676037725
transform 1 0 362940 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3945
timestamp 1676037725
transform 1 0 364044 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3957
timestamp 1676037725
transform 1 0 365148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3969
timestamp 1676037725
transform 1 0 366252 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3975
timestamp 1676037725
transform 1 0 366804 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3977
timestamp 1676037725
transform 1 0 366988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3989
timestamp 1676037725
transform 1 0 368092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4001
timestamp 1676037725
transform 1 0 369196 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4013
timestamp 1676037725
transform 1 0 370300 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4025
timestamp 1676037725
transform 1 0 371404 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4031
timestamp 1676037725
transform 1 0 371956 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4033
timestamp 1676037725
transform 1 0 372140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4045
timestamp 1676037725
transform 1 0 373244 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4057
timestamp 1676037725
transform 1 0 374348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4069
timestamp 1676037725
transform 1 0 375452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4081
timestamp 1676037725
transform 1 0 376556 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4087
timestamp 1676037725
transform 1 0 377108 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4089
timestamp 1676037725
transform 1 0 377292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4101
timestamp 1676037725
transform 1 0 378396 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4113
timestamp 1676037725
transform 1 0 379500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4125
timestamp 1676037725
transform 1 0 380604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4137
timestamp 1676037725
transform 1 0 381708 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4143
timestamp 1676037725
transform 1 0 382260 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4145
timestamp 1676037725
transform 1 0 382444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4157
timestamp 1676037725
transform 1 0 383548 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4169
timestamp 1676037725
transform 1 0 384652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4181
timestamp 1676037725
transform 1 0 385756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4193
timestamp 1676037725
transform 1 0 386860 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4199
timestamp 1676037725
transform 1 0 387412 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4201
timestamp 1676037725
transform 1 0 387596 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4213
timestamp 1676037725
transform 1 0 388700 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4225
timestamp 1676037725
transform 1 0 389804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4237
timestamp 1676037725
transform 1 0 390908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4249
timestamp 1676037725
transform 1 0 392012 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4255
timestamp 1676037725
transform 1 0 392564 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4257
timestamp 1676037725
transform 1 0 392748 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4269
timestamp 1676037725
transform 1 0 393852 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4281
timestamp 1676037725
transform 1 0 394956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4293
timestamp 1676037725
transform 1 0 396060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4305
timestamp 1676037725
transform 1 0 397164 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4311
timestamp 1676037725
transform 1 0 397716 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4313
timestamp 1676037725
transform 1 0 397900 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4325
timestamp 1676037725
transform 1 0 399004 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4337
timestamp 1676037725
transform 1 0 400108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4349
timestamp 1676037725
transform 1 0 401212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4361
timestamp 1676037725
transform 1 0 402316 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4367
timestamp 1676037725
transform 1 0 402868 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4369
timestamp 1676037725
transform 1 0 403052 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4381
timestamp 1676037725
transform 1 0 404156 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4393
timestamp 1676037725
transform 1 0 405260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4405
timestamp 1676037725
transform 1 0 406364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4417
timestamp 1676037725
transform 1 0 407468 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4423
timestamp 1676037725
transform 1 0 408020 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4425
timestamp 1676037725
transform 1 0 408204 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4437
timestamp 1676037725
transform 1 0 409308 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4449
timestamp 1676037725
transform 1 0 410412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4461
timestamp 1676037725
transform 1 0 411516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4473
timestamp 1676037725
transform 1 0 412620 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4479
timestamp 1676037725
transform 1 0 413172 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4481
timestamp 1676037725
transform 1 0 413356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4493
timestamp 1676037725
transform 1 0 414460 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4505
timestamp 1676037725
transform 1 0 415564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4517
timestamp 1676037725
transform 1 0 416668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4529
timestamp 1676037725
transform 1 0 417772 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4535
timestamp 1676037725
transform 1 0 418324 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4537
timestamp 1676037725
transform 1 0 418508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4549
timestamp 1676037725
transform 1 0 419612 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4561
timestamp 1676037725
transform 1 0 420716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4573
timestamp 1676037725
transform 1 0 421820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4585
timestamp 1676037725
transform 1 0 422924 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4591
timestamp 1676037725
transform 1 0 423476 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4593
timestamp 1676037725
transform 1 0 423660 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4605
timestamp 1676037725
transform 1 0 424764 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4617
timestamp 1676037725
transform 1 0 425868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4629
timestamp 1676037725
transform 1 0 426972 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4641
timestamp 1676037725
transform 1 0 428076 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4647
timestamp 1676037725
transform 1 0 428628 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4649
timestamp 1676037725
transform 1 0 428812 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4661
timestamp 1676037725
transform 1 0 429916 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4673
timestamp 1676037725
transform 1 0 431020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4685
timestamp 1676037725
transform 1 0 432124 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4697
timestamp 1676037725
transform 1 0 433228 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4703
timestamp 1676037725
transform 1 0 433780 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4705
timestamp 1676037725
transform 1 0 433964 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4717
timestamp 1676037725
transform 1 0 435068 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4729
timestamp 1676037725
transform 1 0 436172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4741
timestamp 1676037725
transform 1 0 437276 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4753
timestamp 1676037725
transform 1 0 438380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4759
timestamp 1676037725
transform 1 0 438932 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4761
timestamp 1676037725
transform 1 0 439116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4773
timestamp 1676037725
transform 1 0 440220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4785
timestamp 1676037725
transform 1 0 441324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4797
timestamp 1676037725
transform 1 0 442428 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4809
timestamp 1676037725
transform 1 0 443532 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4815
timestamp 1676037725
transform 1 0 444084 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4817
timestamp 1676037725
transform 1 0 444268 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4829
timestamp 1676037725
transform 1 0 445372 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4841
timestamp 1676037725
transform 1 0 446476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4853
timestamp 1676037725
transform 1 0 447580 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4865
timestamp 1676037725
transform 1 0 448684 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4871
timestamp 1676037725
transform 1 0 449236 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4873
timestamp 1676037725
transform 1 0 449420 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4885
timestamp 1676037725
transform 1 0 450524 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4897
timestamp 1676037725
transform 1 0 451628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4909
timestamp 1676037725
transform 1 0 452732 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4921
timestamp 1676037725
transform 1 0 453836 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4927
timestamp 1676037725
transform 1 0 454388 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4929
timestamp 1676037725
transform 1 0 454572 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4941
timestamp 1676037725
transform 1 0 455676 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4953
timestamp 1676037725
transform 1 0 456780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4965
timestamp 1676037725
transform 1 0 457884 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4977
timestamp 1676037725
transform 1 0 458988 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4983
timestamp 1676037725
transform 1 0 459540 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4985
timestamp 1676037725
transform 1 0 459724 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4997
timestamp 1676037725
transform 1 0 460828 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5009
timestamp 1676037725
transform 1 0 461932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5021
timestamp 1676037725
transform 1 0 463036 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5033
timestamp 1676037725
transform 1 0 464140 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5039
timestamp 1676037725
transform 1 0 464692 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5041
timestamp 1676037725
transform 1 0 464876 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5053
timestamp 1676037725
transform 1 0 465980 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5065
timestamp 1676037725
transform 1 0 467084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5077
timestamp 1676037725
transform 1 0 468188 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5089
timestamp 1676037725
transform 1 0 469292 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5095
timestamp 1676037725
transform 1 0 469844 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5097
timestamp 1676037725
transform 1 0 470028 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5109
timestamp 1676037725
transform 1 0 471132 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5121
timestamp 1676037725
transform 1 0 472236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5133
timestamp 1676037725
transform 1 0 473340 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5145
timestamp 1676037725
transform 1 0 474444 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5151
timestamp 1676037725
transform 1 0 474996 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5153
timestamp 1676037725
transform 1 0 475180 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5165
timestamp 1676037725
transform 1 0 476284 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5177
timestamp 1676037725
transform 1 0 477388 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5189
timestamp 1676037725
transform 1 0 478492 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5201
timestamp 1676037725
transform 1 0 479596 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5207
timestamp 1676037725
transform 1 0 480148 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5209
timestamp 1676037725
transform 1 0 480332 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5221
timestamp 1676037725
transform 1 0 481436 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5233
timestamp 1676037725
transform 1 0 482540 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5245
timestamp 1676037725
transform 1 0 483644 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5257
timestamp 1676037725
transform 1 0 484748 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5263
timestamp 1676037725
transform 1 0 485300 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5265
timestamp 1676037725
transform 1 0 485484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5277
timestamp 1676037725
transform 1 0 486588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5289
timestamp 1676037725
transform 1 0 487692 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5301
timestamp 1676037725
transform 1 0 488796 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5313
timestamp 1676037725
transform 1 0 489900 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5319
timestamp 1676037725
transform 1 0 490452 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5321
timestamp 1676037725
transform 1 0 490636 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5333
timestamp 1676037725
transform 1 0 491740 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5345
timestamp 1676037725
transform 1 0 492844 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5357
timestamp 1676037725
transform 1 0 493948 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5369
timestamp 1676037725
transform 1 0 495052 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5375
timestamp 1676037725
transform 1 0 495604 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5377
timestamp 1676037725
transform 1 0 495788 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5389
timestamp 1676037725
transform 1 0 496892 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5401
timestamp 1676037725
transform 1 0 497996 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5413
timestamp 1676037725
transform 1 0 499100 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5425
timestamp 1676037725
transform 1 0 500204 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5431
timestamp 1676037725
transform 1 0 500756 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5433
timestamp 1676037725
transform 1 0 500940 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5445
timestamp 1676037725
transform 1 0 502044 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5457
timestamp 1676037725
transform 1 0 503148 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5469
timestamp 1676037725
transform 1 0 504252 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5481
timestamp 1676037725
transform 1 0 505356 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5487
timestamp 1676037725
transform 1 0 505908 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5489
timestamp 1676037725
transform 1 0 506092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5501
timestamp 1676037725
transform 1 0 507196 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5513
timestamp 1676037725
transform 1 0 508300 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5525
timestamp 1676037725
transform 1 0 509404 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5537
timestamp 1676037725
transform 1 0 510508 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5543
timestamp 1676037725
transform 1 0 511060 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5545
timestamp 1676037725
transform 1 0 511244 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5557
timestamp 1676037725
transform 1 0 512348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5569
timestamp 1676037725
transform 1 0 513452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5581
timestamp 1676037725
transform 1 0 514556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5593
timestamp 1676037725
transform 1 0 515660 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5599
timestamp 1676037725
transform 1 0 516212 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5601
timestamp 1676037725
transform 1 0 516396 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5613
timestamp 1676037725
transform 1 0 517500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5625
timestamp 1676037725
transform 1 0 518604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5637
timestamp 1676037725
transform 1 0 519708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5649
timestamp 1676037725
transform 1 0 520812 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5655
timestamp 1676037725
transform 1 0 521364 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5657
timestamp 1676037725
transform 1 0 521548 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5669
timestamp 1676037725
transform 1 0 522652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5681
timestamp 1676037725
transform 1 0 523756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5693
timestamp 1676037725
transform 1 0 524860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5705
timestamp 1676037725
transform 1 0 525964 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5711
timestamp 1676037725
transform 1 0 526516 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5713
timestamp 1676037725
transform 1 0 526700 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_5725
timestamp 1676037725
transform 1 0 527804 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1676037725
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1676037725
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1676037725
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1676037725
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1676037725
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1676037725
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1676037725
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1676037725
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1676037725
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1676037725
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1676037725
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1676037725
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1676037725
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1676037725
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1676037725
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1676037725
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1676037725
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1676037725
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1676037725
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1676037725
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1676037725
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1676037725
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1676037725
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1676037725
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1676037725
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1676037725
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1676037725
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1676037725
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1676037725
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1676037725
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1676037725
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1676037725
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1676037725
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1676037725
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1676037725
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1676037725
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1676037725
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1676037725
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_781
timestamp 1676037725
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_793
timestamp 1676037725
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 1676037725
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 1676037725
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1676037725
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_825
timestamp 1676037725
transform 1 0 77004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_837
timestamp 1676037725
transform 1 0 78108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_849
timestamp 1676037725
transform 1 0 79212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_861
timestamp 1676037725
transform 1 0 80316 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_867
timestamp 1676037725
transform 1 0 80868 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_869
timestamp 1676037725
transform 1 0 81052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_881
timestamp 1676037725
transform 1 0 82156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_893
timestamp 1676037725
transform 1 0 83260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_905
timestamp 1676037725
transform 1 0 84364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_917
timestamp 1676037725
transform 1 0 85468 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_923
timestamp 1676037725
transform 1 0 86020 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_925
timestamp 1676037725
transform 1 0 86204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_937
timestamp 1676037725
transform 1 0 87308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_949
timestamp 1676037725
transform 1 0 88412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_961
timestamp 1676037725
transform 1 0 89516 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_973
timestamp 1676037725
transform 1 0 90620 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_979
timestamp 1676037725
transform 1 0 91172 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_981
timestamp 1676037725
transform 1 0 91356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_993
timestamp 1676037725
transform 1 0 92460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1005
timestamp 1676037725
transform 1 0 93564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1017
timestamp 1676037725
transform 1 0 94668 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1029
timestamp 1676037725
transform 1 0 95772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1035
timestamp 1676037725
transform 1 0 96324 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1037
timestamp 1676037725
transform 1 0 96508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1049
timestamp 1676037725
transform 1 0 97612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1061
timestamp 1676037725
transform 1 0 98716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1073
timestamp 1676037725
transform 1 0 99820 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1085
timestamp 1676037725
transform 1 0 100924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1091
timestamp 1676037725
transform 1 0 101476 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1093
timestamp 1676037725
transform 1 0 101660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1105
timestamp 1676037725
transform 1 0 102764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1117
timestamp 1676037725
transform 1 0 103868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1129
timestamp 1676037725
transform 1 0 104972 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1141
timestamp 1676037725
transform 1 0 106076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1147
timestamp 1676037725
transform 1 0 106628 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1149
timestamp 1676037725
transform 1 0 106812 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1161
timestamp 1676037725
transform 1 0 107916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1173
timestamp 1676037725
transform 1 0 109020 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1185
timestamp 1676037725
transform 1 0 110124 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1197
timestamp 1676037725
transform 1 0 111228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1203
timestamp 1676037725
transform 1 0 111780 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1205
timestamp 1676037725
transform 1 0 111964 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1217
timestamp 1676037725
transform 1 0 113068 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1229
timestamp 1676037725
transform 1 0 114172 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1241
timestamp 1676037725
transform 1 0 115276 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1244
timestamp 1676037725
transform 1 0 115552 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1250
timestamp 1676037725
transform 1 0 116104 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1254
timestamp 1676037725
transform 1 0 116472 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_1257
timestamp 1676037725
transform 1 0 116748 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1261
timestamp 1676037725
transform 1 0 117116 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1267
timestamp 1676037725
transform 1 0 117668 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1270
timestamp 1676037725
transform 1 0 117944 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1276
timestamp 1676037725
transform 1 0 118496 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1282
timestamp 1676037725
transform 1 0 119048 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1288
timestamp 1676037725
transform 1 0 119600 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1302
timestamp 1676037725
transform 1 0 120888 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1308
timestamp 1676037725
transform 1 0 121440 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1317
timestamp 1676037725
transform 1 0 122268 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1321
timestamp 1676037725
transform 1 0 122636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1333
timestamp 1676037725
transform 1 0 123740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1345
timestamp 1676037725
transform 1 0 124844 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1357
timestamp 1676037725
transform 1 0 125948 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_1369
timestamp 1676037725
transform 1 0 127052 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1373
timestamp 1676037725
transform 1 0 127420 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1385
timestamp 1676037725
transform 1 0 128524 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1397
timestamp 1676037725
transform 1 0 129628 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1409
timestamp 1676037725
transform 1 0 130732 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1421
timestamp 1676037725
transform 1 0 131836 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1427
timestamp 1676037725
transform 1 0 132388 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1429
timestamp 1676037725
transform 1 0 132572 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1441
timestamp 1676037725
transform 1 0 133676 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1453
timestamp 1676037725
transform 1 0 134780 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1465
timestamp 1676037725
transform 1 0 135884 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1477
timestamp 1676037725
transform 1 0 136988 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1483
timestamp 1676037725
transform 1 0 137540 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1485
timestamp 1676037725
transform 1 0 137724 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1497
timestamp 1676037725
transform 1 0 138828 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1509
timestamp 1676037725
transform 1 0 139932 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1521
timestamp 1676037725
transform 1 0 141036 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1533
timestamp 1676037725
transform 1 0 142140 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1539
timestamp 1676037725
transform 1 0 142692 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1541
timestamp 1676037725
transform 1 0 142876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1553
timestamp 1676037725
transform 1 0 143980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1565
timestamp 1676037725
transform 1 0 145084 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1577
timestamp 1676037725
transform 1 0 146188 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1589
timestamp 1676037725
transform 1 0 147292 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1595
timestamp 1676037725
transform 1 0 147844 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1597
timestamp 1676037725
transform 1 0 148028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1609
timestamp 1676037725
transform 1 0 149132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1621
timestamp 1676037725
transform 1 0 150236 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1633
timestamp 1676037725
transform 1 0 151340 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1645
timestamp 1676037725
transform 1 0 152444 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1651
timestamp 1676037725
transform 1 0 152996 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1653
timestamp 1676037725
transform 1 0 153180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1665
timestamp 1676037725
transform 1 0 154284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1677
timestamp 1676037725
transform 1 0 155388 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1689
timestamp 1676037725
transform 1 0 156492 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1701
timestamp 1676037725
transform 1 0 157596 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1707
timestamp 1676037725
transform 1 0 158148 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1709
timestamp 1676037725
transform 1 0 158332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1721
timestamp 1676037725
transform 1 0 159436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1733
timestamp 1676037725
transform 1 0 160540 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1745
timestamp 1676037725
transform 1 0 161644 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1757
timestamp 1676037725
transform 1 0 162748 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1763
timestamp 1676037725
transform 1 0 163300 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1765
timestamp 1676037725
transform 1 0 163484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1777
timestamp 1676037725
transform 1 0 164588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1789
timestamp 1676037725
transform 1 0 165692 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1801
timestamp 1676037725
transform 1 0 166796 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1813
timestamp 1676037725
transform 1 0 167900 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1819
timestamp 1676037725
transform 1 0 168452 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1821
timestamp 1676037725
transform 1 0 168636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1833
timestamp 1676037725
transform 1 0 169740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1845
timestamp 1676037725
transform 1 0 170844 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1857
timestamp 1676037725
transform 1 0 171948 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1869
timestamp 1676037725
transform 1 0 173052 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1875
timestamp 1676037725
transform 1 0 173604 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1877
timestamp 1676037725
transform 1 0 173788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1889
timestamp 1676037725
transform 1 0 174892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1901
timestamp 1676037725
transform 1 0 175996 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1913
timestamp 1676037725
transform 1 0 177100 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1925
timestamp 1676037725
transform 1 0 178204 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1931
timestamp 1676037725
transform 1 0 178756 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1933
timestamp 1676037725
transform 1 0 178940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1945
timestamp 1676037725
transform 1 0 180044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1957
timestamp 1676037725
transform 1 0 181148 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1969
timestamp 1676037725
transform 1 0 182252 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1981
timestamp 1676037725
transform 1 0 183356 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1987
timestamp 1676037725
transform 1 0 183908 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1989
timestamp 1676037725
transform 1 0 184092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2001
timestamp 1676037725
transform 1 0 185196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2013
timestamp 1676037725
transform 1 0 186300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2025
timestamp 1676037725
transform 1 0 187404 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2037
timestamp 1676037725
transform 1 0 188508 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2043
timestamp 1676037725
transform 1 0 189060 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2045
timestamp 1676037725
transform 1 0 189244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2057
timestamp 1676037725
transform 1 0 190348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2069
timestamp 1676037725
transform 1 0 191452 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2081
timestamp 1676037725
transform 1 0 192556 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2093
timestamp 1676037725
transform 1 0 193660 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2099
timestamp 1676037725
transform 1 0 194212 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2101
timestamp 1676037725
transform 1 0 194396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2113
timestamp 1676037725
transform 1 0 195500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2125
timestamp 1676037725
transform 1 0 196604 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2137
timestamp 1676037725
transform 1 0 197708 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2149
timestamp 1676037725
transform 1 0 198812 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2155
timestamp 1676037725
transform 1 0 199364 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2157
timestamp 1676037725
transform 1 0 199548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2169
timestamp 1676037725
transform 1 0 200652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2181
timestamp 1676037725
transform 1 0 201756 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2193
timestamp 1676037725
transform 1 0 202860 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2205
timestamp 1676037725
transform 1 0 203964 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2211
timestamp 1676037725
transform 1 0 204516 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2213
timestamp 1676037725
transform 1 0 204700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2225
timestamp 1676037725
transform 1 0 205804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2237
timestamp 1676037725
transform 1 0 206908 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2249
timestamp 1676037725
transform 1 0 208012 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2261
timestamp 1676037725
transform 1 0 209116 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2267
timestamp 1676037725
transform 1 0 209668 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_2269
timestamp 1676037725
transform 1 0 209852 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2273
timestamp 1676037725
transform 1 0 210220 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_2276
timestamp 1676037725
transform 1 0 210496 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2280
timestamp 1676037725
transform 1 0 210864 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_2283
timestamp 1676037725
transform 1 0 211140 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2289
timestamp 1676037725
transform 1 0 211692 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2295
timestamp 1676037725
transform 1 0 212244 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_2298
timestamp 1676037725
transform 1 0 212520 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_2304
timestamp 1676037725
transform 1 0 213072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_2310
timestamp 1676037725
transform 1 0 213624 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_2316
timestamp 1676037725
transform 1 0 214176 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_2322
timestamp 1676037725
transform 1 0 214728 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2325
timestamp 1676037725
transform 1 0 215004 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2331
timestamp 1676037725
transform 1 0 215556 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_2334
timestamp 1676037725
transform 1 0 215832 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2342
timestamp 1676037725
transform 1 0 216568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_2345
timestamp 1676037725
transform 1 0 216844 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_2351
timestamp 1676037725
transform 1 0 217396 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2357
timestamp 1676037725
transform 1 0 217948 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_2369
timestamp 1676037725
transform 1 0 219052 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_2377
timestamp 1676037725
transform 1 0 219788 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2381
timestamp 1676037725
transform 1 0 220156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2393
timestamp 1676037725
transform 1 0 221260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2405
timestamp 1676037725
transform 1 0 222364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2417
timestamp 1676037725
transform 1 0 223468 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2429
timestamp 1676037725
transform 1 0 224572 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2435
timestamp 1676037725
transform 1 0 225124 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2437
timestamp 1676037725
transform 1 0 225308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2449
timestamp 1676037725
transform 1 0 226412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2461
timestamp 1676037725
transform 1 0 227516 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2473
timestamp 1676037725
transform 1 0 228620 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2485
timestamp 1676037725
transform 1 0 229724 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2491
timestamp 1676037725
transform 1 0 230276 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2493
timestamp 1676037725
transform 1 0 230460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2505
timestamp 1676037725
transform 1 0 231564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2517
timestamp 1676037725
transform 1 0 232668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2529
timestamp 1676037725
transform 1 0 233772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2541
timestamp 1676037725
transform 1 0 234876 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2547
timestamp 1676037725
transform 1 0 235428 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2549
timestamp 1676037725
transform 1 0 235612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2561
timestamp 1676037725
transform 1 0 236716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2573
timestamp 1676037725
transform 1 0 237820 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2585
timestamp 1676037725
transform 1 0 238924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2597
timestamp 1676037725
transform 1 0 240028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2603
timestamp 1676037725
transform 1 0 240580 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2605
timestamp 1676037725
transform 1 0 240764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2617
timestamp 1676037725
transform 1 0 241868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2629
timestamp 1676037725
transform 1 0 242972 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2641
timestamp 1676037725
transform 1 0 244076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2653
timestamp 1676037725
transform 1 0 245180 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2659
timestamp 1676037725
transform 1 0 245732 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2661
timestamp 1676037725
transform 1 0 245916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2673
timestamp 1676037725
transform 1 0 247020 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2685
timestamp 1676037725
transform 1 0 248124 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2697
timestamp 1676037725
transform 1 0 249228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2709
timestamp 1676037725
transform 1 0 250332 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2715
timestamp 1676037725
transform 1 0 250884 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2717
timestamp 1676037725
transform 1 0 251068 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2729
timestamp 1676037725
transform 1 0 252172 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2741
timestamp 1676037725
transform 1 0 253276 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2753
timestamp 1676037725
transform 1 0 254380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2765
timestamp 1676037725
transform 1 0 255484 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2771
timestamp 1676037725
transform 1 0 256036 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2773
timestamp 1676037725
transform 1 0 256220 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2785
timestamp 1676037725
transform 1 0 257324 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2797
timestamp 1676037725
transform 1 0 258428 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2809
timestamp 1676037725
transform 1 0 259532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2821
timestamp 1676037725
transform 1 0 260636 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2827
timestamp 1676037725
transform 1 0 261188 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2829
timestamp 1676037725
transform 1 0 261372 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2841
timestamp 1676037725
transform 1 0 262476 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2853
timestamp 1676037725
transform 1 0 263580 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2865
timestamp 1676037725
transform 1 0 264684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2877
timestamp 1676037725
transform 1 0 265788 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2883
timestamp 1676037725
transform 1 0 266340 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2885
timestamp 1676037725
transform 1 0 266524 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2897
timestamp 1676037725
transform 1 0 267628 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2909
timestamp 1676037725
transform 1 0 268732 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2921
timestamp 1676037725
transform 1 0 269836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2933
timestamp 1676037725
transform 1 0 270940 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2939
timestamp 1676037725
transform 1 0 271492 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2941
timestamp 1676037725
transform 1 0 271676 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2953
timestamp 1676037725
transform 1 0 272780 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2965
timestamp 1676037725
transform 1 0 273884 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2977
timestamp 1676037725
transform 1 0 274988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2989
timestamp 1676037725
transform 1 0 276092 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2995
timestamp 1676037725
transform 1 0 276644 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2997
timestamp 1676037725
transform 1 0 276828 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3009
timestamp 1676037725
transform 1 0 277932 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3021
timestamp 1676037725
transform 1 0 279036 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3033
timestamp 1676037725
transform 1 0 280140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3045
timestamp 1676037725
transform 1 0 281244 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3051
timestamp 1676037725
transform 1 0 281796 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3053
timestamp 1676037725
transform 1 0 281980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3065
timestamp 1676037725
transform 1 0 283084 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3077
timestamp 1676037725
transform 1 0 284188 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3089
timestamp 1676037725
transform 1 0 285292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3101
timestamp 1676037725
transform 1 0 286396 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3107
timestamp 1676037725
transform 1 0 286948 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3109
timestamp 1676037725
transform 1 0 287132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3121
timestamp 1676037725
transform 1 0 288236 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3133
timestamp 1676037725
transform 1 0 289340 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3145
timestamp 1676037725
transform 1 0 290444 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3157
timestamp 1676037725
transform 1 0 291548 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3163
timestamp 1676037725
transform 1 0 292100 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3165
timestamp 1676037725
transform 1 0 292284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3177
timestamp 1676037725
transform 1 0 293388 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3189
timestamp 1676037725
transform 1 0 294492 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3201
timestamp 1676037725
transform 1 0 295596 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3213
timestamp 1676037725
transform 1 0 296700 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3219
timestamp 1676037725
transform 1 0 297252 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3221
timestamp 1676037725
transform 1 0 297436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3233
timestamp 1676037725
transform 1 0 298540 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3245
timestamp 1676037725
transform 1 0 299644 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3257
timestamp 1676037725
transform 1 0 300748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3269
timestamp 1676037725
transform 1 0 301852 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3275
timestamp 1676037725
transform 1 0 302404 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3277
timestamp 1676037725
transform 1 0 302588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3289
timestamp 1676037725
transform 1 0 303692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3301
timestamp 1676037725
transform 1 0 304796 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3309
timestamp 1676037725
transform 1 0 305532 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3312
timestamp 1676037725
transform 1 0 305808 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3318
timestamp 1676037725
transform 1 0 306360 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3324
timestamp 1676037725
transform 1 0 306912 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3330
timestamp 1676037725
transform 1 0 307464 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3333
timestamp 1676037725
transform 1 0 307740 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3343
timestamp 1676037725
transform 1 0 308660 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3349
timestamp 1676037725
transform 1 0 309212 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3355
timestamp 1676037725
transform 1 0 309764 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3363
timestamp 1676037725
transform 1 0 310500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3375
timestamp 1676037725
transform 1 0 311604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3387
timestamp 1676037725
transform 1 0 312708 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3389
timestamp 1676037725
transform 1 0 312892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3401
timestamp 1676037725
transform 1 0 313996 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3413
timestamp 1676037725
transform 1 0 315100 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3425
timestamp 1676037725
transform 1 0 316204 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3437
timestamp 1676037725
transform 1 0 317308 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3443
timestamp 1676037725
transform 1 0 317860 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3445
timestamp 1676037725
transform 1 0 318044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3457
timestamp 1676037725
transform 1 0 319148 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3469
timestamp 1676037725
transform 1 0 320252 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3481
timestamp 1676037725
transform 1 0 321356 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3493
timestamp 1676037725
transform 1 0 322460 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3499
timestamp 1676037725
transform 1 0 323012 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3501
timestamp 1676037725
transform 1 0 323196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3513
timestamp 1676037725
transform 1 0 324300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3525
timestamp 1676037725
transform 1 0 325404 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3537
timestamp 1676037725
transform 1 0 326508 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3549
timestamp 1676037725
transform 1 0 327612 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3555
timestamp 1676037725
transform 1 0 328164 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3557
timestamp 1676037725
transform 1 0 328348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3569
timestamp 1676037725
transform 1 0 329452 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3581
timestamp 1676037725
transform 1 0 330556 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3593
timestamp 1676037725
transform 1 0 331660 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3605
timestamp 1676037725
transform 1 0 332764 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3611
timestamp 1676037725
transform 1 0 333316 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3613
timestamp 1676037725
transform 1 0 333500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3625
timestamp 1676037725
transform 1 0 334604 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3637
timestamp 1676037725
transform 1 0 335708 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3649
timestamp 1676037725
transform 1 0 336812 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3661
timestamp 1676037725
transform 1 0 337916 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3667
timestamp 1676037725
transform 1 0 338468 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3669
timestamp 1676037725
transform 1 0 338652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3681
timestamp 1676037725
transform 1 0 339756 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3693
timestamp 1676037725
transform 1 0 340860 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3705
timestamp 1676037725
transform 1 0 341964 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3717
timestamp 1676037725
transform 1 0 343068 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3723
timestamp 1676037725
transform 1 0 343620 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3725
timestamp 1676037725
transform 1 0 343804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3737
timestamp 1676037725
transform 1 0 344908 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3749
timestamp 1676037725
transform 1 0 346012 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3761
timestamp 1676037725
transform 1 0 347116 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3773
timestamp 1676037725
transform 1 0 348220 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3779
timestamp 1676037725
transform 1 0 348772 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3781
timestamp 1676037725
transform 1 0 348956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3793
timestamp 1676037725
transform 1 0 350060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3805
timestamp 1676037725
transform 1 0 351164 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3817
timestamp 1676037725
transform 1 0 352268 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3829
timestamp 1676037725
transform 1 0 353372 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3835
timestamp 1676037725
transform 1 0 353924 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3837
timestamp 1676037725
transform 1 0 354108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3849
timestamp 1676037725
transform 1 0 355212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3861
timestamp 1676037725
transform 1 0 356316 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3873
timestamp 1676037725
transform 1 0 357420 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3885
timestamp 1676037725
transform 1 0 358524 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3891
timestamp 1676037725
transform 1 0 359076 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3893
timestamp 1676037725
transform 1 0 359260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3905
timestamp 1676037725
transform 1 0 360364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3917
timestamp 1676037725
transform 1 0 361468 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3929
timestamp 1676037725
transform 1 0 362572 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3941
timestamp 1676037725
transform 1 0 363676 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3947
timestamp 1676037725
transform 1 0 364228 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3949
timestamp 1676037725
transform 1 0 364412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3961
timestamp 1676037725
transform 1 0 365516 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3973
timestamp 1676037725
transform 1 0 366620 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3985
timestamp 1676037725
transform 1 0 367724 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3997
timestamp 1676037725
transform 1 0 368828 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4003
timestamp 1676037725
transform 1 0 369380 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4005
timestamp 1676037725
transform 1 0 369564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4017
timestamp 1676037725
transform 1 0 370668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4029
timestamp 1676037725
transform 1 0 371772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4041
timestamp 1676037725
transform 1 0 372876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4053
timestamp 1676037725
transform 1 0 373980 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4059
timestamp 1676037725
transform 1 0 374532 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4061
timestamp 1676037725
transform 1 0 374716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4073
timestamp 1676037725
transform 1 0 375820 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4085
timestamp 1676037725
transform 1 0 376924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4097
timestamp 1676037725
transform 1 0 378028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4109
timestamp 1676037725
transform 1 0 379132 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4115
timestamp 1676037725
transform 1 0 379684 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4117
timestamp 1676037725
transform 1 0 379868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4129
timestamp 1676037725
transform 1 0 380972 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4141
timestamp 1676037725
transform 1 0 382076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4153
timestamp 1676037725
transform 1 0 383180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4165
timestamp 1676037725
transform 1 0 384284 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4171
timestamp 1676037725
transform 1 0 384836 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4173
timestamp 1676037725
transform 1 0 385020 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4185
timestamp 1676037725
transform 1 0 386124 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4197
timestamp 1676037725
transform 1 0 387228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4209
timestamp 1676037725
transform 1 0 388332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4221
timestamp 1676037725
transform 1 0 389436 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4227
timestamp 1676037725
transform 1 0 389988 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4229
timestamp 1676037725
transform 1 0 390172 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4241
timestamp 1676037725
transform 1 0 391276 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4253
timestamp 1676037725
transform 1 0 392380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4265
timestamp 1676037725
transform 1 0 393484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4277
timestamp 1676037725
transform 1 0 394588 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4283
timestamp 1676037725
transform 1 0 395140 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4285
timestamp 1676037725
transform 1 0 395324 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4297
timestamp 1676037725
transform 1 0 396428 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4309
timestamp 1676037725
transform 1 0 397532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4321
timestamp 1676037725
transform 1 0 398636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4333
timestamp 1676037725
transform 1 0 399740 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4339
timestamp 1676037725
transform 1 0 400292 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4341
timestamp 1676037725
transform 1 0 400476 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4353
timestamp 1676037725
transform 1 0 401580 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4365
timestamp 1676037725
transform 1 0 402684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4377
timestamp 1676037725
transform 1 0 403788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4389
timestamp 1676037725
transform 1 0 404892 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4395
timestamp 1676037725
transform 1 0 405444 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4397
timestamp 1676037725
transform 1 0 405628 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4409
timestamp 1676037725
transform 1 0 406732 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4421
timestamp 1676037725
transform 1 0 407836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4433
timestamp 1676037725
transform 1 0 408940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4445
timestamp 1676037725
transform 1 0 410044 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4451
timestamp 1676037725
transform 1 0 410596 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4453
timestamp 1676037725
transform 1 0 410780 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4465
timestamp 1676037725
transform 1 0 411884 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4477
timestamp 1676037725
transform 1 0 412988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4489
timestamp 1676037725
transform 1 0 414092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4501
timestamp 1676037725
transform 1 0 415196 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4507
timestamp 1676037725
transform 1 0 415748 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4509
timestamp 1676037725
transform 1 0 415932 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4521
timestamp 1676037725
transform 1 0 417036 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4533
timestamp 1676037725
transform 1 0 418140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4545
timestamp 1676037725
transform 1 0 419244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4557
timestamp 1676037725
transform 1 0 420348 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4563
timestamp 1676037725
transform 1 0 420900 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4565
timestamp 1676037725
transform 1 0 421084 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4577
timestamp 1676037725
transform 1 0 422188 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4589
timestamp 1676037725
transform 1 0 423292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4601
timestamp 1676037725
transform 1 0 424396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4613
timestamp 1676037725
transform 1 0 425500 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4619
timestamp 1676037725
transform 1 0 426052 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4621
timestamp 1676037725
transform 1 0 426236 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4633
timestamp 1676037725
transform 1 0 427340 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4645
timestamp 1676037725
transform 1 0 428444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4657
timestamp 1676037725
transform 1 0 429548 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4669
timestamp 1676037725
transform 1 0 430652 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4675
timestamp 1676037725
transform 1 0 431204 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4677
timestamp 1676037725
transform 1 0 431388 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4689
timestamp 1676037725
transform 1 0 432492 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4701
timestamp 1676037725
transform 1 0 433596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4713
timestamp 1676037725
transform 1 0 434700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4725
timestamp 1676037725
transform 1 0 435804 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4731
timestamp 1676037725
transform 1 0 436356 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4733
timestamp 1676037725
transform 1 0 436540 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4745
timestamp 1676037725
transform 1 0 437644 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4757
timestamp 1676037725
transform 1 0 438748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4769
timestamp 1676037725
transform 1 0 439852 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4781
timestamp 1676037725
transform 1 0 440956 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4787
timestamp 1676037725
transform 1 0 441508 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4789
timestamp 1676037725
transform 1 0 441692 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4801
timestamp 1676037725
transform 1 0 442796 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4813
timestamp 1676037725
transform 1 0 443900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4825
timestamp 1676037725
transform 1 0 445004 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4837
timestamp 1676037725
transform 1 0 446108 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4843
timestamp 1676037725
transform 1 0 446660 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4845
timestamp 1676037725
transform 1 0 446844 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4857
timestamp 1676037725
transform 1 0 447948 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4869
timestamp 1676037725
transform 1 0 449052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4881
timestamp 1676037725
transform 1 0 450156 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4893
timestamp 1676037725
transform 1 0 451260 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4899
timestamp 1676037725
transform 1 0 451812 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4901
timestamp 1676037725
transform 1 0 451996 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4913
timestamp 1676037725
transform 1 0 453100 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4925
timestamp 1676037725
transform 1 0 454204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4937
timestamp 1676037725
transform 1 0 455308 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4949
timestamp 1676037725
transform 1 0 456412 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4955
timestamp 1676037725
transform 1 0 456964 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4957
timestamp 1676037725
transform 1 0 457148 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4969
timestamp 1676037725
transform 1 0 458252 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4981
timestamp 1676037725
transform 1 0 459356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4993
timestamp 1676037725
transform 1 0 460460 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5005
timestamp 1676037725
transform 1 0 461564 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5011
timestamp 1676037725
transform 1 0 462116 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5013
timestamp 1676037725
transform 1 0 462300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5025
timestamp 1676037725
transform 1 0 463404 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5037
timestamp 1676037725
transform 1 0 464508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5049
timestamp 1676037725
transform 1 0 465612 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5061
timestamp 1676037725
transform 1 0 466716 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5067
timestamp 1676037725
transform 1 0 467268 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5069
timestamp 1676037725
transform 1 0 467452 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5081
timestamp 1676037725
transform 1 0 468556 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5093
timestamp 1676037725
transform 1 0 469660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5105
timestamp 1676037725
transform 1 0 470764 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5117
timestamp 1676037725
transform 1 0 471868 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5123
timestamp 1676037725
transform 1 0 472420 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5125
timestamp 1676037725
transform 1 0 472604 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5137
timestamp 1676037725
transform 1 0 473708 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5149
timestamp 1676037725
transform 1 0 474812 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5161
timestamp 1676037725
transform 1 0 475916 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5173
timestamp 1676037725
transform 1 0 477020 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5179
timestamp 1676037725
transform 1 0 477572 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5181
timestamp 1676037725
transform 1 0 477756 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5193
timestamp 1676037725
transform 1 0 478860 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5205
timestamp 1676037725
transform 1 0 479964 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5217
timestamp 1676037725
transform 1 0 481068 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5229
timestamp 1676037725
transform 1 0 482172 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5235
timestamp 1676037725
transform 1 0 482724 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5237
timestamp 1676037725
transform 1 0 482908 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5249
timestamp 1676037725
transform 1 0 484012 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5261
timestamp 1676037725
transform 1 0 485116 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5273
timestamp 1676037725
transform 1 0 486220 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5285
timestamp 1676037725
transform 1 0 487324 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5291
timestamp 1676037725
transform 1 0 487876 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5293
timestamp 1676037725
transform 1 0 488060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5305
timestamp 1676037725
transform 1 0 489164 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5317
timestamp 1676037725
transform 1 0 490268 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5329
timestamp 1676037725
transform 1 0 491372 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5341
timestamp 1676037725
transform 1 0 492476 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5347
timestamp 1676037725
transform 1 0 493028 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5349
timestamp 1676037725
transform 1 0 493212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5361
timestamp 1676037725
transform 1 0 494316 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5373
timestamp 1676037725
transform 1 0 495420 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5385
timestamp 1676037725
transform 1 0 496524 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5397
timestamp 1676037725
transform 1 0 497628 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5403
timestamp 1676037725
transform 1 0 498180 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5405
timestamp 1676037725
transform 1 0 498364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5417
timestamp 1676037725
transform 1 0 499468 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5429
timestamp 1676037725
transform 1 0 500572 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5441
timestamp 1676037725
transform 1 0 501676 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5453
timestamp 1676037725
transform 1 0 502780 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5459
timestamp 1676037725
transform 1 0 503332 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5461
timestamp 1676037725
transform 1 0 503516 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5473
timestamp 1676037725
transform 1 0 504620 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5485
timestamp 1676037725
transform 1 0 505724 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5497
timestamp 1676037725
transform 1 0 506828 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5509
timestamp 1676037725
transform 1 0 507932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5515
timestamp 1676037725
transform 1 0 508484 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5517
timestamp 1676037725
transform 1 0 508668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5529
timestamp 1676037725
transform 1 0 509772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5541
timestamp 1676037725
transform 1 0 510876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5553
timestamp 1676037725
transform 1 0 511980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5565
timestamp 1676037725
transform 1 0 513084 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5571
timestamp 1676037725
transform 1 0 513636 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5573
timestamp 1676037725
transform 1 0 513820 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5585
timestamp 1676037725
transform 1 0 514924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5597
timestamp 1676037725
transform 1 0 516028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5609
timestamp 1676037725
transform 1 0 517132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5621
timestamp 1676037725
transform 1 0 518236 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5627
timestamp 1676037725
transform 1 0 518788 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5629
timestamp 1676037725
transform 1 0 518972 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5641
timestamp 1676037725
transform 1 0 520076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5653
timestamp 1676037725
transform 1 0 521180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5665
timestamp 1676037725
transform 1 0 522284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5677
timestamp 1676037725
transform 1 0 523388 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5683
timestamp 1676037725
transform 1 0 523940 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5685
timestamp 1676037725
transform 1 0 524124 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5697
timestamp 1676037725
transform 1 0 525228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5709
timestamp 1676037725
transform 1 0 526332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5721
timestamp 1676037725
transform 1 0 527436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1676037725
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1676037725
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1676037725
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1676037725
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1676037725
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1676037725
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1676037725
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1676037725
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1676037725
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1676037725
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1676037725
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1676037725
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1676037725
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1676037725
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1676037725
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1676037725
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1676037725
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1676037725
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1676037725
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1676037725
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1676037725
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1676037725
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1676037725
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1676037725
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1676037725
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1676037725
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1676037725
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1676037725
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1676037725
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1676037725
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1676037725
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1676037725
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1676037725
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1676037725
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1676037725
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1676037725
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 1676037725
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1676037725
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1676037725
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1676037725
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_809
timestamp 1676037725
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_821
timestamp 1676037725
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_833
timestamp 1676037725
transform 1 0 77740 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_839
timestamp 1676037725
transform 1 0 78292 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_841
timestamp 1676037725
transform 1 0 78476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_853
timestamp 1676037725
transform 1 0 79580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_865
timestamp 1676037725
transform 1 0 80684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_877
timestamp 1676037725
transform 1 0 81788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_889
timestamp 1676037725
transform 1 0 82892 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_895
timestamp 1676037725
transform 1 0 83444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_897
timestamp 1676037725
transform 1 0 83628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_909
timestamp 1676037725
transform 1 0 84732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_921
timestamp 1676037725
transform 1 0 85836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_933
timestamp 1676037725
transform 1 0 86940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_945
timestamp 1676037725
transform 1 0 88044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_951
timestamp 1676037725
transform 1 0 88596 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_953
timestamp 1676037725
transform 1 0 88780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_965
timestamp 1676037725
transform 1 0 89884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_977
timestamp 1676037725
transform 1 0 90988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_989
timestamp 1676037725
transform 1 0 92092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1001
timestamp 1676037725
transform 1 0 93196 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1007
timestamp 1676037725
transform 1 0 93748 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1009
timestamp 1676037725
transform 1 0 93932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1021
timestamp 1676037725
transform 1 0 95036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1033
timestamp 1676037725
transform 1 0 96140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1045
timestamp 1676037725
transform 1 0 97244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1057
timestamp 1676037725
transform 1 0 98348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1063
timestamp 1676037725
transform 1 0 98900 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1065
timestamp 1676037725
transform 1 0 99084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1077
timestamp 1676037725
transform 1 0 100188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1089
timestamp 1676037725
transform 1 0 101292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1101
timestamp 1676037725
transform 1 0 102396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1113
timestamp 1676037725
transform 1 0 103500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1119
timestamp 1676037725
transform 1 0 104052 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1121
timestamp 1676037725
transform 1 0 104236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1133
timestamp 1676037725
transform 1 0 105340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1145
timestamp 1676037725
transform 1 0 106444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1157
timestamp 1676037725
transform 1 0 107548 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1169
timestamp 1676037725
transform 1 0 108652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1175
timestamp 1676037725
transform 1 0 109204 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1177
timestamp 1676037725
transform 1 0 109388 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1189
timestamp 1676037725
transform 1 0 110492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1201
timestamp 1676037725
transform 1 0 111596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1213
timestamp 1676037725
transform 1 0 112700 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1225
timestamp 1676037725
transform 1 0 113804 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1231
timestamp 1676037725
transform 1 0 114356 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1233
timestamp 1676037725
transform 1 0 114540 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1245
timestamp 1676037725
transform 1 0 115644 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1253
timestamp 1676037725
transform 1 0 116380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1257
timestamp 1676037725
transform 1 0 116748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1260
timestamp 1676037725
transform 1 0 117024 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1266
timestamp 1676037725
transform 1 0 117576 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1272
timestamp 1676037725
transform 1 0 118128 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1275
timestamp 1676037725
transform 1 0 118404 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1287
timestamp 1676037725
transform 1 0 119508 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1289
timestamp 1676037725
transform 1 0 119692 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1301
timestamp 1676037725
transform 1 0 120796 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1313
timestamp 1676037725
transform 1 0 121900 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1325
timestamp 1676037725
transform 1 0 123004 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1337
timestamp 1676037725
transform 1 0 124108 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1343
timestamp 1676037725
transform 1 0 124660 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1345
timestamp 1676037725
transform 1 0 124844 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1357
timestamp 1676037725
transform 1 0 125948 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1369
timestamp 1676037725
transform 1 0 127052 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1381
timestamp 1676037725
transform 1 0 128156 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1393
timestamp 1676037725
transform 1 0 129260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1399
timestamp 1676037725
transform 1 0 129812 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1401
timestamp 1676037725
transform 1 0 129996 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1413
timestamp 1676037725
transform 1 0 131100 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1425
timestamp 1676037725
transform 1 0 132204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1437
timestamp 1676037725
transform 1 0 133308 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1449
timestamp 1676037725
transform 1 0 134412 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1455
timestamp 1676037725
transform 1 0 134964 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1457
timestamp 1676037725
transform 1 0 135148 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1469
timestamp 1676037725
transform 1 0 136252 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1481
timestamp 1676037725
transform 1 0 137356 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1493
timestamp 1676037725
transform 1 0 138460 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1505
timestamp 1676037725
transform 1 0 139564 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1511
timestamp 1676037725
transform 1 0 140116 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1513
timestamp 1676037725
transform 1 0 140300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1525
timestamp 1676037725
transform 1 0 141404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1537
timestamp 1676037725
transform 1 0 142508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1549
timestamp 1676037725
transform 1 0 143612 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1561
timestamp 1676037725
transform 1 0 144716 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1567
timestamp 1676037725
transform 1 0 145268 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1569
timestamp 1676037725
transform 1 0 145452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1581
timestamp 1676037725
transform 1 0 146556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1593
timestamp 1676037725
transform 1 0 147660 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1605
timestamp 1676037725
transform 1 0 148764 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1617
timestamp 1676037725
transform 1 0 149868 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1623
timestamp 1676037725
transform 1 0 150420 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1625
timestamp 1676037725
transform 1 0 150604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1637
timestamp 1676037725
transform 1 0 151708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1649
timestamp 1676037725
transform 1 0 152812 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1661
timestamp 1676037725
transform 1 0 153916 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1673
timestamp 1676037725
transform 1 0 155020 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1679
timestamp 1676037725
transform 1 0 155572 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1681
timestamp 1676037725
transform 1 0 155756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1693
timestamp 1676037725
transform 1 0 156860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1705
timestamp 1676037725
transform 1 0 157964 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1717
timestamp 1676037725
transform 1 0 159068 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1729
timestamp 1676037725
transform 1 0 160172 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1735
timestamp 1676037725
transform 1 0 160724 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1737
timestamp 1676037725
transform 1 0 160908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1749
timestamp 1676037725
transform 1 0 162012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1761
timestamp 1676037725
transform 1 0 163116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1773
timestamp 1676037725
transform 1 0 164220 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1785
timestamp 1676037725
transform 1 0 165324 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1791
timestamp 1676037725
transform 1 0 165876 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1793
timestamp 1676037725
transform 1 0 166060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1805
timestamp 1676037725
transform 1 0 167164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1817
timestamp 1676037725
transform 1 0 168268 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1829
timestamp 1676037725
transform 1 0 169372 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1841
timestamp 1676037725
transform 1 0 170476 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1847
timestamp 1676037725
transform 1 0 171028 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1849
timestamp 1676037725
transform 1 0 171212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1861
timestamp 1676037725
transform 1 0 172316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1873
timestamp 1676037725
transform 1 0 173420 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1885
timestamp 1676037725
transform 1 0 174524 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1897
timestamp 1676037725
transform 1 0 175628 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1903
timestamp 1676037725
transform 1 0 176180 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1905
timestamp 1676037725
transform 1 0 176364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1917
timestamp 1676037725
transform 1 0 177468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1929
timestamp 1676037725
transform 1 0 178572 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1941
timestamp 1676037725
transform 1 0 179676 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1953
timestamp 1676037725
transform 1 0 180780 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1959
timestamp 1676037725
transform 1 0 181332 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1961
timestamp 1676037725
transform 1 0 181516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1973
timestamp 1676037725
transform 1 0 182620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1985
timestamp 1676037725
transform 1 0 183724 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1997
timestamp 1676037725
transform 1 0 184828 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2009
timestamp 1676037725
transform 1 0 185932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2015
timestamp 1676037725
transform 1 0 186484 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2017
timestamp 1676037725
transform 1 0 186668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2029
timestamp 1676037725
transform 1 0 187772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2041
timestamp 1676037725
transform 1 0 188876 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2053
timestamp 1676037725
transform 1 0 189980 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2065
timestamp 1676037725
transform 1 0 191084 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2071
timestamp 1676037725
transform 1 0 191636 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2073
timestamp 1676037725
transform 1 0 191820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2085
timestamp 1676037725
transform 1 0 192924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2097
timestamp 1676037725
transform 1 0 194028 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2109
timestamp 1676037725
transform 1 0 195132 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2121
timestamp 1676037725
transform 1 0 196236 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2127
timestamp 1676037725
transform 1 0 196788 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2129
timestamp 1676037725
transform 1 0 196972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2141
timestamp 1676037725
transform 1 0 198076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2153
timestamp 1676037725
transform 1 0 199180 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2165
timestamp 1676037725
transform 1 0 200284 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2177
timestamp 1676037725
transform 1 0 201388 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2183
timestamp 1676037725
transform 1 0 201940 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2185
timestamp 1676037725
transform 1 0 202124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2197
timestamp 1676037725
transform 1 0 203228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2209
timestamp 1676037725
transform 1 0 204332 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2221
timestamp 1676037725
transform 1 0 205436 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2233
timestamp 1676037725
transform 1 0 206540 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2239
timestamp 1676037725
transform 1 0 207092 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2241
timestamp 1676037725
transform 1 0 207276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2253
timestamp 1676037725
transform 1 0 208380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2265
timestamp 1676037725
transform 1 0 209484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_2277
timestamp 1676037725
transform 1 0 210588 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_2283
timestamp 1676037725
transform 1 0 211140 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2289
timestamp 1676037725
transform 1 0 211692 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2295
timestamp 1676037725
transform 1 0 212244 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2297
timestamp 1676037725
transform 1 0 212428 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_2311
timestamp 1676037725
transform 1 0 213716 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2315
timestamp 1676037725
transform 1 0 214084 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_2318
timestamp 1676037725
transform 1 0 214360 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_2324
timestamp 1676037725
transform 1 0 214912 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2330
timestamp 1676037725
transform 1 0 215464 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2336
timestamp 1676037725
transform 1 0 216016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_2339
timestamp 1676037725
transform 1 0 216292 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2345
timestamp 1676037725
transform 1 0 216844 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2351
timestamp 1676037725
transform 1 0 217396 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2353
timestamp 1676037725
transform 1 0 217580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2365
timestamp 1676037725
transform 1 0 218684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2377
timestamp 1676037725
transform 1 0 219788 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2389
timestamp 1676037725
transform 1 0 220892 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2401
timestamp 1676037725
transform 1 0 221996 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2407
timestamp 1676037725
transform 1 0 222548 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2409
timestamp 1676037725
transform 1 0 222732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2421
timestamp 1676037725
transform 1 0 223836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2433
timestamp 1676037725
transform 1 0 224940 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2445
timestamp 1676037725
transform 1 0 226044 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2457
timestamp 1676037725
transform 1 0 227148 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2463
timestamp 1676037725
transform 1 0 227700 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2465
timestamp 1676037725
transform 1 0 227884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2477
timestamp 1676037725
transform 1 0 228988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2489
timestamp 1676037725
transform 1 0 230092 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2501
timestamp 1676037725
transform 1 0 231196 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2513
timestamp 1676037725
transform 1 0 232300 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2519
timestamp 1676037725
transform 1 0 232852 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2521
timestamp 1676037725
transform 1 0 233036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2533
timestamp 1676037725
transform 1 0 234140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2545
timestamp 1676037725
transform 1 0 235244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2557
timestamp 1676037725
transform 1 0 236348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2569
timestamp 1676037725
transform 1 0 237452 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2575
timestamp 1676037725
transform 1 0 238004 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2577
timestamp 1676037725
transform 1 0 238188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2589
timestamp 1676037725
transform 1 0 239292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2601
timestamp 1676037725
transform 1 0 240396 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2613
timestamp 1676037725
transform 1 0 241500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2625
timestamp 1676037725
transform 1 0 242604 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2631
timestamp 1676037725
transform 1 0 243156 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2633
timestamp 1676037725
transform 1 0 243340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2645
timestamp 1676037725
transform 1 0 244444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2657
timestamp 1676037725
transform 1 0 245548 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2669
timestamp 1676037725
transform 1 0 246652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2681
timestamp 1676037725
transform 1 0 247756 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2687
timestamp 1676037725
transform 1 0 248308 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2689
timestamp 1676037725
transform 1 0 248492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2701
timestamp 1676037725
transform 1 0 249596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2713
timestamp 1676037725
transform 1 0 250700 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2725
timestamp 1676037725
transform 1 0 251804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2737
timestamp 1676037725
transform 1 0 252908 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2743
timestamp 1676037725
transform 1 0 253460 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2745
timestamp 1676037725
transform 1 0 253644 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2757
timestamp 1676037725
transform 1 0 254748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2769
timestamp 1676037725
transform 1 0 255852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2781
timestamp 1676037725
transform 1 0 256956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2793
timestamp 1676037725
transform 1 0 258060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2799
timestamp 1676037725
transform 1 0 258612 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2801
timestamp 1676037725
transform 1 0 258796 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2813
timestamp 1676037725
transform 1 0 259900 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2825
timestamp 1676037725
transform 1 0 261004 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2837
timestamp 1676037725
transform 1 0 262108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2849
timestamp 1676037725
transform 1 0 263212 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2855
timestamp 1676037725
transform 1 0 263764 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2857
timestamp 1676037725
transform 1 0 263948 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2869
timestamp 1676037725
transform 1 0 265052 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2881
timestamp 1676037725
transform 1 0 266156 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2893
timestamp 1676037725
transform 1 0 267260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2905
timestamp 1676037725
transform 1 0 268364 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2911
timestamp 1676037725
transform 1 0 268916 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2913
timestamp 1676037725
transform 1 0 269100 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2925
timestamp 1676037725
transform 1 0 270204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2937
timestamp 1676037725
transform 1 0 271308 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2949
timestamp 1676037725
transform 1 0 272412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2961
timestamp 1676037725
transform 1 0 273516 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2967
timestamp 1676037725
transform 1 0 274068 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2969
timestamp 1676037725
transform 1 0 274252 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2981
timestamp 1676037725
transform 1 0 275356 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2993
timestamp 1676037725
transform 1 0 276460 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3005
timestamp 1676037725
transform 1 0 277564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3017
timestamp 1676037725
transform 1 0 278668 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3023
timestamp 1676037725
transform 1 0 279220 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3025
timestamp 1676037725
transform 1 0 279404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3037
timestamp 1676037725
transform 1 0 280508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3049
timestamp 1676037725
transform 1 0 281612 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3061
timestamp 1676037725
transform 1 0 282716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3073
timestamp 1676037725
transform 1 0 283820 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3079
timestamp 1676037725
transform 1 0 284372 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3081
timestamp 1676037725
transform 1 0 284556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3093
timestamp 1676037725
transform 1 0 285660 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3105
timestamp 1676037725
transform 1 0 286764 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3117
timestamp 1676037725
transform 1 0 287868 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3129
timestamp 1676037725
transform 1 0 288972 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3135
timestamp 1676037725
transform 1 0 289524 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3137
timestamp 1676037725
transform 1 0 289708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3149
timestamp 1676037725
transform 1 0 290812 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3161
timestamp 1676037725
transform 1 0 291916 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3173
timestamp 1676037725
transform 1 0 293020 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3185
timestamp 1676037725
transform 1 0 294124 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3191
timestamp 1676037725
transform 1 0 294676 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3193
timestamp 1676037725
transform 1 0 294860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3205
timestamp 1676037725
transform 1 0 295964 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3217
timestamp 1676037725
transform 1 0 297068 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3229
timestamp 1676037725
transform 1 0 298172 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3241
timestamp 1676037725
transform 1 0 299276 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3247
timestamp 1676037725
transform 1 0 299828 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3249
timestamp 1676037725
transform 1 0 300012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3261
timestamp 1676037725
transform 1 0 301116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3273
timestamp 1676037725
transform 1 0 302220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3285
timestamp 1676037725
transform 1 0 303324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3297
timestamp 1676037725
transform 1 0 304428 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3303
timestamp 1676037725
transform 1 0 304980 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3305
timestamp 1676037725
transform 1 0 305164 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3313
timestamp 1676037725
transform 1 0 305900 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3318
timestamp 1676037725
transform 1 0 306360 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3324
timestamp 1676037725
transform 1 0 306912 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3332
timestamp 1676037725
transform 1 0 307648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3338
timestamp 1676037725
transform 1 0 308200 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3342
timestamp 1676037725
transform 1 0 308568 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3345
timestamp 1676037725
transform 1 0 308844 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3357
timestamp 1676037725
transform 1 0 309948 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3361
timestamp 1676037725
transform 1 0 310316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3373
timestamp 1676037725
transform 1 0 311420 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3385
timestamp 1676037725
transform 1 0 312524 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3397
timestamp 1676037725
transform 1 0 313628 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3409
timestamp 1676037725
transform 1 0 314732 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3415
timestamp 1676037725
transform 1 0 315284 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3417
timestamp 1676037725
transform 1 0 315468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3429
timestamp 1676037725
transform 1 0 316572 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3441
timestamp 1676037725
transform 1 0 317676 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3453
timestamp 1676037725
transform 1 0 318780 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3465
timestamp 1676037725
transform 1 0 319884 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3471
timestamp 1676037725
transform 1 0 320436 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3473
timestamp 1676037725
transform 1 0 320620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3485
timestamp 1676037725
transform 1 0 321724 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3497
timestamp 1676037725
transform 1 0 322828 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3509
timestamp 1676037725
transform 1 0 323932 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3521
timestamp 1676037725
transform 1 0 325036 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3527
timestamp 1676037725
transform 1 0 325588 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3529
timestamp 1676037725
transform 1 0 325772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3541
timestamp 1676037725
transform 1 0 326876 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3553
timestamp 1676037725
transform 1 0 327980 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3565
timestamp 1676037725
transform 1 0 329084 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3577
timestamp 1676037725
transform 1 0 330188 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3583
timestamp 1676037725
transform 1 0 330740 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3585
timestamp 1676037725
transform 1 0 330924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3597
timestamp 1676037725
transform 1 0 332028 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3609
timestamp 1676037725
transform 1 0 333132 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3621
timestamp 1676037725
transform 1 0 334236 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3633
timestamp 1676037725
transform 1 0 335340 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3639
timestamp 1676037725
transform 1 0 335892 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3641
timestamp 1676037725
transform 1 0 336076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3653
timestamp 1676037725
transform 1 0 337180 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3665
timestamp 1676037725
transform 1 0 338284 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3677
timestamp 1676037725
transform 1 0 339388 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3689
timestamp 1676037725
transform 1 0 340492 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3695
timestamp 1676037725
transform 1 0 341044 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3697
timestamp 1676037725
transform 1 0 341228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3709
timestamp 1676037725
transform 1 0 342332 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3721
timestamp 1676037725
transform 1 0 343436 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3733
timestamp 1676037725
transform 1 0 344540 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3745
timestamp 1676037725
transform 1 0 345644 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3751
timestamp 1676037725
transform 1 0 346196 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3753
timestamp 1676037725
transform 1 0 346380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3765
timestamp 1676037725
transform 1 0 347484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3777
timestamp 1676037725
transform 1 0 348588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3789
timestamp 1676037725
transform 1 0 349692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3801
timestamp 1676037725
transform 1 0 350796 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3807
timestamp 1676037725
transform 1 0 351348 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3809
timestamp 1676037725
transform 1 0 351532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3821
timestamp 1676037725
transform 1 0 352636 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3833
timestamp 1676037725
transform 1 0 353740 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3845
timestamp 1676037725
transform 1 0 354844 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3857
timestamp 1676037725
transform 1 0 355948 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3863
timestamp 1676037725
transform 1 0 356500 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3865
timestamp 1676037725
transform 1 0 356684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3877
timestamp 1676037725
transform 1 0 357788 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3889
timestamp 1676037725
transform 1 0 358892 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3901
timestamp 1676037725
transform 1 0 359996 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3913
timestamp 1676037725
transform 1 0 361100 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3919
timestamp 1676037725
transform 1 0 361652 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3921
timestamp 1676037725
transform 1 0 361836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3933
timestamp 1676037725
transform 1 0 362940 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3945
timestamp 1676037725
transform 1 0 364044 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3957
timestamp 1676037725
transform 1 0 365148 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3969
timestamp 1676037725
transform 1 0 366252 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3975
timestamp 1676037725
transform 1 0 366804 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3977
timestamp 1676037725
transform 1 0 366988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3989
timestamp 1676037725
transform 1 0 368092 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4001
timestamp 1676037725
transform 1 0 369196 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4013
timestamp 1676037725
transform 1 0 370300 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4025
timestamp 1676037725
transform 1 0 371404 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4031
timestamp 1676037725
transform 1 0 371956 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4033
timestamp 1676037725
transform 1 0 372140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4045
timestamp 1676037725
transform 1 0 373244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4057
timestamp 1676037725
transform 1 0 374348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4069
timestamp 1676037725
transform 1 0 375452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4081
timestamp 1676037725
transform 1 0 376556 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4087
timestamp 1676037725
transform 1 0 377108 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4089
timestamp 1676037725
transform 1 0 377292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4101
timestamp 1676037725
transform 1 0 378396 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4113
timestamp 1676037725
transform 1 0 379500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4125
timestamp 1676037725
transform 1 0 380604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4137
timestamp 1676037725
transform 1 0 381708 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4143
timestamp 1676037725
transform 1 0 382260 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4145
timestamp 1676037725
transform 1 0 382444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4157
timestamp 1676037725
transform 1 0 383548 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4169
timestamp 1676037725
transform 1 0 384652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4181
timestamp 1676037725
transform 1 0 385756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4193
timestamp 1676037725
transform 1 0 386860 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4199
timestamp 1676037725
transform 1 0 387412 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4201
timestamp 1676037725
transform 1 0 387596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4213
timestamp 1676037725
transform 1 0 388700 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4225
timestamp 1676037725
transform 1 0 389804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4237
timestamp 1676037725
transform 1 0 390908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4249
timestamp 1676037725
transform 1 0 392012 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4255
timestamp 1676037725
transform 1 0 392564 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4257
timestamp 1676037725
transform 1 0 392748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4269
timestamp 1676037725
transform 1 0 393852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4281
timestamp 1676037725
transform 1 0 394956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4293
timestamp 1676037725
transform 1 0 396060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4305
timestamp 1676037725
transform 1 0 397164 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4311
timestamp 1676037725
transform 1 0 397716 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4313
timestamp 1676037725
transform 1 0 397900 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4325
timestamp 1676037725
transform 1 0 399004 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4337
timestamp 1676037725
transform 1 0 400108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4349
timestamp 1676037725
transform 1 0 401212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4361
timestamp 1676037725
transform 1 0 402316 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4367
timestamp 1676037725
transform 1 0 402868 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4369
timestamp 1676037725
transform 1 0 403052 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4381
timestamp 1676037725
transform 1 0 404156 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4393
timestamp 1676037725
transform 1 0 405260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4405
timestamp 1676037725
transform 1 0 406364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4417
timestamp 1676037725
transform 1 0 407468 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4423
timestamp 1676037725
transform 1 0 408020 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4425
timestamp 1676037725
transform 1 0 408204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4437
timestamp 1676037725
transform 1 0 409308 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4449
timestamp 1676037725
transform 1 0 410412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4461
timestamp 1676037725
transform 1 0 411516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4473
timestamp 1676037725
transform 1 0 412620 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4479
timestamp 1676037725
transform 1 0 413172 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4481
timestamp 1676037725
transform 1 0 413356 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4493
timestamp 1676037725
transform 1 0 414460 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4505
timestamp 1676037725
transform 1 0 415564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4517
timestamp 1676037725
transform 1 0 416668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4529
timestamp 1676037725
transform 1 0 417772 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4535
timestamp 1676037725
transform 1 0 418324 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4537
timestamp 1676037725
transform 1 0 418508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4549
timestamp 1676037725
transform 1 0 419612 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4561
timestamp 1676037725
transform 1 0 420716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4573
timestamp 1676037725
transform 1 0 421820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4585
timestamp 1676037725
transform 1 0 422924 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4591
timestamp 1676037725
transform 1 0 423476 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4593
timestamp 1676037725
transform 1 0 423660 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4605
timestamp 1676037725
transform 1 0 424764 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4617
timestamp 1676037725
transform 1 0 425868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4629
timestamp 1676037725
transform 1 0 426972 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4641
timestamp 1676037725
transform 1 0 428076 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4647
timestamp 1676037725
transform 1 0 428628 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4649
timestamp 1676037725
transform 1 0 428812 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4661
timestamp 1676037725
transform 1 0 429916 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4673
timestamp 1676037725
transform 1 0 431020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4685
timestamp 1676037725
transform 1 0 432124 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4697
timestamp 1676037725
transform 1 0 433228 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4703
timestamp 1676037725
transform 1 0 433780 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4705
timestamp 1676037725
transform 1 0 433964 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4717
timestamp 1676037725
transform 1 0 435068 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4729
timestamp 1676037725
transform 1 0 436172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4741
timestamp 1676037725
transform 1 0 437276 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4753
timestamp 1676037725
transform 1 0 438380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4759
timestamp 1676037725
transform 1 0 438932 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4761
timestamp 1676037725
transform 1 0 439116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4773
timestamp 1676037725
transform 1 0 440220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4785
timestamp 1676037725
transform 1 0 441324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4797
timestamp 1676037725
transform 1 0 442428 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4809
timestamp 1676037725
transform 1 0 443532 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4815
timestamp 1676037725
transform 1 0 444084 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4817
timestamp 1676037725
transform 1 0 444268 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4829
timestamp 1676037725
transform 1 0 445372 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4841
timestamp 1676037725
transform 1 0 446476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4853
timestamp 1676037725
transform 1 0 447580 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4865
timestamp 1676037725
transform 1 0 448684 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4871
timestamp 1676037725
transform 1 0 449236 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4873
timestamp 1676037725
transform 1 0 449420 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4885
timestamp 1676037725
transform 1 0 450524 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4897
timestamp 1676037725
transform 1 0 451628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4909
timestamp 1676037725
transform 1 0 452732 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4921
timestamp 1676037725
transform 1 0 453836 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4927
timestamp 1676037725
transform 1 0 454388 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4929
timestamp 1676037725
transform 1 0 454572 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4941
timestamp 1676037725
transform 1 0 455676 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4953
timestamp 1676037725
transform 1 0 456780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4965
timestamp 1676037725
transform 1 0 457884 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4977
timestamp 1676037725
transform 1 0 458988 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4983
timestamp 1676037725
transform 1 0 459540 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4985
timestamp 1676037725
transform 1 0 459724 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4997
timestamp 1676037725
transform 1 0 460828 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5009
timestamp 1676037725
transform 1 0 461932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5021
timestamp 1676037725
transform 1 0 463036 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5033
timestamp 1676037725
transform 1 0 464140 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5039
timestamp 1676037725
transform 1 0 464692 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5041
timestamp 1676037725
transform 1 0 464876 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5053
timestamp 1676037725
transform 1 0 465980 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5065
timestamp 1676037725
transform 1 0 467084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5077
timestamp 1676037725
transform 1 0 468188 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5089
timestamp 1676037725
transform 1 0 469292 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5095
timestamp 1676037725
transform 1 0 469844 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5097
timestamp 1676037725
transform 1 0 470028 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5109
timestamp 1676037725
transform 1 0 471132 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5121
timestamp 1676037725
transform 1 0 472236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5133
timestamp 1676037725
transform 1 0 473340 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5145
timestamp 1676037725
transform 1 0 474444 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5151
timestamp 1676037725
transform 1 0 474996 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5153
timestamp 1676037725
transform 1 0 475180 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5165
timestamp 1676037725
transform 1 0 476284 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5177
timestamp 1676037725
transform 1 0 477388 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5189
timestamp 1676037725
transform 1 0 478492 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5201
timestamp 1676037725
transform 1 0 479596 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5207
timestamp 1676037725
transform 1 0 480148 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5209
timestamp 1676037725
transform 1 0 480332 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5221
timestamp 1676037725
transform 1 0 481436 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5233
timestamp 1676037725
transform 1 0 482540 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5245
timestamp 1676037725
transform 1 0 483644 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5257
timestamp 1676037725
transform 1 0 484748 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5263
timestamp 1676037725
transform 1 0 485300 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5265
timestamp 1676037725
transform 1 0 485484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5277
timestamp 1676037725
transform 1 0 486588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5289
timestamp 1676037725
transform 1 0 487692 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5301
timestamp 1676037725
transform 1 0 488796 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5313
timestamp 1676037725
transform 1 0 489900 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5319
timestamp 1676037725
transform 1 0 490452 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5321
timestamp 1676037725
transform 1 0 490636 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5333
timestamp 1676037725
transform 1 0 491740 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5345
timestamp 1676037725
transform 1 0 492844 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5357
timestamp 1676037725
transform 1 0 493948 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5369
timestamp 1676037725
transform 1 0 495052 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5375
timestamp 1676037725
transform 1 0 495604 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5377
timestamp 1676037725
transform 1 0 495788 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5389
timestamp 1676037725
transform 1 0 496892 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5401
timestamp 1676037725
transform 1 0 497996 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5413
timestamp 1676037725
transform 1 0 499100 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5425
timestamp 1676037725
transform 1 0 500204 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5431
timestamp 1676037725
transform 1 0 500756 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5433
timestamp 1676037725
transform 1 0 500940 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5445
timestamp 1676037725
transform 1 0 502044 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5457
timestamp 1676037725
transform 1 0 503148 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5469
timestamp 1676037725
transform 1 0 504252 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5481
timestamp 1676037725
transform 1 0 505356 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5487
timestamp 1676037725
transform 1 0 505908 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5489
timestamp 1676037725
transform 1 0 506092 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5501
timestamp 1676037725
transform 1 0 507196 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5513
timestamp 1676037725
transform 1 0 508300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5525
timestamp 1676037725
transform 1 0 509404 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5537
timestamp 1676037725
transform 1 0 510508 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5543
timestamp 1676037725
transform 1 0 511060 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5545
timestamp 1676037725
transform 1 0 511244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5557
timestamp 1676037725
transform 1 0 512348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5569
timestamp 1676037725
transform 1 0 513452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5581
timestamp 1676037725
transform 1 0 514556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5593
timestamp 1676037725
transform 1 0 515660 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5599
timestamp 1676037725
transform 1 0 516212 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5601
timestamp 1676037725
transform 1 0 516396 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5613
timestamp 1676037725
transform 1 0 517500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5625
timestamp 1676037725
transform 1 0 518604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5637
timestamp 1676037725
transform 1 0 519708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5649
timestamp 1676037725
transform 1 0 520812 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5655
timestamp 1676037725
transform 1 0 521364 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5657
timestamp 1676037725
transform 1 0 521548 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5669
timestamp 1676037725
transform 1 0 522652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5681
timestamp 1676037725
transform 1 0 523756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5693
timestamp 1676037725
transform 1 0 524860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5705
timestamp 1676037725
transform 1 0 525964 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5711
timestamp 1676037725
transform 1 0 526516 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5713
timestamp 1676037725
transform 1 0 526700 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_5725
timestamp 1676037725
transform 1 0 527804 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1676037725
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1676037725
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1676037725
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1676037725
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1676037725
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1676037725
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1676037725
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1676037725
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1676037725
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1676037725
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1676037725
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1676037725
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1676037725
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1676037725
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1676037725
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1676037725
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1676037725
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1676037725
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1676037725
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1676037725
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1676037725
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1676037725
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1676037725
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1676037725
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1676037725
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1676037725
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1676037725
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1676037725
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1676037725
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1676037725
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1676037725
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_725
timestamp 1676037725
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_737
timestamp 1676037725
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 1676037725
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1676037725
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1676037725
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1676037725
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_781
timestamp 1676037725
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_793
timestamp 1676037725
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1676037725
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1676037725
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_813
timestamp 1676037725
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_825
timestamp 1676037725
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_837
timestamp 1676037725
transform 1 0 78108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_849
timestamp 1676037725
transform 1 0 79212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_861
timestamp 1676037725
transform 1 0 80316 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_867
timestamp 1676037725
transform 1 0 80868 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_869
timestamp 1676037725
transform 1 0 81052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_881
timestamp 1676037725
transform 1 0 82156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_893
timestamp 1676037725
transform 1 0 83260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_905
timestamp 1676037725
transform 1 0 84364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_917
timestamp 1676037725
transform 1 0 85468 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_923
timestamp 1676037725
transform 1 0 86020 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_925
timestamp 1676037725
transform 1 0 86204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_937
timestamp 1676037725
transform 1 0 87308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_949
timestamp 1676037725
transform 1 0 88412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_961
timestamp 1676037725
transform 1 0 89516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_973
timestamp 1676037725
transform 1 0 90620 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_979
timestamp 1676037725
transform 1 0 91172 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_981
timestamp 1676037725
transform 1 0 91356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_993
timestamp 1676037725
transform 1 0 92460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1005
timestamp 1676037725
transform 1 0 93564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1017
timestamp 1676037725
transform 1 0 94668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1029
timestamp 1676037725
transform 1 0 95772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1035
timestamp 1676037725
transform 1 0 96324 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1037
timestamp 1676037725
transform 1 0 96508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1049
timestamp 1676037725
transform 1 0 97612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1061
timestamp 1676037725
transform 1 0 98716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1073
timestamp 1676037725
transform 1 0 99820 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1085
timestamp 1676037725
transform 1 0 100924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1091
timestamp 1676037725
transform 1 0 101476 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1093
timestamp 1676037725
transform 1 0 101660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1105
timestamp 1676037725
transform 1 0 102764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1117
timestamp 1676037725
transform 1 0 103868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1129
timestamp 1676037725
transform 1 0 104972 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1141
timestamp 1676037725
transform 1 0 106076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1147
timestamp 1676037725
transform 1 0 106628 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1149
timestamp 1676037725
transform 1 0 106812 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1161
timestamp 1676037725
transform 1 0 107916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1173
timestamp 1676037725
transform 1 0 109020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1185
timestamp 1676037725
transform 1 0 110124 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1197
timestamp 1676037725
transform 1 0 111228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1203
timestamp 1676037725
transform 1 0 111780 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1205
timestamp 1676037725
transform 1 0 111964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1217
timestamp 1676037725
transform 1 0 113068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1229
timestamp 1676037725
transform 1 0 114172 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1241
timestamp 1676037725
transform 1 0 115276 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1253
timestamp 1676037725
transform 1 0 116380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1259
timestamp 1676037725
transform 1 0 116932 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1261
timestamp 1676037725
transform 1 0 117116 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1273
timestamp 1676037725
transform 1 0 118220 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1285
timestamp 1676037725
transform 1 0 119324 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1297
timestamp 1676037725
transform 1 0 120428 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1309
timestamp 1676037725
transform 1 0 121532 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1315
timestamp 1676037725
transform 1 0 122084 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1317
timestamp 1676037725
transform 1 0 122268 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1329
timestamp 1676037725
transform 1 0 123372 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1341
timestamp 1676037725
transform 1 0 124476 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1353
timestamp 1676037725
transform 1 0 125580 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1365
timestamp 1676037725
transform 1 0 126684 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1371
timestamp 1676037725
transform 1 0 127236 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1373
timestamp 1676037725
transform 1 0 127420 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1385
timestamp 1676037725
transform 1 0 128524 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1397
timestamp 1676037725
transform 1 0 129628 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1409
timestamp 1676037725
transform 1 0 130732 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1421
timestamp 1676037725
transform 1 0 131836 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1427
timestamp 1676037725
transform 1 0 132388 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1429
timestamp 1676037725
transform 1 0 132572 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1441
timestamp 1676037725
transform 1 0 133676 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1453
timestamp 1676037725
transform 1 0 134780 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1465
timestamp 1676037725
transform 1 0 135884 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1477
timestamp 1676037725
transform 1 0 136988 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1483
timestamp 1676037725
transform 1 0 137540 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1485
timestamp 1676037725
transform 1 0 137724 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1497
timestamp 1676037725
transform 1 0 138828 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1509
timestamp 1676037725
transform 1 0 139932 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1521
timestamp 1676037725
transform 1 0 141036 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1533
timestamp 1676037725
transform 1 0 142140 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1539
timestamp 1676037725
transform 1 0 142692 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1541
timestamp 1676037725
transform 1 0 142876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1553
timestamp 1676037725
transform 1 0 143980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1565
timestamp 1676037725
transform 1 0 145084 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1577
timestamp 1676037725
transform 1 0 146188 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1589
timestamp 1676037725
transform 1 0 147292 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1595
timestamp 1676037725
transform 1 0 147844 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1597
timestamp 1676037725
transform 1 0 148028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1609
timestamp 1676037725
transform 1 0 149132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1621
timestamp 1676037725
transform 1 0 150236 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1633
timestamp 1676037725
transform 1 0 151340 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1645
timestamp 1676037725
transform 1 0 152444 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1651
timestamp 1676037725
transform 1 0 152996 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1653
timestamp 1676037725
transform 1 0 153180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1665
timestamp 1676037725
transform 1 0 154284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1677
timestamp 1676037725
transform 1 0 155388 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1689
timestamp 1676037725
transform 1 0 156492 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1701
timestamp 1676037725
transform 1 0 157596 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1707
timestamp 1676037725
transform 1 0 158148 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1709
timestamp 1676037725
transform 1 0 158332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1721
timestamp 1676037725
transform 1 0 159436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1733
timestamp 1676037725
transform 1 0 160540 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1745
timestamp 1676037725
transform 1 0 161644 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1757
timestamp 1676037725
transform 1 0 162748 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1763
timestamp 1676037725
transform 1 0 163300 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1765
timestamp 1676037725
transform 1 0 163484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1777
timestamp 1676037725
transform 1 0 164588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1789
timestamp 1676037725
transform 1 0 165692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1801
timestamp 1676037725
transform 1 0 166796 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1813
timestamp 1676037725
transform 1 0 167900 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1819
timestamp 1676037725
transform 1 0 168452 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1821
timestamp 1676037725
transform 1 0 168636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1833
timestamp 1676037725
transform 1 0 169740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1845
timestamp 1676037725
transform 1 0 170844 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1857
timestamp 1676037725
transform 1 0 171948 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1869
timestamp 1676037725
transform 1 0 173052 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1875
timestamp 1676037725
transform 1 0 173604 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1877
timestamp 1676037725
transform 1 0 173788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1889
timestamp 1676037725
transform 1 0 174892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1901
timestamp 1676037725
transform 1 0 175996 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1913
timestamp 1676037725
transform 1 0 177100 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1925
timestamp 1676037725
transform 1 0 178204 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1931
timestamp 1676037725
transform 1 0 178756 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1933
timestamp 1676037725
transform 1 0 178940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1945
timestamp 1676037725
transform 1 0 180044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1957
timestamp 1676037725
transform 1 0 181148 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1969
timestamp 1676037725
transform 1 0 182252 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1981
timestamp 1676037725
transform 1 0 183356 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1987
timestamp 1676037725
transform 1 0 183908 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1989
timestamp 1676037725
transform 1 0 184092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2001
timestamp 1676037725
transform 1 0 185196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2013
timestamp 1676037725
transform 1 0 186300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2025
timestamp 1676037725
transform 1 0 187404 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2037
timestamp 1676037725
transform 1 0 188508 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2043
timestamp 1676037725
transform 1 0 189060 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2045
timestamp 1676037725
transform 1 0 189244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2057
timestamp 1676037725
transform 1 0 190348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2069
timestamp 1676037725
transform 1 0 191452 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2081
timestamp 1676037725
transform 1 0 192556 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2093
timestamp 1676037725
transform 1 0 193660 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2099
timestamp 1676037725
transform 1 0 194212 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2101
timestamp 1676037725
transform 1 0 194396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2113
timestamp 1676037725
transform 1 0 195500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2125
timestamp 1676037725
transform 1 0 196604 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2137
timestamp 1676037725
transform 1 0 197708 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2149
timestamp 1676037725
transform 1 0 198812 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2155
timestamp 1676037725
transform 1 0 199364 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2157
timestamp 1676037725
transform 1 0 199548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2169
timestamp 1676037725
transform 1 0 200652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2181
timestamp 1676037725
transform 1 0 201756 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2193
timestamp 1676037725
transform 1 0 202860 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2205
timestamp 1676037725
transform 1 0 203964 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2211
timestamp 1676037725
transform 1 0 204516 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2213
timestamp 1676037725
transform 1 0 204700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2225
timestamp 1676037725
transform 1 0 205804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2237
timestamp 1676037725
transform 1 0 206908 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2249
timestamp 1676037725
transform 1 0 208012 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2261
timestamp 1676037725
transform 1 0 209116 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2267
timestamp 1676037725
transform 1 0 209668 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2269
timestamp 1676037725
transform 1 0 209852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2281
timestamp 1676037725
transform 1 0 210956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2293
timestamp 1676037725
transform 1 0 212060 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2305
timestamp 1676037725
transform 1 0 213164 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2317
timestamp 1676037725
transform 1 0 214268 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2323
timestamp 1676037725
transform 1 0 214820 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2325
timestamp 1676037725
transform 1 0 215004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2337
timestamp 1676037725
transform 1 0 216108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2349
timestamp 1676037725
transform 1 0 217212 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2361
timestamp 1676037725
transform 1 0 218316 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2373
timestamp 1676037725
transform 1 0 219420 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2379
timestamp 1676037725
transform 1 0 219972 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2381
timestamp 1676037725
transform 1 0 220156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2393
timestamp 1676037725
transform 1 0 221260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2405
timestamp 1676037725
transform 1 0 222364 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2417
timestamp 1676037725
transform 1 0 223468 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2429
timestamp 1676037725
transform 1 0 224572 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2435
timestamp 1676037725
transform 1 0 225124 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2437
timestamp 1676037725
transform 1 0 225308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2449
timestamp 1676037725
transform 1 0 226412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2461
timestamp 1676037725
transform 1 0 227516 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2473
timestamp 1676037725
transform 1 0 228620 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2485
timestamp 1676037725
transform 1 0 229724 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2491
timestamp 1676037725
transform 1 0 230276 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2493
timestamp 1676037725
transform 1 0 230460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2505
timestamp 1676037725
transform 1 0 231564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2517
timestamp 1676037725
transform 1 0 232668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2529
timestamp 1676037725
transform 1 0 233772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2541
timestamp 1676037725
transform 1 0 234876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2547
timestamp 1676037725
transform 1 0 235428 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2549
timestamp 1676037725
transform 1 0 235612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2561
timestamp 1676037725
transform 1 0 236716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2573
timestamp 1676037725
transform 1 0 237820 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2585
timestamp 1676037725
transform 1 0 238924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2597
timestamp 1676037725
transform 1 0 240028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2603
timestamp 1676037725
transform 1 0 240580 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2605
timestamp 1676037725
transform 1 0 240764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2617
timestamp 1676037725
transform 1 0 241868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2629
timestamp 1676037725
transform 1 0 242972 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2641
timestamp 1676037725
transform 1 0 244076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2653
timestamp 1676037725
transform 1 0 245180 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2659
timestamp 1676037725
transform 1 0 245732 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2661
timestamp 1676037725
transform 1 0 245916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2673
timestamp 1676037725
transform 1 0 247020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2685
timestamp 1676037725
transform 1 0 248124 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2697
timestamp 1676037725
transform 1 0 249228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2709
timestamp 1676037725
transform 1 0 250332 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2715
timestamp 1676037725
transform 1 0 250884 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2717
timestamp 1676037725
transform 1 0 251068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2729
timestamp 1676037725
transform 1 0 252172 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2741
timestamp 1676037725
transform 1 0 253276 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2753
timestamp 1676037725
transform 1 0 254380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2765
timestamp 1676037725
transform 1 0 255484 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2771
timestamp 1676037725
transform 1 0 256036 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2773
timestamp 1676037725
transform 1 0 256220 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2785
timestamp 1676037725
transform 1 0 257324 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2797
timestamp 1676037725
transform 1 0 258428 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2809
timestamp 1676037725
transform 1 0 259532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2821
timestamp 1676037725
transform 1 0 260636 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2827
timestamp 1676037725
transform 1 0 261188 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2829
timestamp 1676037725
transform 1 0 261372 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2841
timestamp 1676037725
transform 1 0 262476 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2853
timestamp 1676037725
transform 1 0 263580 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2865
timestamp 1676037725
transform 1 0 264684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2877
timestamp 1676037725
transform 1 0 265788 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2883
timestamp 1676037725
transform 1 0 266340 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2885
timestamp 1676037725
transform 1 0 266524 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2897
timestamp 1676037725
transform 1 0 267628 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2909
timestamp 1676037725
transform 1 0 268732 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2921
timestamp 1676037725
transform 1 0 269836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2933
timestamp 1676037725
transform 1 0 270940 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2939
timestamp 1676037725
transform 1 0 271492 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2941
timestamp 1676037725
transform 1 0 271676 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2953
timestamp 1676037725
transform 1 0 272780 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2965
timestamp 1676037725
transform 1 0 273884 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2977
timestamp 1676037725
transform 1 0 274988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2989
timestamp 1676037725
transform 1 0 276092 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2995
timestamp 1676037725
transform 1 0 276644 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2997
timestamp 1676037725
transform 1 0 276828 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3009
timestamp 1676037725
transform 1 0 277932 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3021
timestamp 1676037725
transform 1 0 279036 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3033
timestamp 1676037725
transform 1 0 280140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3045
timestamp 1676037725
transform 1 0 281244 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3051
timestamp 1676037725
transform 1 0 281796 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3053
timestamp 1676037725
transform 1 0 281980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3065
timestamp 1676037725
transform 1 0 283084 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3077
timestamp 1676037725
transform 1 0 284188 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3089
timestamp 1676037725
transform 1 0 285292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3101
timestamp 1676037725
transform 1 0 286396 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3107
timestamp 1676037725
transform 1 0 286948 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3109
timestamp 1676037725
transform 1 0 287132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3121
timestamp 1676037725
transform 1 0 288236 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3133
timestamp 1676037725
transform 1 0 289340 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3145
timestamp 1676037725
transform 1 0 290444 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3157
timestamp 1676037725
transform 1 0 291548 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3163
timestamp 1676037725
transform 1 0 292100 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3165
timestamp 1676037725
transform 1 0 292284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3177
timestamp 1676037725
transform 1 0 293388 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3189
timestamp 1676037725
transform 1 0 294492 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3201
timestamp 1676037725
transform 1 0 295596 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3213
timestamp 1676037725
transform 1 0 296700 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3219
timestamp 1676037725
transform 1 0 297252 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3221
timestamp 1676037725
transform 1 0 297436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3233
timestamp 1676037725
transform 1 0 298540 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3245
timestamp 1676037725
transform 1 0 299644 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3257
timestamp 1676037725
transform 1 0 300748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3269
timestamp 1676037725
transform 1 0 301852 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3275
timestamp 1676037725
transform 1 0 302404 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3277
timestamp 1676037725
transform 1 0 302588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3289
timestamp 1676037725
transform 1 0 303692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3301
timestamp 1676037725
transform 1 0 304796 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3313
timestamp 1676037725
transform 1 0 305900 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3325
timestamp 1676037725
transform 1 0 307004 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3331
timestamp 1676037725
transform 1 0 307556 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3333
timestamp 1676037725
transform 1 0 307740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3345
timestamp 1676037725
transform 1 0 308844 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3357
timestamp 1676037725
transform 1 0 309948 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3369
timestamp 1676037725
transform 1 0 311052 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3381
timestamp 1676037725
transform 1 0 312156 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3387
timestamp 1676037725
transform 1 0 312708 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3389
timestamp 1676037725
transform 1 0 312892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3401
timestamp 1676037725
transform 1 0 313996 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3413
timestamp 1676037725
transform 1 0 315100 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3425
timestamp 1676037725
transform 1 0 316204 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3437
timestamp 1676037725
transform 1 0 317308 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3443
timestamp 1676037725
transform 1 0 317860 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3445
timestamp 1676037725
transform 1 0 318044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3457
timestamp 1676037725
transform 1 0 319148 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3469
timestamp 1676037725
transform 1 0 320252 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3481
timestamp 1676037725
transform 1 0 321356 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3493
timestamp 1676037725
transform 1 0 322460 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3499
timestamp 1676037725
transform 1 0 323012 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3501
timestamp 1676037725
transform 1 0 323196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3513
timestamp 1676037725
transform 1 0 324300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3525
timestamp 1676037725
transform 1 0 325404 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3537
timestamp 1676037725
transform 1 0 326508 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3549
timestamp 1676037725
transform 1 0 327612 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3555
timestamp 1676037725
transform 1 0 328164 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3557
timestamp 1676037725
transform 1 0 328348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3569
timestamp 1676037725
transform 1 0 329452 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3581
timestamp 1676037725
transform 1 0 330556 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3593
timestamp 1676037725
transform 1 0 331660 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3605
timestamp 1676037725
transform 1 0 332764 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3611
timestamp 1676037725
transform 1 0 333316 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3613
timestamp 1676037725
transform 1 0 333500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3625
timestamp 1676037725
transform 1 0 334604 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3637
timestamp 1676037725
transform 1 0 335708 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3649
timestamp 1676037725
transform 1 0 336812 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3661
timestamp 1676037725
transform 1 0 337916 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3667
timestamp 1676037725
transform 1 0 338468 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3669
timestamp 1676037725
transform 1 0 338652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3681
timestamp 1676037725
transform 1 0 339756 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3693
timestamp 1676037725
transform 1 0 340860 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3705
timestamp 1676037725
transform 1 0 341964 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3717
timestamp 1676037725
transform 1 0 343068 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3723
timestamp 1676037725
transform 1 0 343620 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3725
timestamp 1676037725
transform 1 0 343804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3737
timestamp 1676037725
transform 1 0 344908 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3749
timestamp 1676037725
transform 1 0 346012 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3761
timestamp 1676037725
transform 1 0 347116 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3773
timestamp 1676037725
transform 1 0 348220 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3779
timestamp 1676037725
transform 1 0 348772 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3781
timestamp 1676037725
transform 1 0 348956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3793
timestamp 1676037725
transform 1 0 350060 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3805
timestamp 1676037725
transform 1 0 351164 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3817
timestamp 1676037725
transform 1 0 352268 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3829
timestamp 1676037725
transform 1 0 353372 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3835
timestamp 1676037725
transform 1 0 353924 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3837
timestamp 1676037725
transform 1 0 354108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3849
timestamp 1676037725
transform 1 0 355212 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3861
timestamp 1676037725
transform 1 0 356316 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3873
timestamp 1676037725
transform 1 0 357420 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3885
timestamp 1676037725
transform 1 0 358524 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3891
timestamp 1676037725
transform 1 0 359076 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3893
timestamp 1676037725
transform 1 0 359260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3905
timestamp 1676037725
transform 1 0 360364 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3917
timestamp 1676037725
transform 1 0 361468 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3929
timestamp 1676037725
transform 1 0 362572 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3941
timestamp 1676037725
transform 1 0 363676 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3947
timestamp 1676037725
transform 1 0 364228 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3949
timestamp 1676037725
transform 1 0 364412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3961
timestamp 1676037725
transform 1 0 365516 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3973
timestamp 1676037725
transform 1 0 366620 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3985
timestamp 1676037725
transform 1 0 367724 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3997
timestamp 1676037725
transform 1 0 368828 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4003
timestamp 1676037725
transform 1 0 369380 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4005
timestamp 1676037725
transform 1 0 369564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4017
timestamp 1676037725
transform 1 0 370668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4029
timestamp 1676037725
transform 1 0 371772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4041
timestamp 1676037725
transform 1 0 372876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4053
timestamp 1676037725
transform 1 0 373980 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4059
timestamp 1676037725
transform 1 0 374532 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4061
timestamp 1676037725
transform 1 0 374716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4073
timestamp 1676037725
transform 1 0 375820 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4085
timestamp 1676037725
transform 1 0 376924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4097
timestamp 1676037725
transform 1 0 378028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4109
timestamp 1676037725
transform 1 0 379132 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4115
timestamp 1676037725
transform 1 0 379684 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4117
timestamp 1676037725
transform 1 0 379868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4129
timestamp 1676037725
transform 1 0 380972 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4141
timestamp 1676037725
transform 1 0 382076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4153
timestamp 1676037725
transform 1 0 383180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4165
timestamp 1676037725
transform 1 0 384284 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4171
timestamp 1676037725
transform 1 0 384836 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4173
timestamp 1676037725
transform 1 0 385020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4185
timestamp 1676037725
transform 1 0 386124 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4197
timestamp 1676037725
transform 1 0 387228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4209
timestamp 1676037725
transform 1 0 388332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4221
timestamp 1676037725
transform 1 0 389436 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4227
timestamp 1676037725
transform 1 0 389988 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4229
timestamp 1676037725
transform 1 0 390172 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4241
timestamp 1676037725
transform 1 0 391276 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4253
timestamp 1676037725
transform 1 0 392380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4265
timestamp 1676037725
transform 1 0 393484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4277
timestamp 1676037725
transform 1 0 394588 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4283
timestamp 1676037725
transform 1 0 395140 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4285
timestamp 1676037725
transform 1 0 395324 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4297
timestamp 1676037725
transform 1 0 396428 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4309
timestamp 1676037725
transform 1 0 397532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4321
timestamp 1676037725
transform 1 0 398636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4333
timestamp 1676037725
transform 1 0 399740 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4339
timestamp 1676037725
transform 1 0 400292 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4341
timestamp 1676037725
transform 1 0 400476 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4353
timestamp 1676037725
transform 1 0 401580 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4365
timestamp 1676037725
transform 1 0 402684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4377
timestamp 1676037725
transform 1 0 403788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4389
timestamp 1676037725
transform 1 0 404892 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4395
timestamp 1676037725
transform 1 0 405444 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4397
timestamp 1676037725
transform 1 0 405628 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4409
timestamp 1676037725
transform 1 0 406732 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4421
timestamp 1676037725
transform 1 0 407836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4433
timestamp 1676037725
transform 1 0 408940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4445
timestamp 1676037725
transform 1 0 410044 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4451
timestamp 1676037725
transform 1 0 410596 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4453
timestamp 1676037725
transform 1 0 410780 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4465
timestamp 1676037725
transform 1 0 411884 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4477
timestamp 1676037725
transform 1 0 412988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4489
timestamp 1676037725
transform 1 0 414092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4501
timestamp 1676037725
transform 1 0 415196 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4507
timestamp 1676037725
transform 1 0 415748 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4509
timestamp 1676037725
transform 1 0 415932 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4521
timestamp 1676037725
transform 1 0 417036 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4533
timestamp 1676037725
transform 1 0 418140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4545
timestamp 1676037725
transform 1 0 419244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4557
timestamp 1676037725
transform 1 0 420348 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4563
timestamp 1676037725
transform 1 0 420900 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4565
timestamp 1676037725
transform 1 0 421084 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4577
timestamp 1676037725
transform 1 0 422188 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4589
timestamp 1676037725
transform 1 0 423292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4601
timestamp 1676037725
transform 1 0 424396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4613
timestamp 1676037725
transform 1 0 425500 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4619
timestamp 1676037725
transform 1 0 426052 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4621
timestamp 1676037725
transform 1 0 426236 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4633
timestamp 1676037725
transform 1 0 427340 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4645
timestamp 1676037725
transform 1 0 428444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4657
timestamp 1676037725
transform 1 0 429548 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4669
timestamp 1676037725
transform 1 0 430652 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4675
timestamp 1676037725
transform 1 0 431204 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4677
timestamp 1676037725
transform 1 0 431388 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4689
timestamp 1676037725
transform 1 0 432492 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4701
timestamp 1676037725
transform 1 0 433596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4713
timestamp 1676037725
transform 1 0 434700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4725
timestamp 1676037725
transform 1 0 435804 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4731
timestamp 1676037725
transform 1 0 436356 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4733
timestamp 1676037725
transform 1 0 436540 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4745
timestamp 1676037725
transform 1 0 437644 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4757
timestamp 1676037725
transform 1 0 438748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4769
timestamp 1676037725
transform 1 0 439852 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4781
timestamp 1676037725
transform 1 0 440956 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4787
timestamp 1676037725
transform 1 0 441508 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4789
timestamp 1676037725
transform 1 0 441692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4801
timestamp 1676037725
transform 1 0 442796 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4813
timestamp 1676037725
transform 1 0 443900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4825
timestamp 1676037725
transform 1 0 445004 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4837
timestamp 1676037725
transform 1 0 446108 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4843
timestamp 1676037725
transform 1 0 446660 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4845
timestamp 1676037725
transform 1 0 446844 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4857
timestamp 1676037725
transform 1 0 447948 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4869
timestamp 1676037725
transform 1 0 449052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4881
timestamp 1676037725
transform 1 0 450156 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4893
timestamp 1676037725
transform 1 0 451260 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4899
timestamp 1676037725
transform 1 0 451812 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4901
timestamp 1676037725
transform 1 0 451996 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4913
timestamp 1676037725
transform 1 0 453100 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4925
timestamp 1676037725
transform 1 0 454204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4937
timestamp 1676037725
transform 1 0 455308 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4949
timestamp 1676037725
transform 1 0 456412 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4955
timestamp 1676037725
transform 1 0 456964 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4957
timestamp 1676037725
transform 1 0 457148 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4969
timestamp 1676037725
transform 1 0 458252 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4981
timestamp 1676037725
transform 1 0 459356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4993
timestamp 1676037725
transform 1 0 460460 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5005
timestamp 1676037725
transform 1 0 461564 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5011
timestamp 1676037725
transform 1 0 462116 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5013
timestamp 1676037725
transform 1 0 462300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5025
timestamp 1676037725
transform 1 0 463404 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5037
timestamp 1676037725
transform 1 0 464508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5049
timestamp 1676037725
transform 1 0 465612 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5061
timestamp 1676037725
transform 1 0 466716 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5067
timestamp 1676037725
transform 1 0 467268 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5069
timestamp 1676037725
transform 1 0 467452 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5081
timestamp 1676037725
transform 1 0 468556 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5093
timestamp 1676037725
transform 1 0 469660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5105
timestamp 1676037725
transform 1 0 470764 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5117
timestamp 1676037725
transform 1 0 471868 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5123
timestamp 1676037725
transform 1 0 472420 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5125
timestamp 1676037725
transform 1 0 472604 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5137
timestamp 1676037725
transform 1 0 473708 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5149
timestamp 1676037725
transform 1 0 474812 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5161
timestamp 1676037725
transform 1 0 475916 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5173
timestamp 1676037725
transform 1 0 477020 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5179
timestamp 1676037725
transform 1 0 477572 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5181
timestamp 1676037725
transform 1 0 477756 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5193
timestamp 1676037725
transform 1 0 478860 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5205
timestamp 1676037725
transform 1 0 479964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5217
timestamp 1676037725
transform 1 0 481068 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5229
timestamp 1676037725
transform 1 0 482172 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5235
timestamp 1676037725
transform 1 0 482724 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5237
timestamp 1676037725
transform 1 0 482908 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5249
timestamp 1676037725
transform 1 0 484012 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5261
timestamp 1676037725
transform 1 0 485116 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5273
timestamp 1676037725
transform 1 0 486220 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5285
timestamp 1676037725
transform 1 0 487324 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5291
timestamp 1676037725
transform 1 0 487876 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5293
timestamp 1676037725
transform 1 0 488060 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5305
timestamp 1676037725
transform 1 0 489164 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5317
timestamp 1676037725
transform 1 0 490268 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5329
timestamp 1676037725
transform 1 0 491372 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5341
timestamp 1676037725
transform 1 0 492476 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5347
timestamp 1676037725
transform 1 0 493028 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5349
timestamp 1676037725
transform 1 0 493212 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5361
timestamp 1676037725
transform 1 0 494316 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5373
timestamp 1676037725
transform 1 0 495420 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5385
timestamp 1676037725
transform 1 0 496524 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5397
timestamp 1676037725
transform 1 0 497628 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5403
timestamp 1676037725
transform 1 0 498180 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5405
timestamp 1676037725
transform 1 0 498364 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5417
timestamp 1676037725
transform 1 0 499468 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5429
timestamp 1676037725
transform 1 0 500572 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5441
timestamp 1676037725
transform 1 0 501676 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5453
timestamp 1676037725
transform 1 0 502780 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5459
timestamp 1676037725
transform 1 0 503332 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5461
timestamp 1676037725
transform 1 0 503516 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5473
timestamp 1676037725
transform 1 0 504620 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5485
timestamp 1676037725
transform 1 0 505724 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5497
timestamp 1676037725
transform 1 0 506828 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5509
timestamp 1676037725
transform 1 0 507932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5515
timestamp 1676037725
transform 1 0 508484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5517
timestamp 1676037725
transform 1 0 508668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5529
timestamp 1676037725
transform 1 0 509772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5541
timestamp 1676037725
transform 1 0 510876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5553
timestamp 1676037725
transform 1 0 511980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5565
timestamp 1676037725
transform 1 0 513084 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5571
timestamp 1676037725
transform 1 0 513636 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5573
timestamp 1676037725
transform 1 0 513820 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5585
timestamp 1676037725
transform 1 0 514924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5597
timestamp 1676037725
transform 1 0 516028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5609
timestamp 1676037725
transform 1 0 517132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5621
timestamp 1676037725
transform 1 0 518236 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5627
timestamp 1676037725
transform 1 0 518788 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5629
timestamp 1676037725
transform 1 0 518972 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5641
timestamp 1676037725
transform 1 0 520076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5653
timestamp 1676037725
transform 1 0 521180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5665
timestamp 1676037725
transform 1 0 522284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5677
timestamp 1676037725
transform 1 0 523388 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5683
timestamp 1676037725
transform 1 0 523940 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5685
timestamp 1676037725
transform 1 0 524124 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5697
timestamp 1676037725
transform 1 0 525228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5709
timestamp 1676037725
transform 1 0 526332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5721
timestamp 1676037725
transform 1 0 527436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1676037725
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1676037725
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1676037725
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1676037725
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1676037725
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1676037725
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1676037725
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1676037725
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1676037725
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1676037725
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1676037725
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1676037725
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1676037725
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1676037725
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1676037725
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1676037725
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1676037725
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1676037725
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1676037725
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1676037725
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1676037725
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1676037725
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1676037725
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1676037725
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1676037725
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1676037725
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1676037725
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1676037725
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1676037725
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1676037725
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_729
timestamp 1676037725
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_741
timestamp 1676037725
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_753
timestamp 1676037725
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_765
timestamp 1676037725
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1676037725
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1676037725
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_785
timestamp 1676037725
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_797
timestamp 1676037725
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_809
timestamp 1676037725
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_821
timestamp 1676037725
transform 1 0 76636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_833
timestamp 1676037725
transform 1 0 77740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_839
timestamp 1676037725
transform 1 0 78292 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_841
timestamp 1676037725
transform 1 0 78476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_853
timestamp 1676037725
transform 1 0 79580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_865
timestamp 1676037725
transform 1 0 80684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_877
timestamp 1676037725
transform 1 0 81788 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_889
timestamp 1676037725
transform 1 0 82892 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_895
timestamp 1676037725
transform 1 0 83444 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_897
timestamp 1676037725
transform 1 0 83628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_909
timestamp 1676037725
transform 1 0 84732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_921
timestamp 1676037725
transform 1 0 85836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_933
timestamp 1676037725
transform 1 0 86940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_945
timestamp 1676037725
transform 1 0 88044 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_951
timestamp 1676037725
transform 1 0 88596 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_953
timestamp 1676037725
transform 1 0 88780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_965
timestamp 1676037725
transform 1 0 89884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_977
timestamp 1676037725
transform 1 0 90988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_989
timestamp 1676037725
transform 1 0 92092 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1001
timestamp 1676037725
transform 1 0 93196 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1007
timestamp 1676037725
transform 1 0 93748 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1009
timestamp 1676037725
transform 1 0 93932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1021
timestamp 1676037725
transform 1 0 95036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1033
timestamp 1676037725
transform 1 0 96140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1045
timestamp 1676037725
transform 1 0 97244 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1057
timestamp 1676037725
transform 1 0 98348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1063
timestamp 1676037725
transform 1 0 98900 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1065
timestamp 1676037725
transform 1 0 99084 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1077
timestamp 1676037725
transform 1 0 100188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1089
timestamp 1676037725
transform 1 0 101292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1101
timestamp 1676037725
transform 1 0 102396 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1113
timestamp 1676037725
transform 1 0 103500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1119
timestamp 1676037725
transform 1 0 104052 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1121
timestamp 1676037725
transform 1 0 104236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1133
timestamp 1676037725
transform 1 0 105340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1145
timestamp 1676037725
transform 1 0 106444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1157
timestamp 1676037725
transform 1 0 107548 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1169
timestamp 1676037725
transform 1 0 108652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1175
timestamp 1676037725
transform 1 0 109204 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1177
timestamp 1676037725
transform 1 0 109388 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1189
timestamp 1676037725
transform 1 0 110492 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1201
timestamp 1676037725
transform 1 0 111596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1213
timestamp 1676037725
transform 1 0 112700 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1225
timestamp 1676037725
transform 1 0 113804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1231
timestamp 1676037725
transform 1 0 114356 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1233
timestamp 1676037725
transform 1 0 114540 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1245
timestamp 1676037725
transform 1 0 115644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1257
timestamp 1676037725
transform 1 0 116748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1269
timestamp 1676037725
transform 1 0 117852 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1281
timestamp 1676037725
transform 1 0 118956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1287
timestamp 1676037725
transform 1 0 119508 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1289
timestamp 1676037725
transform 1 0 119692 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1301
timestamp 1676037725
transform 1 0 120796 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1313
timestamp 1676037725
transform 1 0 121900 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1325
timestamp 1676037725
transform 1 0 123004 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1337
timestamp 1676037725
transform 1 0 124108 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1343
timestamp 1676037725
transform 1 0 124660 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1345
timestamp 1676037725
transform 1 0 124844 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1357
timestamp 1676037725
transform 1 0 125948 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1369
timestamp 1676037725
transform 1 0 127052 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1381
timestamp 1676037725
transform 1 0 128156 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1393
timestamp 1676037725
transform 1 0 129260 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1399
timestamp 1676037725
transform 1 0 129812 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1401
timestamp 1676037725
transform 1 0 129996 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1413
timestamp 1676037725
transform 1 0 131100 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1425
timestamp 1676037725
transform 1 0 132204 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1437
timestamp 1676037725
transform 1 0 133308 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1449
timestamp 1676037725
transform 1 0 134412 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1455
timestamp 1676037725
transform 1 0 134964 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1457
timestamp 1676037725
transform 1 0 135148 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1469
timestamp 1676037725
transform 1 0 136252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1481
timestamp 1676037725
transform 1 0 137356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1493
timestamp 1676037725
transform 1 0 138460 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1505
timestamp 1676037725
transform 1 0 139564 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1511
timestamp 1676037725
transform 1 0 140116 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1513
timestamp 1676037725
transform 1 0 140300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1525
timestamp 1676037725
transform 1 0 141404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1537
timestamp 1676037725
transform 1 0 142508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1549
timestamp 1676037725
transform 1 0 143612 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1561
timestamp 1676037725
transform 1 0 144716 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1567
timestamp 1676037725
transform 1 0 145268 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1569
timestamp 1676037725
transform 1 0 145452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1581
timestamp 1676037725
transform 1 0 146556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1593
timestamp 1676037725
transform 1 0 147660 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1605
timestamp 1676037725
transform 1 0 148764 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1617
timestamp 1676037725
transform 1 0 149868 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1623
timestamp 1676037725
transform 1 0 150420 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1625
timestamp 1676037725
transform 1 0 150604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1637
timestamp 1676037725
transform 1 0 151708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1649
timestamp 1676037725
transform 1 0 152812 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1661
timestamp 1676037725
transform 1 0 153916 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1673
timestamp 1676037725
transform 1 0 155020 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1679
timestamp 1676037725
transform 1 0 155572 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1681
timestamp 1676037725
transform 1 0 155756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1693
timestamp 1676037725
transform 1 0 156860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1705
timestamp 1676037725
transform 1 0 157964 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1717
timestamp 1676037725
transform 1 0 159068 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1729
timestamp 1676037725
transform 1 0 160172 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1735
timestamp 1676037725
transform 1 0 160724 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1737
timestamp 1676037725
transform 1 0 160908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1749
timestamp 1676037725
transform 1 0 162012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1761
timestamp 1676037725
transform 1 0 163116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1773
timestamp 1676037725
transform 1 0 164220 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1785
timestamp 1676037725
transform 1 0 165324 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1791
timestamp 1676037725
transform 1 0 165876 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1793
timestamp 1676037725
transform 1 0 166060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1805
timestamp 1676037725
transform 1 0 167164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1817
timestamp 1676037725
transform 1 0 168268 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1829
timestamp 1676037725
transform 1 0 169372 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1841
timestamp 1676037725
transform 1 0 170476 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1847
timestamp 1676037725
transform 1 0 171028 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1849
timestamp 1676037725
transform 1 0 171212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1861
timestamp 1676037725
transform 1 0 172316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1873
timestamp 1676037725
transform 1 0 173420 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1885
timestamp 1676037725
transform 1 0 174524 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1897
timestamp 1676037725
transform 1 0 175628 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1903
timestamp 1676037725
transform 1 0 176180 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1905
timestamp 1676037725
transform 1 0 176364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1917
timestamp 1676037725
transform 1 0 177468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1929
timestamp 1676037725
transform 1 0 178572 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1941
timestamp 1676037725
transform 1 0 179676 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1953
timestamp 1676037725
transform 1 0 180780 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1959
timestamp 1676037725
transform 1 0 181332 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1961
timestamp 1676037725
transform 1 0 181516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1973
timestamp 1676037725
transform 1 0 182620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1985
timestamp 1676037725
transform 1 0 183724 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1997
timestamp 1676037725
transform 1 0 184828 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2009
timestamp 1676037725
transform 1 0 185932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2015
timestamp 1676037725
transform 1 0 186484 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2017
timestamp 1676037725
transform 1 0 186668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2029
timestamp 1676037725
transform 1 0 187772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2041
timestamp 1676037725
transform 1 0 188876 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2053
timestamp 1676037725
transform 1 0 189980 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2065
timestamp 1676037725
transform 1 0 191084 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2071
timestamp 1676037725
transform 1 0 191636 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2073
timestamp 1676037725
transform 1 0 191820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2085
timestamp 1676037725
transform 1 0 192924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2097
timestamp 1676037725
transform 1 0 194028 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2109
timestamp 1676037725
transform 1 0 195132 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2121
timestamp 1676037725
transform 1 0 196236 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2127
timestamp 1676037725
transform 1 0 196788 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2129
timestamp 1676037725
transform 1 0 196972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2141
timestamp 1676037725
transform 1 0 198076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2153
timestamp 1676037725
transform 1 0 199180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2165
timestamp 1676037725
transform 1 0 200284 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2177
timestamp 1676037725
transform 1 0 201388 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2183
timestamp 1676037725
transform 1 0 201940 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2185
timestamp 1676037725
transform 1 0 202124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2197
timestamp 1676037725
transform 1 0 203228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2209
timestamp 1676037725
transform 1 0 204332 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2221
timestamp 1676037725
transform 1 0 205436 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2233
timestamp 1676037725
transform 1 0 206540 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2239
timestamp 1676037725
transform 1 0 207092 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2241
timestamp 1676037725
transform 1 0 207276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2253
timestamp 1676037725
transform 1 0 208380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2265
timestamp 1676037725
transform 1 0 209484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2277
timestamp 1676037725
transform 1 0 210588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2289
timestamp 1676037725
transform 1 0 211692 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2295
timestamp 1676037725
transform 1 0 212244 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2297
timestamp 1676037725
transform 1 0 212428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2309
timestamp 1676037725
transform 1 0 213532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2321
timestamp 1676037725
transform 1 0 214636 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2333
timestamp 1676037725
transform 1 0 215740 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2345
timestamp 1676037725
transform 1 0 216844 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2351
timestamp 1676037725
transform 1 0 217396 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2353
timestamp 1676037725
transform 1 0 217580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2365
timestamp 1676037725
transform 1 0 218684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2377
timestamp 1676037725
transform 1 0 219788 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2389
timestamp 1676037725
transform 1 0 220892 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2401
timestamp 1676037725
transform 1 0 221996 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2407
timestamp 1676037725
transform 1 0 222548 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2409
timestamp 1676037725
transform 1 0 222732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2421
timestamp 1676037725
transform 1 0 223836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2433
timestamp 1676037725
transform 1 0 224940 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2445
timestamp 1676037725
transform 1 0 226044 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2457
timestamp 1676037725
transform 1 0 227148 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2463
timestamp 1676037725
transform 1 0 227700 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2465
timestamp 1676037725
transform 1 0 227884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2477
timestamp 1676037725
transform 1 0 228988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2489
timestamp 1676037725
transform 1 0 230092 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2501
timestamp 1676037725
transform 1 0 231196 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2513
timestamp 1676037725
transform 1 0 232300 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2519
timestamp 1676037725
transform 1 0 232852 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2521
timestamp 1676037725
transform 1 0 233036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2533
timestamp 1676037725
transform 1 0 234140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2545
timestamp 1676037725
transform 1 0 235244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2557
timestamp 1676037725
transform 1 0 236348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2569
timestamp 1676037725
transform 1 0 237452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2575
timestamp 1676037725
transform 1 0 238004 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2577
timestamp 1676037725
transform 1 0 238188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2589
timestamp 1676037725
transform 1 0 239292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2601
timestamp 1676037725
transform 1 0 240396 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2613
timestamp 1676037725
transform 1 0 241500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2625
timestamp 1676037725
transform 1 0 242604 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2631
timestamp 1676037725
transform 1 0 243156 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2633
timestamp 1676037725
transform 1 0 243340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2645
timestamp 1676037725
transform 1 0 244444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2657
timestamp 1676037725
transform 1 0 245548 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2669
timestamp 1676037725
transform 1 0 246652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2681
timestamp 1676037725
transform 1 0 247756 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2687
timestamp 1676037725
transform 1 0 248308 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2689
timestamp 1676037725
transform 1 0 248492 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2701
timestamp 1676037725
transform 1 0 249596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2713
timestamp 1676037725
transform 1 0 250700 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2725
timestamp 1676037725
transform 1 0 251804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2737
timestamp 1676037725
transform 1 0 252908 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2743
timestamp 1676037725
transform 1 0 253460 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2745
timestamp 1676037725
transform 1 0 253644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2757
timestamp 1676037725
transform 1 0 254748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2769
timestamp 1676037725
transform 1 0 255852 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2781
timestamp 1676037725
transform 1 0 256956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2793
timestamp 1676037725
transform 1 0 258060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2799
timestamp 1676037725
transform 1 0 258612 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2801
timestamp 1676037725
transform 1 0 258796 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2813
timestamp 1676037725
transform 1 0 259900 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2825
timestamp 1676037725
transform 1 0 261004 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2837
timestamp 1676037725
transform 1 0 262108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2849
timestamp 1676037725
transform 1 0 263212 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2855
timestamp 1676037725
transform 1 0 263764 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2857
timestamp 1676037725
transform 1 0 263948 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2869
timestamp 1676037725
transform 1 0 265052 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2881
timestamp 1676037725
transform 1 0 266156 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2893
timestamp 1676037725
transform 1 0 267260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2905
timestamp 1676037725
transform 1 0 268364 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2911
timestamp 1676037725
transform 1 0 268916 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2913
timestamp 1676037725
transform 1 0 269100 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2925
timestamp 1676037725
transform 1 0 270204 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2937
timestamp 1676037725
transform 1 0 271308 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2949
timestamp 1676037725
transform 1 0 272412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2961
timestamp 1676037725
transform 1 0 273516 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2967
timestamp 1676037725
transform 1 0 274068 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2969
timestamp 1676037725
transform 1 0 274252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2981
timestamp 1676037725
transform 1 0 275356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2993
timestamp 1676037725
transform 1 0 276460 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3005
timestamp 1676037725
transform 1 0 277564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3017
timestamp 1676037725
transform 1 0 278668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3023
timestamp 1676037725
transform 1 0 279220 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3025
timestamp 1676037725
transform 1 0 279404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3037
timestamp 1676037725
transform 1 0 280508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3049
timestamp 1676037725
transform 1 0 281612 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3061
timestamp 1676037725
transform 1 0 282716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3073
timestamp 1676037725
transform 1 0 283820 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3079
timestamp 1676037725
transform 1 0 284372 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3081
timestamp 1676037725
transform 1 0 284556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3093
timestamp 1676037725
transform 1 0 285660 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3105
timestamp 1676037725
transform 1 0 286764 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3117
timestamp 1676037725
transform 1 0 287868 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3129
timestamp 1676037725
transform 1 0 288972 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3135
timestamp 1676037725
transform 1 0 289524 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3137
timestamp 1676037725
transform 1 0 289708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3149
timestamp 1676037725
transform 1 0 290812 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3161
timestamp 1676037725
transform 1 0 291916 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3173
timestamp 1676037725
transform 1 0 293020 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3185
timestamp 1676037725
transform 1 0 294124 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3191
timestamp 1676037725
transform 1 0 294676 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3193
timestamp 1676037725
transform 1 0 294860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3205
timestamp 1676037725
transform 1 0 295964 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3217
timestamp 1676037725
transform 1 0 297068 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3229
timestamp 1676037725
transform 1 0 298172 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3241
timestamp 1676037725
transform 1 0 299276 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3247
timestamp 1676037725
transform 1 0 299828 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3249
timestamp 1676037725
transform 1 0 300012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3261
timestamp 1676037725
transform 1 0 301116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3273
timestamp 1676037725
transform 1 0 302220 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3285
timestamp 1676037725
transform 1 0 303324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3297
timestamp 1676037725
transform 1 0 304428 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3303
timestamp 1676037725
transform 1 0 304980 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3305
timestamp 1676037725
transform 1 0 305164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3317
timestamp 1676037725
transform 1 0 306268 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3329
timestamp 1676037725
transform 1 0 307372 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3341
timestamp 1676037725
transform 1 0 308476 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3353
timestamp 1676037725
transform 1 0 309580 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3359
timestamp 1676037725
transform 1 0 310132 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3361
timestamp 1676037725
transform 1 0 310316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3373
timestamp 1676037725
transform 1 0 311420 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3385
timestamp 1676037725
transform 1 0 312524 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3397
timestamp 1676037725
transform 1 0 313628 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3409
timestamp 1676037725
transform 1 0 314732 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3415
timestamp 1676037725
transform 1 0 315284 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3417
timestamp 1676037725
transform 1 0 315468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3429
timestamp 1676037725
transform 1 0 316572 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3441
timestamp 1676037725
transform 1 0 317676 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3453
timestamp 1676037725
transform 1 0 318780 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3465
timestamp 1676037725
transform 1 0 319884 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3471
timestamp 1676037725
transform 1 0 320436 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3473
timestamp 1676037725
transform 1 0 320620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3485
timestamp 1676037725
transform 1 0 321724 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3497
timestamp 1676037725
transform 1 0 322828 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3509
timestamp 1676037725
transform 1 0 323932 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3521
timestamp 1676037725
transform 1 0 325036 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3527
timestamp 1676037725
transform 1 0 325588 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3529
timestamp 1676037725
transform 1 0 325772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3541
timestamp 1676037725
transform 1 0 326876 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3553
timestamp 1676037725
transform 1 0 327980 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3565
timestamp 1676037725
transform 1 0 329084 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3577
timestamp 1676037725
transform 1 0 330188 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3583
timestamp 1676037725
transform 1 0 330740 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3585
timestamp 1676037725
transform 1 0 330924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3597
timestamp 1676037725
transform 1 0 332028 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3609
timestamp 1676037725
transform 1 0 333132 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3621
timestamp 1676037725
transform 1 0 334236 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3633
timestamp 1676037725
transform 1 0 335340 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3639
timestamp 1676037725
transform 1 0 335892 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3641
timestamp 1676037725
transform 1 0 336076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3653
timestamp 1676037725
transform 1 0 337180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3665
timestamp 1676037725
transform 1 0 338284 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3677
timestamp 1676037725
transform 1 0 339388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3689
timestamp 1676037725
transform 1 0 340492 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3695
timestamp 1676037725
transform 1 0 341044 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3697
timestamp 1676037725
transform 1 0 341228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3709
timestamp 1676037725
transform 1 0 342332 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3721
timestamp 1676037725
transform 1 0 343436 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3733
timestamp 1676037725
transform 1 0 344540 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3745
timestamp 1676037725
transform 1 0 345644 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3751
timestamp 1676037725
transform 1 0 346196 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3753
timestamp 1676037725
transform 1 0 346380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3765
timestamp 1676037725
transform 1 0 347484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3777
timestamp 1676037725
transform 1 0 348588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3789
timestamp 1676037725
transform 1 0 349692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3801
timestamp 1676037725
transform 1 0 350796 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3807
timestamp 1676037725
transform 1 0 351348 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3809
timestamp 1676037725
transform 1 0 351532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3821
timestamp 1676037725
transform 1 0 352636 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3833
timestamp 1676037725
transform 1 0 353740 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3845
timestamp 1676037725
transform 1 0 354844 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3857
timestamp 1676037725
transform 1 0 355948 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3863
timestamp 1676037725
transform 1 0 356500 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3865
timestamp 1676037725
transform 1 0 356684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3877
timestamp 1676037725
transform 1 0 357788 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3889
timestamp 1676037725
transform 1 0 358892 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3901
timestamp 1676037725
transform 1 0 359996 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3913
timestamp 1676037725
transform 1 0 361100 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3919
timestamp 1676037725
transform 1 0 361652 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3921
timestamp 1676037725
transform 1 0 361836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3933
timestamp 1676037725
transform 1 0 362940 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3945
timestamp 1676037725
transform 1 0 364044 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3957
timestamp 1676037725
transform 1 0 365148 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3969
timestamp 1676037725
transform 1 0 366252 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3975
timestamp 1676037725
transform 1 0 366804 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3977
timestamp 1676037725
transform 1 0 366988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3989
timestamp 1676037725
transform 1 0 368092 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4001
timestamp 1676037725
transform 1 0 369196 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4013
timestamp 1676037725
transform 1 0 370300 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4025
timestamp 1676037725
transform 1 0 371404 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4031
timestamp 1676037725
transform 1 0 371956 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4033
timestamp 1676037725
transform 1 0 372140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4045
timestamp 1676037725
transform 1 0 373244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4057
timestamp 1676037725
transform 1 0 374348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4069
timestamp 1676037725
transform 1 0 375452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4081
timestamp 1676037725
transform 1 0 376556 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4087
timestamp 1676037725
transform 1 0 377108 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4089
timestamp 1676037725
transform 1 0 377292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4101
timestamp 1676037725
transform 1 0 378396 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4113
timestamp 1676037725
transform 1 0 379500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4125
timestamp 1676037725
transform 1 0 380604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4137
timestamp 1676037725
transform 1 0 381708 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4143
timestamp 1676037725
transform 1 0 382260 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4145
timestamp 1676037725
transform 1 0 382444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4157
timestamp 1676037725
transform 1 0 383548 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4169
timestamp 1676037725
transform 1 0 384652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4181
timestamp 1676037725
transform 1 0 385756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4193
timestamp 1676037725
transform 1 0 386860 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4199
timestamp 1676037725
transform 1 0 387412 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4201
timestamp 1676037725
transform 1 0 387596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4213
timestamp 1676037725
transform 1 0 388700 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4225
timestamp 1676037725
transform 1 0 389804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4237
timestamp 1676037725
transform 1 0 390908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4249
timestamp 1676037725
transform 1 0 392012 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4255
timestamp 1676037725
transform 1 0 392564 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4257
timestamp 1676037725
transform 1 0 392748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4269
timestamp 1676037725
transform 1 0 393852 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4281
timestamp 1676037725
transform 1 0 394956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4293
timestamp 1676037725
transform 1 0 396060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4305
timestamp 1676037725
transform 1 0 397164 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4311
timestamp 1676037725
transform 1 0 397716 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4313
timestamp 1676037725
transform 1 0 397900 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4325
timestamp 1676037725
transform 1 0 399004 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4337
timestamp 1676037725
transform 1 0 400108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4349
timestamp 1676037725
transform 1 0 401212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4361
timestamp 1676037725
transform 1 0 402316 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4367
timestamp 1676037725
transform 1 0 402868 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4369
timestamp 1676037725
transform 1 0 403052 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4381
timestamp 1676037725
transform 1 0 404156 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4393
timestamp 1676037725
transform 1 0 405260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4405
timestamp 1676037725
transform 1 0 406364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4417
timestamp 1676037725
transform 1 0 407468 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4423
timestamp 1676037725
transform 1 0 408020 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4425
timestamp 1676037725
transform 1 0 408204 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4437
timestamp 1676037725
transform 1 0 409308 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4449
timestamp 1676037725
transform 1 0 410412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4461
timestamp 1676037725
transform 1 0 411516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4473
timestamp 1676037725
transform 1 0 412620 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4479
timestamp 1676037725
transform 1 0 413172 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4481
timestamp 1676037725
transform 1 0 413356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4493
timestamp 1676037725
transform 1 0 414460 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4505
timestamp 1676037725
transform 1 0 415564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4517
timestamp 1676037725
transform 1 0 416668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4529
timestamp 1676037725
transform 1 0 417772 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4535
timestamp 1676037725
transform 1 0 418324 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4537
timestamp 1676037725
transform 1 0 418508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4549
timestamp 1676037725
transform 1 0 419612 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4561
timestamp 1676037725
transform 1 0 420716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4573
timestamp 1676037725
transform 1 0 421820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4585
timestamp 1676037725
transform 1 0 422924 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4591
timestamp 1676037725
transform 1 0 423476 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4593
timestamp 1676037725
transform 1 0 423660 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4605
timestamp 1676037725
transform 1 0 424764 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4617
timestamp 1676037725
transform 1 0 425868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4629
timestamp 1676037725
transform 1 0 426972 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4641
timestamp 1676037725
transform 1 0 428076 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4647
timestamp 1676037725
transform 1 0 428628 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4649
timestamp 1676037725
transform 1 0 428812 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4661
timestamp 1676037725
transform 1 0 429916 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4673
timestamp 1676037725
transform 1 0 431020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4685
timestamp 1676037725
transform 1 0 432124 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4697
timestamp 1676037725
transform 1 0 433228 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4703
timestamp 1676037725
transform 1 0 433780 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4705
timestamp 1676037725
transform 1 0 433964 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4717
timestamp 1676037725
transform 1 0 435068 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4729
timestamp 1676037725
transform 1 0 436172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4741
timestamp 1676037725
transform 1 0 437276 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4753
timestamp 1676037725
transform 1 0 438380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4759
timestamp 1676037725
transform 1 0 438932 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4761
timestamp 1676037725
transform 1 0 439116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4773
timestamp 1676037725
transform 1 0 440220 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4785
timestamp 1676037725
transform 1 0 441324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4797
timestamp 1676037725
transform 1 0 442428 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4809
timestamp 1676037725
transform 1 0 443532 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4815
timestamp 1676037725
transform 1 0 444084 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4817
timestamp 1676037725
transform 1 0 444268 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4829
timestamp 1676037725
transform 1 0 445372 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4841
timestamp 1676037725
transform 1 0 446476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4853
timestamp 1676037725
transform 1 0 447580 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4865
timestamp 1676037725
transform 1 0 448684 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4871
timestamp 1676037725
transform 1 0 449236 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4873
timestamp 1676037725
transform 1 0 449420 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4885
timestamp 1676037725
transform 1 0 450524 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4897
timestamp 1676037725
transform 1 0 451628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4909
timestamp 1676037725
transform 1 0 452732 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4921
timestamp 1676037725
transform 1 0 453836 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4927
timestamp 1676037725
transform 1 0 454388 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4929
timestamp 1676037725
transform 1 0 454572 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4941
timestamp 1676037725
transform 1 0 455676 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4953
timestamp 1676037725
transform 1 0 456780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4965
timestamp 1676037725
transform 1 0 457884 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4977
timestamp 1676037725
transform 1 0 458988 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4983
timestamp 1676037725
transform 1 0 459540 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4985
timestamp 1676037725
transform 1 0 459724 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4997
timestamp 1676037725
transform 1 0 460828 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5009
timestamp 1676037725
transform 1 0 461932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5021
timestamp 1676037725
transform 1 0 463036 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5033
timestamp 1676037725
transform 1 0 464140 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5039
timestamp 1676037725
transform 1 0 464692 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5041
timestamp 1676037725
transform 1 0 464876 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5053
timestamp 1676037725
transform 1 0 465980 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5065
timestamp 1676037725
transform 1 0 467084 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5077
timestamp 1676037725
transform 1 0 468188 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5089
timestamp 1676037725
transform 1 0 469292 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5095
timestamp 1676037725
transform 1 0 469844 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5097
timestamp 1676037725
transform 1 0 470028 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5109
timestamp 1676037725
transform 1 0 471132 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5121
timestamp 1676037725
transform 1 0 472236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5133
timestamp 1676037725
transform 1 0 473340 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5145
timestamp 1676037725
transform 1 0 474444 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5151
timestamp 1676037725
transform 1 0 474996 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5153
timestamp 1676037725
transform 1 0 475180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5165
timestamp 1676037725
transform 1 0 476284 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5177
timestamp 1676037725
transform 1 0 477388 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5189
timestamp 1676037725
transform 1 0 478492 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5201
timestamp 1676037725
transform 1 0 479596 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5207
timestamp 1676037725
transform 1 0 480148 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5209
timestamp 1676037725
transform 1 0 480332 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5221
timestamp 1676037725
transform 1 0 481436 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5233
timestamp 1676037725
transform 1 0 482540 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5245
timestamp 1676037725
transform 1 0 483644 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5257
timestamp 1676037725
transform 1 0 484748 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5263
timestamp 1676037725
transform 1 0 485300 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5265
timestamp 1676037725
transform 1 0 485484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5277
timestamp 1676037725
transform 1 0 486588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5289
timestamp 1676037725
transform 1 0 487692 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5301
timestamp 1676037725
transform 1 0 488796 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5313
timestamp 1676037725
transform 1 0 489900 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5319
timestamp 1676037725
transform 1 0 490452 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5321
timestamp 1676037725
transform 1 0 490636 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5333
timestamp 1676037725
transform 1 0 491740 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5345
timestamp 1676037725
transform 1 0 492844 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5357
timestamp 1676037725
transform 1 0 493948 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5369
timestamp 1676037725
transform 1 0 495052 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5375
timestamp 1676037725
transform 1 0 495604 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5377
timestamp 1676037725
transform 1 0 495788 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5389
timestamp 1676037725
transform 1 0 496892 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5401
timestamp 1676037725
transform 1 0 497996 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5413
timestamp 1676037725
transform 1 0 499100 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5425
timestamp 1676037725
transform 1 0 500204 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5431
timestamp 1676037725
transform 1 0 500756 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5433
timestamp 1676037725
transform 1 0 500940 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5445
timestamp 1676037725
transform 1 0 502044 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5457
timestamp 1676037725
transform 1 0 503148 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5469
timestamp 1676037725
transform 1 0 504252 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5481
timestamp 1676037725
transform 1 0 505356 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5487
timestamp 1676037725
transform 1 0 505908 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5489
timestamp 1676037725
transform 1 0 506092 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5501
timestamp 1676037725
transform 1 0 507196 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5513
timestamp 1676037725
transform 1 0 508300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5525
timestamp 1676037725
transform 1 0 509404 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5537
timestamp 1676037725
transform 1 0 510508 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5543
timestamp 1676037725
transform 1 0 511060 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5545
timestamp 1676037725
transform 1 0 511244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5557
timestamp 1676037725
transform 1 0 512348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5569
timestamp 1676037725
transform 1 0 513452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5581
timestamp 1676037725
transform 1 0 514556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5593
timestamp 1676037725
transform 1 0 515660 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5599
timestamp 1676037725
transform 1 0 516212 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5601
timestamp 1676037725
transform 1 0 516396 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5613
timestamp 1676037725
transform 1 0 517500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5625
timestamp 1676037725
transform 1 0 518604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5637
timestamp 1676037725
transform 1 0 519708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5649
timestamp 1676037725
transform 1 0 520812 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5655
timestamp 1676037725
transform 1 0 521364 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5657
timestamp 1676037725
transform 1 0 521548 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5669
timestamp 1676037725
transform 1 0 522652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5681
timestamp 1676037725
transform 1 0 523756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5693
timestamp 1676037725
transform 1 0 524860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5705
timestamp 1676037725
transform 1 0 525964 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5711
timestamp 1676037725
transform 1 0 526516 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5713
timestamp 1676037725
transform 1 0 526700 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_5725
timestamp 1676037725
transform 1 0 527804 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1676037725
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1676037725
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1676037725
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1676037725
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1676037725
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1676037725
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1676037725
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1676037725
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1676037725
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1676037725
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1676037725
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1676037725
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1676037725
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1676037725
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1676037725
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1676037725
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1676037725
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1676037725
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1676037725
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1676037725
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1676037725
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1676037725
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1676037725
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1676037725
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1676037725
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1676037725
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1676037725
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1676037725
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1676037725
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1676037725
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1676037725
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_725
timestamp 1676037725
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_737
timestamp 1676037725
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1676037725
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1676037725
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_757
timestamp 1676037725
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_769
timestamp 1676037725
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_781
timestamp 1676037725
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_793
timestamp 1676037725
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1676037725
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1676037725
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_813
timestamp 1676037725
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_825
timestamp 1676037725
transform 1 0 77004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_837
timestamp 1676037725
transform 1 0 78108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_849
timestamp 1676037725
transform 1 0 79212 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_861
timestamp 1676037725
transform 1 0 80316 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_867
timestamp 1676037725
transform 1 0 80868 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_869
timestamp 1676037725
transform 1 0 81052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_881
timestamp 1676037725
transform 1 0 82156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_893
timestamp 1676037725
transform 1 0 83260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_905
timestamp 1676037725
transform 1 0 84364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_917
timestamp 1676037725
transform 1 0 85468 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_923
timestamp 1676037725
transform 1 0 86020 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_925
timestamp 1676037725
transform 1 0 86204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_937
timestamp 1676037725
transform 1 0 87308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_949
timestamp 1676037725
transform 1 0 88412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_961
timestamp 1676037725
transform 1 0 89516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_973
timestamp 1676037725
transform 1 0 90620 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_979
timestamp 1676037725
transform 1 0 91172 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_981
timestamp 1676037725
transform 1 0 91356 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_993
timestamp 1676037725
transform 1 0 92460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1005
timestamp 1676037725
transform 1 0 93564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1017
timestamp 1676037725
transform 1 0 94668 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1029
timestamp 1676037725
transform 1 0 95772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1035
timestamp 1676037725
transform 1 0 96324 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1037
timestamp 1676037725
transform 1 0 96508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1049
timestamp 1676037725
transform 1 0 97612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1061
timestamp 1676037725
transform 1 0 98716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1073
timestamp 1676037725
transform 1 0 99820 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1085
timestamp 1676037725
transform 1 0 100924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1091
timestamp 1676037725
transform 1 0 101476 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1093
timestamp 1676037725
transform 1 0 101660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1105
timestamp 1676037725
transform 1 0 102764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1117
timestamp 1676037725
transform 1 0 103868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1129
timestamp 1676037725
transform 1 0 104972 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1141
timestamp 1676037725
transform 1 0 106076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1147
timestamp 1676037725
transform 1 0 106628 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1149
timestamp 1676037725
transform 1 0 106812 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1161
timestamp 1676037725
transform 1 0 107916 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1173
timestamp 1676037725
transform 1 0 109020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1185
timestamp 1676037725
transform 1 0 110124 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1197
timestamp 1676037725
transform 1 0 111228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1203
timestamp 1676037725
transform 1 0 111780 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1205
timestamp 1676037725
transform 1 0 111964 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1217
timestamp 1676037725
transform 1 0 113068 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1229
timestamp 1676037725
transform 1 0 114172 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1241
timestamp 1676037725
transform 1 0 115276 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1253
timestamp 1676037725
transform 1 0 116380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1259
timestamp 1676037725
transform 1 0 116932 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1261
timestamp 1676037725
transform 1 0 117116 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1273
timestamp 1676037725
transform 1 0 118220 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1285
timestamp 1676037725
transform 1 0 119324 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1297
timestamp 1676037725
transform 1 0 120428 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1309
timestamp 1676037725
transform 1 0 121532 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1315
timestamp 1676037725
transform 1 0 122084 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1317
timestamp 1676037725
transform 1 0 122268 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1329
timestamp 1676037725
transform 1 0 123372 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1341
timestamp 1676037725
transform 1 0 124476 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1353
timestamp 1676037725
transform 1 0 125580 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1365
timestamp 1676037725
transform 1 0 126684 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1371
timestamp 1676037725
transform 1 0 127236 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1373
timestamp 1676037725
transform 1 0 127420 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1385
timestamp 1676037725
transform 1 0 128524 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1397
timestamp 1676037725
transform 1 0 129628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1409
timestamp 1676037725
transform 1 0 130732 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1421
timestamp 1676037725
transform 1 0 131836 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1427
timestamp 1676037725
transform 1 0 132388 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1429
timestamp 1676037725
transform 1 0 132572 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1441
timestamp 1676037725
transform 1 0 133676 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1453
timestamp 1676037725
transform 1 0 134780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1465
timestamp 1676037725
transform 1 0 135884 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1477
timestamp 1676037725
transform 1 0 136988 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1483
timestamp 1676037725
transform 1 0 137540 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1485
timestamp 1676037725
transform 1 0 137724 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1497
timestamp 1676037725
transform 1 0 138828 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1509
timestamp 1676037725
transform 1 0 139932 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1521
timestamp 1676037725
transform 1 0 141036 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1533
timestamp 1676037725
transform 1 0 142140 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1539
timestamp 1676037725
transform 1 0 142692 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1541
timestamp 1676037725
transform 1 0 142876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1553
timestamp 1676037725
transform 1 0 143980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1565
timestamp 1676037725
transform 1 0 145084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1577
timestamp 1676037725
transform 1 0 146188 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1589
timestamp 1676037725
transform 1 0 147292 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1595
timestamp 1676037725
transform 1 0 147844 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1597
timestamp 1676037725
transform 1 0 148028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1609
timestamp 1676037725
transform 1 0 149132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1621
timestamp 1676037725
transform 1 0 150236 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1633
timestamp 1676037725
transform 1 0 151340 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1645
timestamp 1676037725
transform 1 0 152444 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1651
timestamp 1676037725
transform 1 0 152996 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1653
timestamp 1676037725
transform 1 0 153180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1665
timestamp 1676037725
transform 1 0 154284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1677
timestamp 1676037725
transform 1 0 155388 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1689
timestamp 1676037725
transform 1 0 156492 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1701
timestamp 1676037725
transform 1 0 157596 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1707
timestamp 1676037725
transform 1 0 158148 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1709
timestamp 1676037725
transform 1 0 158332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1721
timestamp 1676037725
transform 1 0 159436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1733
timestamp 1676037725
transform 1 0 160540 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1745
timestamp 1676037725
transform 1 0 161644 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1757
timestamp 1676037725
transform 1 0 162748 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1763
timestamp 1676037725
transform 1 0 163300 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1765
timestamp 1676037725
transform 1 0 163484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1777
timestamp 1676037725
transform 1 0 164588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1789
timestamp 1676037725
transform 1 0 165692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1801
timestamp 1676037725
transform 1 0 166796 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1813
timestamp 1676037725
transform 1 0 167900 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1819
timestamp 1676037725
transform 1 0 168452 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1821
timestamp 1676037725
transform 1 0 168636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1833
timestamp 1676037725
transform 1 0 169740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1845
timestamp 1676037725
transform 1 0 170844 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1857
timestamp 1676037725
transform 1 0 171948 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1869
timestamp 1676037725
transform 1 0 173052 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1875
timestamp 1676037725
transform 1 0 173604 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1877
timestamp 1676037725
transform 1 0 173788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1889
timestamp 1676037725
transform 1 0 174892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1901
timestamp 1676037725
transform 1 0 175996 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1913
timestamp 1676037725
transform 1 0 177100 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1925
timestamp 1676037725
transform 1 0 178204 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1931
timestamp 1676037725
transform 1 0 178756 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1933
timestamp 1676037725
transform 1 0 178940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1945
timestamp 1676037725
transform 1 0 180044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1957
timestamp 1676037725
transform 1 0 181148 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1969
timestamp 1676037725
transform 1 0 182252 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1981
timestamp 1676037725
transform 1 0 183356 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1987
timestamp 1676037725
transform 1 0 183908 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1989
timestamp 1676037725
transform 1 0 184092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2001
timestamp 1676037725
transform 1 0 185196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2013
timestamp 1676037725
transform 1 0 186300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2025
timestamp 1676037725
transform 1 0 187404 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2037
timestamp 1676037725
transform 1 0 188508 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2043
timestamp 1676037725
transform 1 0 189060 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2045
timestamp 1676037725
transform 1 0 189244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2057
timestamp 1676037725
transform 1 0 190348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2069
timestamp 1676037725
transform 1 0 191452 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2081
timestamp 1676037725
transform 1 0 192556 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2093
timestamp 1676037725
transform 1 0 193660 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2099
timestamp 1676037725
transform 1 0 194212 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2101
timestamp 1676037725
transform 1 0 194396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2113
timestamp 1676037725
transform 1 0 195500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2125
timestamp 1676037725
transform 1 0 196604 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2137
timestamp 1676037725
transform 1 0 197708 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2149
timestamp 1676037725
transform 1 0 198812 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2155
timestamp 1676037725
transform 1 0 199364 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2157
timestamp 1676037725
transform 1 0 199548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2169
timestamp 1676037725
transform 1 0 200652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2181
timestamp 1676037725
transform 1 0 201756 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2193
timestamp 1676037725
transform 1 0 202860 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2205
timestamp 1676037725
transform 1 0 203964 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2211
timestamp 1676037725
transform 1 0 204516 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2213
timestamp 1676037725
transform 1 0 204700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2225
timestamp 1676037725
transform 1 0 205804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2237
timestamp 1676037725
transform 1 0 206908 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2249
timestamp 1676037725
transform 1 0 208012 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2261
timestamp 1676037725
transform 1 0 209116 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2267
timestamp 1676037725
transform 1 0 209668 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2269
timestamp 1676037725
transform 1 0 209852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2281
timestamp 1676037725
transform 1 0 210956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2293
timestamp 1676037725
transform 1 0 212060 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2305
timestamp 1676037725
transform 1 0 213164 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2317
timestamp 1676037725
transform 1 0 214268 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2323
timestamp 1676037725
transform 1 0 214820 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2325
timestamp 1676037725
transform 1 0 215004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2337
timestamp 1676037725
transform 1 0 216108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2349
timestamp 1676037725
transform 1 0 217212 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2361
timestamp 1676037725
transform 1 0 218316 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2373
timestamp 1676037725
transform 1 0 219420 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2379
timestamp 1676037725
transform 1 0 219972 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2381
timestamp 1676037725
transform 1 0 220156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2393
timestamp 1676037725
transform 1 0 221260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2405
timestamp 1676037725
transform 1 0 222364 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2417
timestamp 1676037725
transform 1 0 223468 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2429
timestamp 1676037725
transform 1 0 224572 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2435
timestamp 1676037725
transform 1 0 225124 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2437
timestamp 1676037725
transform 1 0 225308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2449
timestamp 1676037725
transform 1 0 226412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2461
timestamp 1676037725
transform 1 0 227516 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2473
timestamp 1676037725
transform 1 0 228620 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2485
timestamp 1676037725
transform 1 0 229724 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2491
timestamp 1676037725
transform 1 0 230276 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2493
timestamp 1676037725
transform 1 0 230460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2505
timestamp 1676037725
transform 1 0 231564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2517
timestamp 1676037725
transform 1 0 232668 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2529
timestamp 1676037725
transform 1 0 233772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2541
timestamp 1676037725
transform 1 0 234876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2547
timestamp 1676037725
transform 1 0 235428 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2549
timestamp 1676037725
transform 1 0 235612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2561
timestamp 1676037725
transform 1 0 236716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2573
timestamp 1676037725
transform 1 0 237820 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2585
timestamp 1676037725
transform 1 0 238924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2597
timestamp 1676037725
transform 1 0 240028 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2603
timestamp 1676037725
transform 1 0 240580 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2605
timestamp 1676037725
transform 1 0 240764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2617
timestamp 1676037725
transform 1 0 241868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2629
timestamp 1676037725
transform 1 0 242972 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2641
timestamp 1676037725
transform 1 0 244076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2653
timestamp 1676037725
transform 1 0 245180 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2659
timestamp 1676037725
transform 1 0 245732 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2661
timestamp 1676037725
transform 1 0 245916 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2673
timestamp 1676037725
transform 1 0 247020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2685
timestamp 1676037725
transform 1 0 248124 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2697
timestamp 1676037725
transform 1 0 249228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2709
timestamp 1676037725
transform 1 0 250332 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2715
timestamp 1676037725
transform 1 0 250884 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2717
timestamp 1676037725
transform 1 0 251068 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2729
timestamp 1676037725
transform 1 0 252172 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2741
timestamp 1676037725
transform 1 0 253276 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2753
timestamp 1676037725
transform 1 0 254380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2765
timestamp 1676037725
transform 1 0 255484 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2771
timestamp 1676037725
transform 1 0 256036 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2773
timestamp 1676037725
transform 1 0 256220 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2785
timestamp 1676037725
transform 1 0 257324 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2797
timestamp 1676037725
transform 1 0 258428 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2809
timestamp 1676037725
transform 1 0 259532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2821
timestamp 1676037725
transform 1 0 260636 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2827
timestamp 1676037725
transform 1 0 261188 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2829
timestamp 1676037725
transform 1 0 261372 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2841
timestamp 1676037725
transform 1 0 262476 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2853
timestamp 1676037725
transform 1 0 263580 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2865
timestamp 1676037725
transform 1 0 264684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2877
timestamp 1676037725
transform 1 0 265788 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2883
timestamp 1676037725
transform 1 0 266340 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2885
timestamp 1676037725
transform 1 0 266524 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2897
timestamp 1676037725
transform 1 0 267628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2909
timestamp 1676037725
transform 1 0 268732 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2921
timestamp 1676037725
transform 1 0 269836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2933
timestamp 1676037725
transform 1 0 270940 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2939
timestamp 1676037725
transform 1 0 271492 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2941
timestamp 1676037725
transform 1 0 271676 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2953
timestamp 1676037725
transform 1 0 272780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2965
timestamp 1676037725
transform 1 0 273884 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2977
timestamp 1676037725
transform 1 0 274988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2989
timestamp 1676037725
transform 1 0 276092 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2995
timestamp 1676037725
transform 1 0 276644 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2997
timestamp 1676037725
transform 1 0 276828 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3009
timestamp 1676037725
transform 1 0 277932 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3021
timestamp 1676037725
transform 1 0 279036 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3033
timestamp 1676037725
transform 1 0 280140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3045
timestamp 1676037725
transform 1 0 281244 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3051
timestamp 1676037725
transform 1 0 281796 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3053
timestamp 1676037725
transform 1 0 281980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3065
timestamp 1676037725
transform 1 0 283084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3077
timestamp 1676037725
transform 1 0 284188 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3089
timestamp 1676037725
transform 1 0 285292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3101
timestamp 1676037725
transform 1 0 286396 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3107
timestamp 1676037725
transform 1 0 286948 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3109
timestamp 1676037725
transform 1 0 287132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3121
timestamp 1676037725
transform 1 0 288236 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3133
timestamp 1676037725
transform 1 0 289340 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3145
timestamp 1676037725
transform 1 0 290444 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3157
timestamp 1676037725
transform 1 0 291548 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3163
timestamp 1676037725
transform 1 0 292100 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3165
timestamp 1676037725
transform 1 0 292284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3177
timestamp 1676037725
transform 1 0 293388 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3189
timestamp 1676037725
transform 1 0 294492 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3201
timestamp 1676037725
transform 1 0 295596 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3213
timestamp 1676037725
transform 1 0 296700 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3219
timestamp 1676037725
transform 1 0 297252 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3221
timestamp 1676037725
transform 1 0 297436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3233
timestamp 1676037725
transform 1 0 298540 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3245
timestamp 1676037725
transform 1 0 299644 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3257
timestamp 1676037725
transform 1 0 300748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3269
timestamp 1676037725
transform 1 0 301852 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3275
timestamp 1676037725
transform 1 0 302404 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3277
timestamp 1676037725
transform 1 0 302588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3289
timestamp 1676037725
transform 1 0 303692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3301
timestamp 1676037725
transform 1 0 304796 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3313
timestamp 1676037725
transform 1 0 305900 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3325
timestamp 1676037725
transform 1 0 307004 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3331
timestamp 1676037725
transform 1 0 307556 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3333
timestamp 1676037725
transform 1 0 307740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3345
timestamp 1676037725
transform 1 0 308844 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3357
timestamp 1676037725
transform 1 0 309948 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3369
timestamp 1676037725
transform 1 0 311052 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3381
timestamp 1676037725
transform 1 0 312156 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3387
timestamp 1676037725
transform 1 0 312708 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3389
timestamp 1676037725
transform 1 0 312892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3401
timestamp 1676037725
transform 1 0 313996 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3413
timestamp 1676037725
transform 1 0 315100 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3425
timestamp 1676037725
transform 1 0 316204 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3437
timestamp 1676037725
transform 1 0 317308 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3443
timestamp 1676037725
transform 1 0 317860 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3445
timestamp 1676037725
transform 1 0 318044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3457
timestamp 1676037725
transform 1 0 319148 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3469
timestamp 1676037725
transform 1 0 320252 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3481
timestamp 1676037725
transform 1 0 321356 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3493
timestamp 1676037725
transform 1 0 322460 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3499
timestamp 1676037725
transform 1 0 323012 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3501
timestamp 1676037725
transform 1 0 323196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3513
timestamp 1676037725
transform 1 0 324300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3525
timestamp 1676037725
transform 1 0 325404 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3537
timestamp 1676037725
transform 1 0 326508 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3549
timestamp 1676037725
transform 1 0 327612 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3555
timestamp 1676037725
transform 1 0 328164 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3557
timestamp 1676037725
transform 1 0 328348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3569
timestamp 1676037725
transform 1 0 329452 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3581
timestamp 1676037725
transform 1 0 330556 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3593
timestamp 1676037725
transform 1 0 331660 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3605
timestamp 1676037725
transform 1 0 332764 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3611
timestamp 1676037725
transform 1 0 333316 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3613
timestamp 1676037725
transform 1 0 333500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3625
timestamp 1676037725
transform 1 0 334604 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3637
timestamp 1676037725
transform 1 0 335708 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3649
timestamp 1676037725
transform 1 0 336812 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3661
timestamp 1676037725
transform 1 0 337916 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3667
timestamp 1676037725
transform 1 0 338468 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3669
timestamp 1676037725
transform 1 0 338652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3681
timestamp 1676037725
transform 1 0 339756 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3693
timestamp 1676037725
transform 1 0 340860 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3705
timestamp 1676037725
transform 1 0 341964 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3717
timestamp 1676037725
transform 1 0 343068 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3723
timestamp 1676037725
transform 1 0 343620 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3725
timestamp 1676037725
transform 1 0 343804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3737
timestamp 1676037725
transform 1 0 344908 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3749
timestamp 1676037725
transform 1 0 346012 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3761
timestamp 1676037725
transform 1 0 347116 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3773
timestamp 1676037725
transform 1 0 348220 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3779
timestamp 1676037725
transform 1 0 348772 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3781
timestamp 1676037725
transform 1 0 348956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3793
timestamp 1676037725
transform 1 0 350060 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3805
timestamp 1676037725
transform 1 0 351164 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3817
timestamp 1676037725
transform 1 0 352268 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3829
timestamp 1676037725
transform 1 0 353372 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3835
timestamp 1676037725
transform 1 0 353924 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3837
timestamp 1676037725
transform 1 0 354108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3849
timestamp 1676037725
transform 1 0 355212 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3861
timestamp 1676037725
transform 1 0 356316 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3873
timestamp 1676037725
transform 1 0 357420 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3885
timestamp 1676037725
transform 1 0 358524 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3891
timestamp 1676037725
transform 1 0 359076 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3893
timestamp 1676037725
transform 1 0 359260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3905
timestamp 1676037725
transform 1 0 360364 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3917
timestamp 1676037725
transform 1 0 361468 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3929
timestamp 1676037725
transform 1 0 362572 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3941
timestamp 1676037725
transform 1 0 363676 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3947
timestamp 1676037725
transform 1 0 364228 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3949
timestamp 1676037725
transform 1 0 364412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3961
timestamp 1676037725
transform 1 0 365516 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3973
timestamp 1676037725
transform 1 0 366620 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3985
timestamp 1676037725
transform 1 0 367724 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3997
timestamp 1676037725
transform 1 0 368828 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4003
timestamp 1676037725
transform 1 0 369380 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4005
timestamp 1676037725
transform 1 0 369564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4017
timestamp 1676037725
transform 1 0 370668 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4029
timestamp 1676037725
transform 1 0 371772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4041
timestamp 1676037725
transform 1 0 372876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4053
timestamp 1676037725
transform 1 0 373980 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4059
timestamp 1676037725
transform 1 0 374532 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4061
timestamp 1676037725
transform 1 0 374716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4073
timestamp 1676037725
transform 1 0 375820 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4085
timestamp 1676037725
transform 1 0 376924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4097
timestamp 1676037725
transform 1 0 378028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4109
timestamp 1676037725
transform 1 0 379132 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4115
timestamp 1676037725
transform 1 0 379684 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4117
timestamp 1676037725
transform 1 0 379868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4129
timestamp 1676037725
transform 1 0 380972 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4141
timestamp 1676037725
transform 1 0 382076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4153
timestamp 1676037725
transform 1 0 383180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4165
timestamp 1676037725
transform 1 0 384284 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4171
timestamp 1676037725
transform 1 0 384836 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4173
timestamp 1676037725
transform 1 0 385020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4185
timestamp 1676037725
transform 1 0 386124 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4197
timestamp 1676037725
transform 1 0 387228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4209
timestamp 1676037725
transform 1 0 388332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4221
timestamp 1676037725
transform 1 0 389436 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4227
timestamp 1676037725
transform 1 0 389988 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4229
timestamp 1676037725
transform 1 0 390172 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4241
timestamp 1676037725
transform 1 0 391276 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4253
timestamp 1676037725
transform 1 0 392380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4265
timestamp 1676037725
transform 1 0 393484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4277
timestamp 1676037725
transform 1 0 394588 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4283
timestamp 1676037725
transform 1 0 395140 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4285
timestamp 1676037725
transform 1 0 395324 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4297
timestamp 1676037725
transform 1 0 396428 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4309
timestamp 1676037725
transform 1 0 397532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4321
timestamp 1676037725
transform 1 0 398636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4333
timestamp 1676037725
transform 1 0 399740 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4339
timestamp 1676037725
transform 1 0 400292 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4341
timestamp 1676037725
transform 1 0 400476 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4353
timestamp 1676037725
transform 1 0 401580 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4365
timestamp 1676037725
transform 1 0 402684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4377
timestamp 1676037725
transform 1 0 403788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4389
timestamp 1676037725
transform 1 0 404892 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4395
timestamp 1676037725
transform 1 0 405444 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4397
timestamp 1676037725
transform 1 0 405628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4409
timestamp 1676037725
transform 1 0 406732 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4421
timestamp 1676037725
transform 1 0 407836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4433
timestamp 1676037725
transform 1 0 408940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4445
timestamp 1676037725
transform 1 0 410044 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4451
timestamp 1676037725
transform 1 0 410596 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4453
timestamp 1676037725
transform 1 0 410780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4465
timestamp 1676037725
transform 1 0 411884 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4477
timestamp 1676037725
transform 1 0 412988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4489
timestamp 1676037725
transform 1 0 414092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4501
timestamp 1676037725
transform 1 0 415196 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4507
timestamp 1676037725
transform 1 0 415748 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4509
timestamp 1676037725
transform 1 0 415932 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4521
timestamp 1676037725
transform 1 0 417036 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4533
timestamp 1676037725
transform 1 0 418140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4545
timestamp 1676037725
transform 1 0 419244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4557
timestamp 1676037725
transform 1 0 420348 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4563
timestamp 1676037725
transform 1 0 420900 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4565
timestamp 1676037725
transform 1 0 421084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4577
timestamp 1676037725
transform 1 0 422188 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4589
timestamp 1676037725
transform 1 0 423292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4601
timestamp 1676037725
transform 1 0 424396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4613
timestamp 1676037725
transform 1 0 425500 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4619
timestamp 1676037725
transform 1 0 426052 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4621
timestamp 1676037725
transform 1 0 426236 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4633
timestamp 1676037725
transform 1 0 427340 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4645
timestamp 1676037725
transform 1 0 428444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4657
timestamp 1676037725
transform 1 0 429548 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4669
timestamp 1676037725
transform 1 0 430652 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4675
timestamp 1676037725
transform 1 0 431204 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4677
timestamp 1676037725
transform 1 0 431388 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4689
timestamp 1676037725
transform 1 0 432492 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4701
timestamp 1676037725
transform 1 0 433596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4713
timestamp 1676037725
transform 1 0 434700 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4725
timestamp 1676037725
transform 1 0 435804 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4731
timestamp 1676037725
transform 1 0 436356 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4733
timestamp 1676037725
transform 1 0 436540 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4745
timestamp 1676037725
transform 1 0 437644 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4757
timestamp 1676037725
transform 1 0 438748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4769
timestamp 1676037725
transform 1 0 439852 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4781
timestamp 1676037725
transform 1 0 440956 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4787
timestamp 1676037725
transform 1 0 441508 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4789
timestamp 1676037725
transform 1 0 441692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4801
timestamp 1676037725
transform 1 0 442796 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4813
timestamp 1676037725
transform 1 0 443900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4825
timestamp 1676037725
transform 1 0 445004 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4837
timestamp 1676037725
transform 1 0 446108 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4843
timestamp 1676037725
transform 1 0 446660 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4845
timestamp 1676037725
transform 1 0 446844 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4857
timestamp 1676037725
transform 1 0 447948 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4869
timestamp 1676037725
transform 1 0 449052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4881
timestamp 1676037725
transform 1 0 450156 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4893
timestamp 1676037725
transform 1 0 451260 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4899
timestamp 1676037725
transform 1 0 451812 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4901
timestamp 1676037725
transform 1 0 451996 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4913
timestamp 1676037725
transform 1 0 453100 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4925
timestamp 1676037725
transform 1 0 454204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4937
timestamp 1676037725
transform 1 0 455308 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4949
timestamp 1676037725
transform 1 0 456412 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4955
timestamp 1676037725
transform 1 0 456964 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4957
timestamp 1676037725
transform 1 0 457148 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4969
timestamp 1676037725
transform 1 0 458252 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4981
timestamp 1676037725
transform 1 0 459356 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4993
timestamp 1676037725
transform 1 0 460460 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5005
timestamp 1676037725
transform 1 0 461564 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5011
timestamp 1676037725
transform 1 0 462116 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5013
timestamp 1676037725
transform 1 0 462300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5025
timestamp 1676037725
transform 1 0 463404 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5037
timestamp 1676037725
transform 1 0 464508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5049
timestamp 1676037725
transform 1 0 465612 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5061
timestamp 1676037725
transform 1 0 466716 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5067
timestamp 1676037725
transform 1 0 467268 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5069
timestamp 1676037725
transform 1 0 467452 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5081
timestamp 1676037725
transform 1 0 468556 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5093
timestamp 1676037725
transform 1 0 469660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5105
timestamp 1676037725
transform 1 0 470764 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5117
timestamp 1676037725
transform 1 0 471868 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5123
timestamp 1676037725
transform 1 0 472420 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5125
timestamp 1676037725
transform 1 0 472604 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5137
timestamp 1676037725
transform 1 0 473708 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5149
timestamp 1676037725
transform 1 0 474812 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5161
timestamp 1676037725
transform 1 0 475916 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5173
timestamp 1676037725
transform 1 0 477020 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5179
timestamp 1676037725
transform 1 0 477572 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5181
timestamp 1676037725
transform 1 0 477756 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5193
timestamp 1676037725
transform 1 0 478860 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5205
timestamp 1676037725
transform 1 0 479964 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5217
timestamp 1676037725
transform 1 0 481068 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5229
timestamp 1676037725
transform 1 0 482172 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5235
timestamp 1676037725
transform 1 0 482724 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5237
timestamp 1676037725
transform 1 0 482908 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5249
timestamp 1676037725
transform 1 0 484012 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5261
timestamp 1676037725
transform 1 0 485116 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5273
timestamp 1676037725
transform 1 0 486220 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5285
timestamp 1676037725
transform 1 0 487324 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5291
timestamp 1676037725
transform 1 0 487876 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5293
timestamp 1676037725
transform 1 0 488060 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5305
timestamp 1676037725
transform 1 0 489164 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5317
timestamp 1676037725
transform 1 0 490268 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5329
timestamp 1676037725
transform 1 0 491372 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5341
timestamp 1676037725
transform 1 0 492476 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5347
timestamp 1676037725
transform 1 0 493028 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5349
timestamp 1676037725
transform 1 0 493212 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5361
timestamp 1676037725
transform 1 0 494316 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5373
timestamp 1676037725
transform 1 0 495420 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5385
timestamp 1676037725
transform 1 0 496524 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5397
timestamp 1676037725
transform 1 0 497628 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5403
timestamp 1676037725
transform 1 0 498180 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5405
timestamp 1676037725
transform 1 0 498364 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5417
timestamp 1676037725
transform 1 0 499468 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5429
timestamp 1676037725
transform 1 0 500572 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5441
timestamp 1676037725
transform 1 0 501676 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5453
timestamp 1676037725
transform 1 0 502780 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5459
timestamp 1676037725
transform 1 0 503332 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5461
timestamp 1676037725
transform 1 0 503516 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5473
timestamp 1676037725
transform 1 0 504620 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5485
timestamp 1676037725
transform 1 0 505724 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5497
timestamp 1676037725
transform 1 0 506828 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5509
timestamp 1676037725
transform 1 0 507932 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5515
timestamp 1676037725
transform 1 0 508484 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5517
timestamp 1676037725
transform 1 0 508668 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5529
timestamp 1676037725
transform 1 0 509772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5541
timestamp 1676037725
transform 1 0 510876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5553
timestamp 1676037725
transform 1 0 511980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5565
timestamp 1676037725
transform 1 0 513084 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5571
timestamp 1676037725
transform 1 0 513636 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5573
timestamp 1676037725
transform 1 0 513820 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5585
timestamp 1676037725
transform 1 0 514924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5597
timestamp 1676037725
transform 1 0 516028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5609
timestamp 1676037725
transform 1 0 517132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5621
timestamp 1676037725
transform 1 0 518236 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5627
timestamp 1676037725
transform 1 0 518788 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5629
timestamp 1676037725
transform 1 0 518972 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5641
timestamp 1676037725
transform 1 0 520076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5653
timestamp 1676037725
transform 1 0 521180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5665
timestamp 1676037725
transform 1 0 522284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5677
timestamp 1676037725
transform 1 0 523388 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5683
timestamp 1676037725
transform 1 0 523940 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5685
timestamp 1676037725
transform 1 0 524124 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5697
timestamp 1676037725
transform 1 0 525228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5709
timestamp 1676037725
transform 1 0 526332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5721
timestamp 1676037725
transform 1 0 527436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_29
timestamp 1676037725
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_41
timestamp 1676037725
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1676037725
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_85
timestamp 1676037725
transform 1 0 8924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_97
timestamp 1676037725
transform 1 0 10028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1676037725
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_141
timestamp 1676037725
transform 1 0 14076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_153
timestamp 1676037725
transform 1 0 15180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1676037725
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_197
timestamp 1676037725
transform 1 0 19228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_209
timestamp 1676037725
transform 1 0 20332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp 1676037725
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_253
timestamp 1676037725
transform 1 0 24380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_265
timestamp 1676037725
transform 1 0 25484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1676037725
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_309
timestamp 1676037725
transform 1 0 29532 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_321
timestamp 1676037725
transform 1 0 30636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp 1676037725
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1676037725
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_361
timestamp 1676037725
transform 1 0 34316 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_365
timestamp 1676037725
transform 1 0 34684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_377
timestamp 1676037725
transform 1 0 35788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_389
timestamp 1676037725
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1676037725
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_417
timestamp 1676037725
transform 1 0 39468 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_421
timestamp 1676037725
transform 1 0 39836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_433
timestamp 1676037725
transform 1 0 40940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_445
timestamp 1676037725
transform 1 0 42044 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_473
timestamp 1676037725
transform 1 0 44620 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_477
timestamp 1676037725
transform 1 0 44988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_489
timestamp 1676037725
transform 1 0 46092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_501
timestamp 1676037725
transform 1 0 47196 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1676037725
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_529
timestamp 1676037725
transform 1 0 49772 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_533
timestamp 1676037725
transform 1 0 50140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_545
timestamp 1676037725
transform 1 0 51244 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_557
timestamp 1676037725
transform 1 0 52348 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1676037725
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1676037725
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_585
timestamp 1676037725
transform 1 0 54924 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_589
timestamp 1676037725
transform 1 0 55292 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_601
timestamp 1676037725
transform 1 0 56396 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_613
timestamp 1676037725
transform 1 0 57500 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1676037725
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1676037725
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_641
timestamp 1676037725
transform 1 0 60076 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_645
timestamp 1676037725
transform 1 0 60444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_657
timestamp 1676037725
transform 1 0 61548 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_669
timestamp 1676037725
transform 1 0 62652 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1676037725
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1676037725
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_697
timestamp 1676037725
transform 1 0 65228 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_701
timestamp 1676037725
transform 1 0 65596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_713
timestamp 1676037725
transform 1 0 66700 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_725
timestamp 1676037725
transform 1 0 67804 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_729
timestamp 1676037725
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_741
timestamp 1676037725
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_753
timestamp 1676037725
transform 1 0 70380 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_757
timestamp 1676037725
transform 1 0 70748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_769
timestamp 1676037725
transform 1 0 71852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_781
timestamp 1676037725
transform 1 0 72956 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_785
timestamp 1676037725
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_797
timestamp 1676037725
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_809
timestamp 1676037725
transform 1 0 75532 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_813
timestamp 1676037725
transform 1 0 75900 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_825
timestamp 1676037725
transform 1 0 77004 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_837
timestamp 1676037725
transform 1 0 78108 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_841
timestamp 1676037725
transform 1 0 78476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_853
timestamp 1676037725
transform 1 0 79580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_865
timestamp 1676037725
transform 1 0 80684 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_869
timestamp 1676037725
transform 1 0 81052 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_881
timestamp 1676037725
transform 1 0 82156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_893
timestamp 1676037725
transform 1 0 83260 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_897
timestamp 1676037725
transform 1 0 83628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_909
timestamp 1676037725
transform 1 0 84732 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_921
timestamp 1676037725
transform 1 0 85836 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_925
timestamp 1676037725
transform 1 0 86204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_937
timestamp 1676037725
transform 1 0 87308 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_949
timestamp 1676037725
transform 1 0 88412 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_953
timestamp 1676037725
transform 1 0 88780 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_965
timestamp 1676037725
transform 1 0 89884 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_977
timestamp 1676037725
transform 1 0 90988 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_981
timestamp 1676037725
transform 1 0 91356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_993
timestamp 1676037725
transform 1 0 92460 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1005
timestamp 1676037725
transform 1 0 93564 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1009
timestamp 1676037725
transform 1 0 93932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1021
timestamp 1676037725
transform 1 0 95036 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1033
timestamp 1676037725
transform 1 0 96140 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1037
timestamp 1676037725
transform 1 0 96508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1049
timestamp 1676037725
transform 1 0 97612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1061
timestamp 1676037725
transform 1 0 98716 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1065
timestamp 1676037725
transform 1 0 99084 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1077
timestamp 1676037725
transform 1 0 100188 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1089
timestamp 1676037725
transform 1 0 101292 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1093
timestamp 1676037725
transform 1 0 101660 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1105
timestamp 1676037725
transform 1 0 102764 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1117
timestamp 1676037725
transform 1 0 103868 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1121
timestamp 1676037725
transform 1 0 104236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1133
timestamp 1676037725
transform 1 0 105340 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1145
timestamp 1676037725
transform 1 0 106444 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1149
timestamp 1676037725
transform 1 0 106812 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1161
timestamp 1676037725
transform 1 0 107916 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1173
timestamp 1676037725
transform 1 0 109020 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1177
timestamp 1676037725
transform 1 0 109388 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1189
timestamp 1676037725
transform 1 0 110492 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1201
timestamp 1676037725
transform 1 0 111596 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1205
timestamp 1676037725
transform 1 0 111964 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1217
timestamp 1676037725
transform 1 0 113068 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1229
timestamp 1676037725
transform 1 0 114172 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1233
timestamp 1676037725
transform 1 0 114540 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1245
timestamp 1676037725
transform 1 0 115644 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1257
timestamp 1676037725
transform 1 0 116748 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1261
timestamp 1676037725
transform 1 0 117116 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1273
timestamp 1676037725
transform 1 0 118220 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1285
timestamp 1676037725
transform 1 0 119324 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1289
timestamp 1676037725
transform 1 0 119692 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1301
timestamp 1676037725
transform 1 0 120796 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1313
timestamp 1676037725
transform 1 0 121900 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1317
timestamp 1676037725
transform 1 0 122268 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1329
timestamp 1676037725
transform 1 0 123372 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1341
timestamp 1676037725
transform 1 0 124476 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1345
timestamp 1676037725
transform 1 0 124844 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1357
timestamp 1676037725
transform 1 0 125948 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1369
timestamp 1676037725
transform 1 0 127052 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1373
timestamp 1676037725
transform 1 0 127420 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1385
timestamp 1676037725
transform 1 0 128524 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1397
timestamp 1676037725
transform 1 0 129628 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1401
timestamp 1676037725
transform 1 0 129996 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1413
timestamp 1676037725
transform 1 0 131100 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1425
timestamp 1676037725
transform 1 0 132204 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1429
timestamp 1676037725
transform 1 0 132572 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1441
timestamp 1676037725
transform 1 0 133676 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1453
timestamp 1676037725
transform 1 0 134780 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1457
timestamp 1676037725
transform 1 0 135148 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1469
timestamp 1676037725
transform 1 0 136252 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1481
timestamp 1676037725
transform 1 0 137356 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1485
timestamp 1676037725
transform 1 0 137724 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1497
timestamp 1676037725
transform 1 0 138828 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1509
timestamp 1676037725
transform 1 0 139932 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1513
timestamp 1676037725
transform 1 0 140300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1525
timestamp 1676037725
transform 1 0 141404 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1537
timestamp 1676037725
transform 1 0 142508 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1541
timestamp 1676037725
transform 1 0 142876 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1553
timestamp 1676037725
transform 1 0 143980 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1565
timestamp 1676037725
transform 1 0 145084 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1569
timestamp 1676037725
transform 1 0 145452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1581
timestamp 1676037725
transform 1 0 146556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1593
timestamp 1676037725
transform 1 0 147660 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1597
timestamp 1676037725
transform 1 0 148028 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1609
timestamp 1676037725
transform 1 0 149132 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1621
timestamp 1676037725
transform 1 0 150236 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1625
timestamp 1676037725
transform 1 0 150604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1637
timestamp 1676037725
transform 1 0 151708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1649
timestamp 1676037725
transform 1 0 152812 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1653
timestamp 1676037725
transform 1 0 153180 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1665
timestamp 1676037725
transform 1 0 154284 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1677
timestamp 1676037725
transform 1 0 155388 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1681
timestamp 1676037725
transform 1 0 155756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1693
timestamp 1676037725
transform 1 0 156860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1705
timestamp 1676037725
transform 1 0 157964 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1709
timestamp 1676037725
transform 1 0 158332 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1721
timestamp 1676037725
transform 1 0 159436 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1733
timestamp 1676037725
transform 1 0 160540 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1737
timestamp 1676037725
transform 1 0 160908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1749
timestamp 1676037725
transform 1 0 162012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1761
timestamp 1676037725
transform 1 0 163116 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1765
timestamp 1676037725
transform 1 0 163484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1777
timestamp 1676037725
transform 1 0 164588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1789
timestamp 1676037725
transform 1 0 165692 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1793
timestamp 1676037725
transform 1 0 166060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1805
timestamp 1676037725
transform 1 0 167164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1817
timestamp 1676037725
transform 1 0 168268 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1821
timestamp 1676037725
transform 1 0 168636 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1833
timestamp 1676037725
transform 1 0 169740 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1845
timestamp 1676037725
transform 1 0 170844 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1849
timestamp 1676037725
transform 1 0 171212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1861
timestamp 1676037725
transform 1 0 172316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1873
timestamp 1676037725
transform 1 0 173420 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1877
timestamp 1676037725
transform 1 0 173788 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1889
timestamp 1676037725
transform 1 0 174892 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1901
timestamp 1676037725
transform 1 0 175996 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1905
timestamp 1676037725
transform 1 0 176364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1917
timestamp 1676037725
transform 1 0 177468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1929
timestamp 1676037725
transform 1 0 178572 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1933
timestamp 1676037725
transform 1 0 178940 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1945
timestamp 1676037725
transform 1 0 180044 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1957
timestamp 1676037725
transform 1 0 181148 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1961
timestamp 1676037725
transform 1 0 181516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1973
timestamp 1676037725
transform 1 0 182620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1985
timestamp 1676037725
transform 1 0 183724 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1989
timestamp 1676037725
transform 1 0 184092 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2001
timestamp 1676037725
transform 1 0 185196 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2013
timestamp 1676037725
transform 1 0 186300 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2017
timestamp 1676037725
transform 1 0 186668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2029
timestamp 1676037725
transform 1 0 187772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2041
timestamp 1676037725
transform 1 0 188876 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2045
timestamp 1676037725
transform 1 0 189244 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2057
timestamp 1676037725
transform 1 0 190348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2069
timestamp 1676037725
transform 1 0 191452 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2073
timestamp 1676037725
transform 1 0 191820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2085
timestamp 1676037725
transform 1 0 192924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2097
timestamp 1676037725
transform 1 0 194028 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2101
timestamp 1676037725
transform 1 0 194396 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2113
timestamp 1676037725
transform 1 0 195500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2125
timestamp 1676037725
transform 1 0 196604 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2129
timestamp 1676037725
transform 1 0 196972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2141
timestamp 1676037725
transform 1 0 198076 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2153
timestamp 1676037725
transform 1 0 199180 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2157
timestamp 1676037725
transform 1 0 199548 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2169
timestamp 1676037725
transform 1 0 200652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2181
timestamp 1676037725
transform 1 0 201756 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2185
timestamp 1676037725
transform 1 0 202124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2197
timestamp 1676037725
transform 1 0 203228 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2209
timestamp 1676037725
transform 1 0 204332 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2213
timestamp 1676037725
transform 1 0 204700 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2225
timestamp 1676037725
transform 1 0 205804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2237
timestamp 1676037725
transform 1 0 206908 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2241
timestamp 1676037725
transform 1 0 207276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2253
timestamp 1676037725
transform 1 0 208380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2265
timestamp 1676037725
transform 1 0 209484 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2269
timestamp 1676037725
transform 1 0 209852 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2281
timestamp 1676037725
transform 1 0 210956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2293
timestamp 1676037725
transform 1 0 212060 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2297
timestamp 1676037725
transform 1 0 212428 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2309
timestamp 1676037725
transform 1 0 213532 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2321
timestamp 1676037725
transform 1 0 214636 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2325
timestamp 1676037725
transform 1 0 215004 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2337
timestamp 1676037725
transform 1 0 216108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2349
timestamp 1676037725
transform 1 0 217212 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2353
timestamp 1676037725
transform 1 0 217580 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2365
timestamp 1676037725
transform 1 0 218684 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2377
timestamp 1676037725
transform 1 0 219788 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2381
timestamp 1676037725
transform 1 0 220156 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2393
timestamp 1676037725
transform 1 0 221260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2405
timestamp 1676037725
transform 1 0 222364 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2409
timestamp 1676037725
transform 1 0 222732 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2421
timestamp 1676037725
transform 1 0 223836 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2433
timestamp 1676037725
transform 1 0 224940 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2437
timestamp 1676037725
transform 1 0 225308 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2449
timestamp 1676037725
transform 1 0 226412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2461
timestamp 1676037725
transform 1 0 227516 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2465
timestamp 1676037725
transform 1 0 227884 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2477
timestamp 1676037725
transform 1 0 228988 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2489
timestamp 1676037725
transform 1 0 230092 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2493
timestamp 1676037725
transform 1 0 230460 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2505
timestamp 1676037725
transform 1 0 231564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2517
timestamp 1676037725
transform 1 0 232668 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2521
timestamp 1676037725
transform 1 0 233036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2533
timestamp 1676037725
transform 1 0 234140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2545
timestamp 1676037725
transform 1 0 235244 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2549
timestamp 1676037725
transform 1 0 235612 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2561
timestamp 1676037725
transform 1 0 236716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2573
timestamp 1676037725
transform 1 0 237820 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2577
timestamp 1676037725
transform 1 0 238188 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2589
timestamp 1676037725
transform 1 0 239292 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2601
timestamp 1676037725
transform 1 0 240396 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2605
timestamp 1676037725
transform 1 0 240764 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2617
timestamp 1676037725
transform 1 0 241868 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2629
timestamp 1676037725
transform 1 0 242972 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2633
timestamp 1676037725
transform 1 0 243340 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2645
timestamp 1676037725
transform 1 0 244444 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2657
timestamp 1676037725
transform 1 0 245548 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2661
timestamp 1676037725
transform 1 0 245916 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2673
timestamp 1676037725
transform 1 0 247020 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2685
timestamp 1676037725
transform 1 0 248124 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2689
timestamp 1676037725
transform 1 0 248492 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2701
timestamp 1676037725
transform 1 0 249596 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2713
timestamp 1676037725
transform 1 0 250700 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2717
timestamp 1676037725
transform 1 0 251068 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2729
timestamp 1676037725
transform 1 0 252172 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2741
timestamp 1676037725
transform 1 0 253276 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2745
timestamp 1676037725
transform 1 0 253644 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2757
timestamp 1676037725
transform 1 0 254748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2769
timestamp 1676037725
transform 1 0 255852 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2773
timestamp 1676037725
transform 1 0 256220 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2785
timestamp 1676037725
transform 1 0 257324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2797
timestamp 1676037725
transform 1 0 258428 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2801
timestamp 1676037725
transform 1 0 258796 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2813
timestamp 1676037725
transform 1 0 259900 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2825
timestamp 1676037725
transform 1 0 261004 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2829
timestamp 1676037725
transform 1 0 261372 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2841
timestamp 1676037725
transform 1 0 262476 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2853
timestamp 1676037725
transform 1 0 263580 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2857
timestamp 1676037725
transform 1 0 263948 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2869
timestamp 1676037725
transform 1 0 265052 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2881
timestamp 1676037725
transform 1 0 266156 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2885
timestamp 1676037725
transform 1 0 266524 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2897
timestamp 1676037725
transform 1 0 267628 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2909
timestamp 1676037725
transform 1 0 268732 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2913
timestamp 1676037725
transform 1 0 269100 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2925
timestamp 1676037725
transform 1 0 270204 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2937
timestamp 1676037725
transform 1 0 271308 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2941
timestamp 1676037725
transform 1 0 271676 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2953
timestamp 1676037725
transform 1 0 272780 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2965
timestamp 1676037725
transform 1 0 273884 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2969
timestamp 1676037725
transform 1 0 274252 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2981
timestamp 1676037725
transform 1 0 275356 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2993
timestamp 1676037725
transform 1 0 276460 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2997
timestamp 1676037725
transform 1 0 276828 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3009
timestamp 1676037725
transform 1 0 277932 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3021
timestamp 1676037725
transform 1 0 279036 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3025
timestamp 1676037725
transform 1 0 279404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3037
timestamp 1676037725
transform 1 0 280508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3049
timestamp 1676037725
transform 1 0 281612 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3053
timestamp 1676037725
transform 1 0 281980 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3065
timestamp 1676037725
transform 1 0 283084 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3077
timestamp 1676037725
transform 1 0 284188 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3081
timestamp 1676037725
transform 1 0 284556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3093
timestamp 1676037725
transform 1 0 285660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3105
timestamp 1676037725
transform 1 0 286764 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3109
timestamp 1676037725
transform 1 0 287132 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3121
timestamp 1676037725
transform 1 0 288236 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3133
timestamp 1676037725
transform 1 0 289340 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3137
timestamp 1676037725
transform 1 0 289708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3149
timestamp 1676037725
transform 1 0 290812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3161
timestamp 1676037725
transform 1 0 291916 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3165
timestamp 1676037725
transform 1 0 292284 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3177
timestamp 1676037725
transform 1 0 293388 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3189
timestamp 1676037725
transform 1 0 294492 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3193
timestamp 1676037725
transform 1 0 294860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3205
timestamp 1676037725
transform 1 0 295964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3217
timestamp 1676037725
transform 1 0 297068 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3221
timestamp 1676037725
transform 1 0 297436 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3233
timestamp 1676037725
transform 1 0 298540 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3245
timestamp 1676037725
transform 1 0 299644 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3249
timestamp 1676037725
transform 1 0 300012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3261
timestamp 1676037725
transform 1 0 301116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3273
timestamp 1676037725
transform 1 0 302220 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3277
timestamp 1676037725
transform 1 0 302588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3289
timestamp 1676037725
transform 1 0 303692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3301
timestamp 1676037725
transform 1 0 304796 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3305
timestamp 1676037725
transform 1 0 305164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3317
timestamp 1676037725
transform 1 0 306268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3329
timestamp 1676037725
transform 1 0 307372 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3333
timestamp 1676037725
transform 1 0 307740 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3345
timestamp 1676037725
transform 1 0 308844 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3357
timestamp 1676037725
transform 1 0 309948 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3361
timestamp 1676037725
transform 1 0 310316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3373
timestamp 1676037725
transform 1 0 311420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3385
timestamp 1676037725
transform 1 0 312524 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3389
timestamp 1676037725
transform 1 0 312892 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3401
timestamp 1676037725
transform 1 0 313996 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3413
timestamp 1676037725
transform 1 0 315100 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3417
timestamp 1676037725
transform 1 0 315468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3429
timestamp 1676037725
transform 1 0 316572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3441
timestamp 1676037725
transform 1 0 317676 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3445
timestamp 1676037725
transform 1 0 318044 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3457
timestamp 1676037725
transform 1 0 319148 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3469
timestamp 1676037725
transform 1 0 320252 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3473
timestamp 1676037725
transform 1 0 320620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3485
timestamp 1676037725
transform 1 0 321724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3497
timestamp 1676037725
transform 1 0 322828 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3501
timestamp 1676037725
transform 1 0 323196 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3513
timestamp 1676037725
transform 1 0 324300 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3525
timestamp 1676037725
transform 1 0 325404 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3529
timestamp 1676037725
transform 1 0 325772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3541
timestamp 1676037725
transform 1 0 326876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3553
timestamp 1676037725
transform 1 0 327980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3557
timestamp 1676037725
transform 1 0 328348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3569
timestamp 1676037725
transform 1 0 329452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3581
timestamp 1676037725
transform 1 0 330556 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3585
timestamp 1676037725
transform 1 0 330924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3597
timestamp 1676037725
transform 1 0 332028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3609
timestamp 1676037725
transform 1 0 333132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3613
timestamp 1676037725
transform 1 0 333500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3625
timestamp 1676037725
transform 1 0 334604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3637
timestamp 1676037725
transform 1 0 335708 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3641
timestamp 1676037725
transform 1 0 336076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3653
timestamp 1676037725
transform 1 0 337180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3665
timestamp 1676037725
transform 1 0 338284 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3669
timestamp 1676037725
transform 1 0 338652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3681
timestamp 1676037725
transform 1 0 339756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3693
timestamp 1676037725
transform 1 0 340860 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3697
timestamp 1676037725
transform 1 0 341228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3709
timestamp 1676037725
transform 1 0 342332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3721
timestamp 1676037725
transform 1 0 343436 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3725
timestamp 1676037725
transform 1 0 343804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3737
timestamp 1676037725
transform 1 0 344908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3749
timestamp 1676037725
transform 1 0 346012 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3753
timestamp 1676037725
transform 1 0 346380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3765
timestamp 1676037725
transform 1 0 347484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3777
timestamp 1676037725
transform 1 0 348588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3781
timestamp 1676037725
transform 1 0 348956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3793
timestamp 1676037725
transform 1 0 350060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3805
timestamp 1676037725
transform 1 0 351164 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3809
timestamp 1676037725
transform 1 0 351532 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3821
timestamp 1676037725
transform 1 0 352636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3833
timestamp 1676037725
transform 1 0 353740 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3837
timestamp 1676037725
transform 1 0 354108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3849
timestamp 1676037725
transform 1 0 355212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3861
timestamp 1676037725
transform 1 0 356316 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3865
timestamp 1676037725
transform 1 0 356684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3877
timestamp 1676037725
transform 1 0 357788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3889
timestamp 1676037725
transform 1 0 358892 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3893
timestamp 1676037725
transform 1 0 359260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3905
timestamp 1676037725
transform 1 0 360364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3917
timestamp 1676037725
transform 1 0 361468 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3921
timestamp 1676037725
transform 1 0 361836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3933
timestamp 1676037725
transform 1 0 362940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3945
timestamp 1676037725
transform 1 0 364044 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3949
timestamp 1676037725
transform 1 0 364412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3961
timestamp 1676037725
transform 1 0 365516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3973
timestamp 1676037725
transform 1 0 366620 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3977
timestamp 1676037725
transform 1 0 366988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3989
timestamp 1676037725
transform 1 0 368092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4001
timestamp 1676037725
transform 1 0 369196 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4005
timestamp 1676037725
transform 1 0 369564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4017
timestamp 1676037725
transform 1 0 370668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4029
timestamp 1676037725
transform 1 0 371772 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4033
timestamp 1676037725
transform 1 0 372140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4045
timestamp 1676037725
transform 1 0 373244 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4057
timestamp 1676037725
transform 1 0 374348 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4061
timestamp 1676037725
transform 1 0 374716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4073
timestamp 1676037725
transform 1 0 375820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4085
timestamp 1676037725
transform 1 0 376924 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4089
timestamp 1676037725
transform 1 0 377292 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4101
timestamp 1676037725
transform 1 0 378396 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4113
timestamp 1676037725
transform 1 0 379500 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4117
timestamp 1676037725
transform 1 0 379868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4129
timestamp 1676037725
transform 1 0 380972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4141
timestamp 1676037725
transform 1 0 382076 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4145
timestamp 1676037725
transform 1 0 382444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4157
timestamp 1676037725
transform 1 0 383548 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4169
timestamp 1676037725
transform 1 0 384652 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4173
timestamp 1676037725
transform 1 0 385020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4185
timestamp 1676037725
transform 1 0 386124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4197
timestamp 1676037725
transform 1 0 387228 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4201
timestamp 1676037725
transform 1 0 387596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4213
timestamp 1676037725
transform 1 0 388700 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4225
timestamp 1676037725
transform 1 0 389804 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4229
timestamp 1676037725
transform 1 0 390172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4241
timestamp 1676037725
transform 1 0 391276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4253
timestamp 1676037725
transform 1 0 392380 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4257
timestamp 1676037725
transform 1 0 392748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4269
timestamp 1676037725
transform 1 0 393852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4281
timestamp 1676037725
transform 1 0 394956 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4285
timestamp 1676037725
transform 1 0 395324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4297
timestamp 1676037725
transform 1 0 396428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4309
timestamp 1676037725
transform 1 0 397532 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4313
timestamp 1676037725
transform 1 0 397900 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4325
timestamp 1676037725
transform 1 0 399004 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4337
timestamp 1676037725
transform 1 0 400108 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4341
timestamp 1676037725
transform 1 0 400476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4353
timestamp 1676037725
transform 1 0 401580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4365
timestamp 1676037725
transform 1 0 402684 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4369
timestamp 1676037725
transform 1 0 403052 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4381
timestamp 1676037725
transform 1 0 404156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4393
timestamp 1676037725
transform 1 0 405260 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4397
timestamp 1676037725
transform 1 0 405628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4409
timestamp 1676037725
transform 1 0 406732 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4421
timestamp 1676037725
transform 1 0 407836 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4425
timestamp 1676037725
transform 1 0 408204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4437
timestamp 1676037725
transform 1 0 409308 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4449
timestamp 1676037725
transform 1 0 410412 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4453
timestamp 1676037725
transform 1 0 410780 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4465
timestamp 1676037725
transform 1 0 411884 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4477
timestamp 1676037725
transform 1 0 412988 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4481
timestamp 1676037725
transform 1 0 413356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4493
timestamp 1676037725
transform 1 0 414460 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4505
timestamp 1676037725
transform 1 0 415564 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4509
timestamp 1676037725
transform 1 0 415932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4521
timestamp 1676037725
transform 1 0 417036 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4533
timestamp 1676037725
transform 1 0 418140 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4537
timestamp 1676037725
transform 1 0 418508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4549
timestamp 1676037725
transform 1 0 419612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4561
timestamp 1676037725
transform 1 0 420716 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4565
timestamp 1676037725
transform 1 0 421084 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4577
timestamp 1676037725
transform 1 0 422188 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4589
timestamp 1676037725
transform 1 0 423292 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4593
timestamp 1676037725
transform 1 0 423660 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4605
timestamp 1676037725
transform 1 0 424764 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4617
timestamp 1676037725
transform 1 0 425868 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4621
timestamp 1676037725
transform 1 0 426236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4633
timestamp 1676037725
transform 1 0 427340 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4645
timestamp 1676037725
transform 1 0 428444 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4649
timestamp 1676037725
transform 1 0 428812 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4661
timestamp 1676037725
transform 1 0 429916 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4673
timestamp 1676037725
transform 1 0 431020 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4677
timestamp 1676037725
transform 1 0 431388 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4689
timestamp 1676037725
transform 1 0 432492 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4701
timestamp 1676037725
transform 1 0 433596 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4705
timestamp 1676037725
transform 1 0 433964 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4717
timestamp 1676037725
transform 1 0 435068 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4729
timestamp 1676037725
transform 1 0 436172 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4733
timestamp 1676037725
transform 1 0 436540 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4745
timestamp 1676037725
transform 1 0 437644 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4757
timestamp 1676037725
transform 1 0 438748 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4761
timestamp 1676037725
transform 1 0 439116 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4773
timestamp 1676037725
transform 1 0 440220 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4785
timestamp 1676037725
transform 1 0 441324 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4789
timestamp 1676037725
transform 1 0 441692 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4801
timestamp 1676037725
transform 1 0 442796 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4813
timestamp 1676037725
transform 1 0 443900 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4817
timestamp 1676037725
transform 1 0 444268 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4829
timestamp 1676037725
transform 1 0 445372 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4841
timestamp 1676037725
transform 1 0 446476 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4845
timestamp 1676037725
transform 1 0 446844 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4857
timestamp 1676037725
transform 1 0 447948 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4869
timestamp 1676037725
transform 1 0 449052 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4873
timestamp 1676037725
transform 1 0 449420 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4885
timestamp 1676037725
transform 1 0 450524 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4897
timestamp 1676037725
transform 1 0 451628 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4901
timestamp 1676037725
transform 1 0 451996 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4913
timestamp 1676037725
transform 1 0 453100 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4925
timestamp 1676037725
transform 1 0 454204 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4929
timestamp 1676037725
transform 1 0 454572 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4941
timestamp 1676037725
transform 1 0 455676 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4953
timestamp 1676037725
transform 1 0 456780 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4957
timestamp 1676037725
transform 1 0 457148 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4969
timestamp 1676037725
transform 1 0 458252 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4981
timestamp 1676037725
transform 1 0 459356 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4985
timestamp 1676037725
transform 1 0 459724 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4997
timestamp 1676037725
transform 1 0 460828 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5009
timestamp 1676037725
transform 1 0 461932 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5013
timestamp 1676037725
transform 1 0 462300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5025
timestamp 1676037725
transform 1 0 463404 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5037
timestamp 1676037725
transform 1 0 464508 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5041
timestamp 1676037725
transform 1 0 464876 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5053
timestamp 1676037725
transform 1 0 465980 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5065
timestamp 1676037725
transform 1 0 467084 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5069
timestamp 1676037725
transform 1 0 467452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5081
timestamp 1676037725
transform 1 0 468556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5093
timestamp 1676037725
transform 1 0 469660 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5097
timestamp 1676037725
transform 1 0 470028 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5109
timestamp 1676037725
transform 1 0 471132 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5121
timestamp 1676037725
transform 1 0 472236 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5125
timestamp 1676037725
transform 1 0 472604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5137
timestamp 1676037725
transform 1 0 473708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5149
timestamp 1676037725
transform 1 0 474812 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5153
timestamp 1676037725
transform 1 0 475180 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5165
timestamp 1676037725
transform 1 0 476284 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5177
timestamp 1676037725
transform 1 0 477388 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5181
timestamp 1676037725
transform 1 0 477756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5193
timestamp 1676037725
transform 1 0 478860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5205
timestamp 1676037725
transform 1 0 479964 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5209
timestamp 1676037725
transform 1 0 480332 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5221
timestamp 1676037725
transform 1 0 481436 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5233
timestamp 1676037725
transform 1 0 482540 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5237
timestamp 1676037725
transform 1 0 482908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5249
timestamp 1676037725
transform 1 0 484012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5261
timestamp 1676037725
transform 1 0 485116 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5265
timestamp 1676037725
transform 1 0 485484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5277
timestamp 1676037725
transform 1 0 486588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5289
timestamp 1676037725
transform 1 0 487692 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5293
timestamp 1676037725
transform 1 0 488060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5305
timestamp 1676037725
transform 1 0 489164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5317
timestamp 1676037725
transform 1 0 490268 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5321
timestamp 1676037725
transform 1 0 490636 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5333
timestamp 1676037725
transform 1 0 491740 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5345
timestamp 1676037725
transform 1 0 492844 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5349
timestamp 1676037725
transform 1 0 493212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5361
timestamp 1676037725
transform 1 0 494316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5373
timestamp 1676037725
transform 1 0 495420 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5377
timestamp 1676037725
transform 1 0 495788 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5389
timestamp 1676037725
transform 1 0 496892 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5401
timestamp 1676037725
transform 1 0 497996 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5405
timestamp 1676037725
transform 1 0 498364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5417
timestamp 1676037725
transform 1 0 499468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5429
timestamp 1676037725
transform 1 0 500572 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5433
timestamp 1676037725
transform 1 0 500940 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5445
timestamp 1676037725
transform 1 0 502044 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5457
timestamp 1676037725
transform 1 0 503148 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5461
timestamp 1676037725
transform 1 0 503516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5473
timestamp 1676037725
transform 1 0 504620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5485
timestamp 1676037725
transform 1 0 505724 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5489
timestamp 1676037725
transform 1 0 506092 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5501
timestamp 1676037725
transform 1 0 507196 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5513
timestamp 1676037725
transform 1 0 508300 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5517
timestamp 1676037725
transform 1 0 508668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5529
timestamp 1676037725
transform 1 0 509772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5541
timestamp 1676037725
transform 1 0 510876 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5545
timestamp 1676037725
transform 1 0 511244 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5557
timestamp 1676037725
transform 1 0 512348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5569
timestamp 1676037725
transform 1 0 513452 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5573
timestamp 1676037725
transform 1 0 513820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5585
timestamp 1676037725
transform 1 0 514924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5597
timestamp 1676037725
transform 1 0 516028 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5601
timestamp 1676037725
transform 1 0 516396 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5613
timestamp 1676037725
transform 1 0 517500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5625
timestamp 1676037725
transform 1 0 518604 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5629
timestamp 1676037725
transform 1 0 518972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5641
timestamp 1676037725
transform 1 0 520076 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5653
timestamp 1676037725
transform 1 0 521180 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5657
timestamp 1676037725
transform 1 0 521548 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5669
timestamp 1676037725
transform 1 0 522652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5681
timestamp 1676037725
transform 1 0 523756 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5685
timestamp 1676037725
transform 1 0 524124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5697
timestamp 1676037725
transform 1 0 525228 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5709
timestamp 1676037725
transform 1 0 526332 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5713
timestamp 1676037725
transform 1 0 526700 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_5725
timestamp 1676037725
transform 1 0 527804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 528816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 528816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 528816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 528816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 528816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 528816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 528816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 528816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 528816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 528816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1676037725
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1676037725
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1676037725
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1676037725
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1676037725
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1676037725
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1676037725
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1676037725
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1676037725
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1676037725
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1676037725
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1676037725
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1676037725
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1676037725
transform 1 0 83536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1676037725
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1676037725
transform 1 0 88688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1676037725
transform 1 0 91264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1676037725
transform 1 0 93840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1676037725
transform 1 0 96416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1676037725
transform 1 0 98992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1676037725
transform 1 0 101568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1676037725
transform 1 0 104144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1676037725
transform 1 0 106720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1676037725
transform 1 0 109296 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1676037725
transform 1 0 111872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1676037725
transform 1 0 114448 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1676037725
transform 1 0 117024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1676037725
transform 1 0 119600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1676037725
transform 1 0 122176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1676037725
transform 1 0 124752 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1676037725
transform 1 0 127328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1676037725
transform 1 0 129904 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1676037725
transform 1 0 132480 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1676037725
transform 1 0 135056 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1676037725
transform 1 0 137632 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 140208 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 142784 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 145360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 147936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 150512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 153088 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 155664 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 158240 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 160816 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 163392 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 165968 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 168544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 171120 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 173696 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 176272 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 178848 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 181424 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 184000 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 186576 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 189152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 191728 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 194304 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 196880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 199456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 202032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 204608 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 207184 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 209760 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 212336 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 214912 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 217488 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 220064 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 222640 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 225216 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 227792 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 230368 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 232944 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 235520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 238096 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 240672 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 243248 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 245824 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 248400 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 250976 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 253552 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 256128 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 258704 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 261280 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 263856 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 266432 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 269008 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 271584 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 274160 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 276736 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 279312 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 281888 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 284464 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 287040 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 289616 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 292192 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 294768 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 297344 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 299920 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 302496 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 305072 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 307648 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 310224 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 312800 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 315376 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 317952 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 320528 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 323104 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 325680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 328256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 330832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 333408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 335984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 338560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 341136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 343712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 346288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 348864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 351440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 354016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 356592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 359168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 361744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 364320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 366896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 369472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 372048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 374624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 377200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 379776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 382352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 384928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 387504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 390080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 392656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 395232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 397808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 400384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 402960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 405536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 408112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 410688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 413264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 415840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 418416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 420992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 423568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 426144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 428720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 431296 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 433872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 436448 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 439024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 441600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 444176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 446752 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 449328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 451904 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 454480 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 457056 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 459632 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 462208 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 464784 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 467360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 469936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 472512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 475088 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 477664 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 480240 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 482816 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 485392 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 487968 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 490544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 493120 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 495696 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 498272 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 500848 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 503424 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 506000 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 508576 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 511152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 513728 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 516304 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 518880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 521456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 524032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 526608 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 88688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 93840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 98992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 104144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 109296 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 114448 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 119600 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 124752 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 129904 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 135056 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 140208 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 145360 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 150512 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 155664 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 160816 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 165968 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 171120 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 176272 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 181424 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 186576 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 191728 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 196880 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 202032 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 207184 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 212336 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 217488 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 222640 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 227792 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 232944 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 238096 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 243248 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 248400 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 253552 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 258704 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 263856 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 269008 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 274160 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 279312 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 284464 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 289616 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 294768 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 299920 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 305072 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 310224 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 315376 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 320528 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 325680 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 330832 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 335984 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 341136 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 346288 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 351440 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 356592 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 361744 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 366896 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 372048 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 377200 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 382352 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 387504 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 392656 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 397808 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 402960 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 408112 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 413264 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 418416 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 423568 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 428720 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 433872 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 439024 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 444176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 449328 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 454480 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 459632 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 464784 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 469936 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 475088 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 480240 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 485392 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 490544 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 495696 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 500848 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 506000 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 511152 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 516304 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 521456 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 526608 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 91264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 96416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 101568 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 106720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 111872 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 117024 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 122176 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 127328 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 132480 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 137632 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 142784 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 147936 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 153088 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 158240 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 163392 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 168544 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 173696 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 178848 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 184000 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 189152 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 194304 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 199456 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 204608 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 209760 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 214912 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 220064 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 225216 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 230368 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 235520 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 240672 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 245824 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 250976 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 256128 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 261280 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 266432 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 271584 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 276736 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 281888 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 287040 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 292192 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 297344 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 302496 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 307648 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 312800 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 317952 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 323104 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 328256 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 333408 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 338560 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 343712 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 348864 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 354016 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 359168 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 364320 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 369472 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 374624 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 379776 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 384928 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 390080 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 395232 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 400384 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 405536 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 410688 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 415840 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 420992 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 426144 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 431296 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 436448 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 441600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 446752 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 451904 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 457056 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 462208 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 467360 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 472512 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 477664 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 482816 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 487968 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 493120 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 498272 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 503424 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 508576 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 513728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 518880 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 524032 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 88688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 93840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 98992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 104144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 109296 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 114448 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 119600 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 124752 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 129904 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 135056 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 140208 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 145360 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 150512 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 155664 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 160816 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 165968 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 171120 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 176272 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 181424 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 186576 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 191728 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 196880 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 202032 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 207184 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 212336 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 217488 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 222640 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 227792 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 232944 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 238096 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 243248 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 248400 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 253552 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 258704 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 263856 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 269008 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 274160 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 279312 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 284464 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 289616 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 294768 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 299920 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 305072 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 310224 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 315376 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 320528 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 325680 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 330832 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 335984 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 341136 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 346288 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 351440 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 356592 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 361744 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 366896 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 372048 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 377200 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 382352 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 387504 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 392656 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 397808 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 402960 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 408112 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 413264 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 418416 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 423568 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 428720 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 433872 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 439024 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 444176 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 449328 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 454480 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 459632 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 464784 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 469936 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 475088 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 480240 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 485392 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 490544 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 495696 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 500848 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 506000 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 511152 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 516304 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 521456 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 526608 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 91264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 96416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 101568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 106720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 111872 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 117024 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 122176 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 127328 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 132480 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 137632 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 142784 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 147936 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 153088 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 158240 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 163392 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 168544 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 173696 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 178848 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 184000 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 189152 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 194304 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 199456 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 204608 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 209760 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 214912 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 220064 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 225216 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 230368 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 235520 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 240672 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 245824 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 250976 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 256128 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 261280 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 266432 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 271584 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 276736 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 281888 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 287040 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 292192 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 297344 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 302496 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 307648 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 312800 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 317952 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 323104 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 328256 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 333408 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 338560 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 343712 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 348864 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 354016 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 359168 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 364320 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 369472 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 374624 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 379776 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 384928 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 390080 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 395232 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 400384 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 405536 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 410688 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 415840 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 420992 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 426144 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 431296 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 436448 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 441600 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 446752 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 451904 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 457056 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 462208 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 467360 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 472512 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 477664 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 482816 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 487968 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 493120 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 498272 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 503424 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 508576 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 513728 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 518880 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 524032 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1676037725
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1676037725
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1676037725
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1676037725
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1676037725
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1676037725
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1676037725
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1676037725
transform 1 0 88688 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1676037725
transform 1 0 93840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1676037725
transform 1 0 98992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1676037725
transform 1 0 104144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1676037725
transform 1 0 109296 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1676037725
transform 1 0 114448 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1676037725
transform 1 0 119600 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1676037725
transform 1 0 124752 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1676037725
transform 1 0 129904 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1676037725
transform 1 0 135056 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1676037725
transform 1 0 140208 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1676037725
transform 1 0 145360 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1676037725
transform 1 0 150512 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1676037725
transform 1 0 155664 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1676037725
transform 1 0 160816 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1676037725
transform 1 0 165968 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1676037725
transform 1 0 171120 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1676037725
transform 1 0 176272 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1676037725
transform 1 0 181424 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1676037725
transform 1 0 186576 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1676037725
transform 1 0 191728 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1676037725
transform 1 0 196880 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1676037725
transform 1 0 202032 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1676037725
transform 1 0 207184 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1676037725
transform 1 0 212336 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1676037725
transform 1 0 217488 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1676037725
transform 1 0 222640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1676037725
transform 1 0 227792 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1676037725
transform 1 0 232944 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1676037725
transform 1 0 238096 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1676037725
transform 1 0 243248 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1676037725
transform 1 0 248400 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1676037725
transform 1 0 253552 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1676037725
transform 1 0 258704 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1676037725
transform 1 0 263856 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1676037725
transform 1 0 269008 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1676037725
transform 1 0 274160 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1676037725
transform 1 0 279312 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1676037725
transform 1 0 284464 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1676037725
transform 1 0 289616 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1676037725
transform 1 0 294768 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1676037725
transform 1 0 299920 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1676037725
transform 1 0 305072 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1676037725
transform 1 0 310224 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1676037725
transform 1 0 315376 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1676037725
transform 1 0 320528 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1676037725
transform 1 0 325680 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1676037725
transform 1 0 330832 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1676037725
transform 1 0 335984 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1676037725
transform 1 0 341136 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1676037725
transform 1 0 346288 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1676037725
transform 1 0 351440 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1676037725
transform 1 0 356592 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1676037725
transform 1 0 361744 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1676037725
transform 1 0 366896 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1676037725
transform 1 0 372048 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1676037725
transform 1 0 377200 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1676037725
transform 1 0 382352 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1676037725
transform 1 0 387504 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1676037725
transform 1 0 392656 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1676037725
transform 1 0 397808 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1676037725
transform 1 0 402960 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1676037725
transform 1 0 408112 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1676037725
transform 1 0 413264 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1676037725
transform 1 0 418416 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1676037725
transform 1 0 423568 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1676037725
transform 1 0 428720 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1676037725
transform 1 0 433872 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1676037725
transform 1 0 439024 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1676037725
transform 1 0 444176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1676037725
transform 1 0 449328 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1676037725
transform 1 0 454480 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1676037725
transform 1 0 459632 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1676037725
transform 1 0 464784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1676037725
transform 1 0 469936 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1676037725
transform 1 0 475088 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1676037725
transform 1 0 480240 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1676037725
transform 1 0 485392 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1676037725
transform 1 0 490544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1676037725
transform 1 0 495696 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1676037725
transform 1 0 500848 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1676037725
transform 1 0 506000 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1676037725
transform 1 0 511152 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1676037725
transform 1 0 516304 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1676037725
transform 1 0 521456 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1676037725
transform 1 0 526608 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1676037725
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1676037725
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1676037725
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1676037725
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1676037725
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1676037725
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1676037725
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1676037725
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1676037725
transform 1 0 91264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1676037725
transform 1 0 96416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1676037725
transform 1 0 101568 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1676037725
transform 1 0 106720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1676037725
transform 1 0 111872 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1676037725
transform 1 0 117024 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1676037725
transform 1 0 122176 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1676037725
transform 1 0 127328 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1676037725
transform 1 0 132480 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1676037725
transform 1 0 137632 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1676037725
transform 1 0 142784 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1676037725
transform 1 0 147936 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1676037725
transform 1 0 153088 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1676037725
transform 1 0 158240 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1676037725
transform 1 0 163392 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1676037725
transform 1 0 168544 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1676037725
transform 1 0 173696 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1676037725
transform 1 0 178848 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1676037725
transform 1 0 184000 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1676037725
transform 1 0 189152 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1676037725
transform 1 0 194304 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1676037725
transform 1 0 199456 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1676037725
transform 1 0 204608 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1676037725
transform 1 0 209760 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1676037725
transform 1 0 214912 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1676037725
transform 1 0 220064 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1676037725
transform 1 0 225216 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1676037725
transform 1 0 230368 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1676037725
transform 1 0 235520 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1676037725
transform 1 0 240672 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1676037725
transform 1 0 245824 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1676037725
transform 1 0 250976 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1676037725
transform 1 0 256128 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1676037725
transform 1 0 261280 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1676037725
transform 1 0 266432 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1676037725
transform 1 0 271584 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1676037725
transform 1 0 276736 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1676037725
transform 1 0 281888 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1676037725
transform 1 0 287040 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1676037725
transform 1 0 292192 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1676037725
transform 1 0 297344 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1676037725
transform 1 0 302496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1676037725
transform 1 0 307648 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1676037725
transform 1 0 312800 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1676037725
transform 1 0 317952 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1676037725
transform 1 0 323104 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1676037725
transform 1 0 328256 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1676037725
transform 1 0 333408 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1676037725
transform 1 0 338560 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1676037725
transform 1 0 343712 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1676037725
transform 1 0 348864 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1676037725
transform 1 0 354016 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1676037725
transform 1 0 359168 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1676037725
transform 1 0 364320 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1676037725
transform 1 0 369472 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1676037725
transform 1 0 374624 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1676037725
transform 1 0 379776 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1676037725
transform 1 0 384928 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1676037725
transform 1 0 390080 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1676037725
transform 1 0 395232 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1676037725
transform 1 0 400384 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1676037725
transform 1 0 405536 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1676037725
transform 1 0 410688 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1676037725
transform 1 0 415840 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1676037725
transform 1 0 420992 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1676037725
transform 1 0 426144 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1676037725
transform 1 0 431296 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1676037725
transform 1 0 436448 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1676037725
transform 1 0 441600 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1676037725
transform 1 0 446752 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1676037725
transform 1 0 451904 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1676037725
transform 1 0 457056 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1676037725
transform 1 0 462208 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1676037725
transform 1 0 467360 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1676037725
transform 1 0 472512 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1676037725
transform 1 0 477664 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1676037725
transform 1 0 482816 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1676037725
transform 1 0 487968 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1676037725
transform 1 0 493120 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1676037725
transform 1 0 498272 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1676037725
transform 1 0 503424 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1676037725
transform 1 0 508576 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1676037725
transform 1 0 513728 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1676037725
transform 1 0 518880 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1676037725
transform 1 0 524032 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1676037725
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1676037725
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1676037725
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1676037725
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1676037725
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1676037725
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1676037725
transform 1 0 83536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1676037725
transform 1 0 88688 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1676037725
transform 1 0 93840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1676037725
transform 1 0 98992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1676037725
transform 1 0 104144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1676037725
transform 1 0 109296 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1676037725
transform 1 0 114448 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1676037725
transform 1 0 119600 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1676037725
transform 1 0 124752 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1676037725
transform 1 0 129904 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1676037725
transform 1 0 135056 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1676037725
transform 1 0 140208 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1676037725
transform 1 0 145360 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1676037725
transform 1 0 150512 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1676037725
transform 1 0 155664 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1676037725
transform 1 0 160816 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1676037725
transform 1 0 165968 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1676037725
transform 1 0 171120 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1676037725
transform 1 0 176272 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1676037725
transform 1 0 181424 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1676037725
transform 1 0 186576 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1676037725
transform 1 0 191728 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1676037725
transform 1 0 196880 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1676037725
transform 1 0 202032 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1676037725
transform 1 0 207184 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1676037725
transform 1 0 212336 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1676037725
transform 1 0 217488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1676037725
transform 1 0 222640 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1676037725
transform 1 0 227792 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1676037725
transform 1 0 232944 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1676037725
transform 1 0 238096 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1676037725
transform 1 0 243248 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1676037725
transform 1 0 248400 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1676037725
transform 1 0 253552 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1676037725
transform 1 0 258704 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1676037725
transform 1 0 263856 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1676037725
transform 1 0 269008 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1676037725
transform 1 0 274160 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1676037725
transform 1 0 279312 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1676037725
transform 1 0 284464 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1676037725
transform 1 0 289616 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1676037725
transform 1 0 294768 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1676037725
transform 1 0 299920 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1676037725
transform 1 0 305072 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1676037725
transform 1 0 310224 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1676037725
transform 1 0 315376 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1676037725
transform 1 0 320528 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1676037725
transform 1 0 325680 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1676037725
transform 1 0 330832 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1676037725
transform 1 0 335984 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1676037725
transform 1 0 341136 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1676037725
transform 1 0 346288 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1676037725
transform 1 0 351440 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1676037725
transform 1 0 356592 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1676037725
transform 1 0 361744 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1676037725
transform 1 0 366896 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1676037725
transform 1 0 372048 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1676037725
transform 1 0 377200 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1676037725
transform 1 0 382352 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1676037725
transform 1 0 387504 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1676037725
transform 1 0 392656 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1676037725
transform 1 0 397808 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1676037725
transform 1 0 402960 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1676037725
transform 1 0 408112 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1676037725
transform 1 0 413264 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1676037725
transform 1 0 418416 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1676037725
transform 1 0 423568 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1676037725
transform 1 0 428720 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1676037725
transform 1 0 433872 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1676037725
transform 1 0 439024 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1676037725
transform 1 0 444176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1676037725
transform 1 0 449328 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1676037725
transform 1 0 454480 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1676037725
transform 1 0 459632 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1676037725
transform 1 0 464784 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1676037725
transform 1 0 469936 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1676037725
transform 1 0 475088 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1676037725
transform 1 0 480240 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1676037725
transform 1 0 485392 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1676037725
transform 1 0 490544 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1676037725
transform 1 0 495696 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1676037725
transform 1 0 500848 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1676037725
transform 1 0 506000 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1676037725
transform 1 0 511152 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1676037725
transform 1 0 516304 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1676037725
transform 1 0 521456 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1676037725
transform 1 0 526608 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1676037725
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1676037725
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1676037725
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1676037725
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1676037725
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1676037725
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1676037725
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1676037725
transform 1 0 86112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1676037725
transform 1 0 91264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1676037725
transform 1 0 96416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1676037725
transform 1 0 101568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1676037725
transform 1 0 106720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1676037725
transform 1 0 111872 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1676037725
transform 1 0 117024 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1676037725
transform 1 0 122176 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1676037725
transform 1 0 127328 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1676037725
transform 1 0 132480 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1676037725
transform 1 0 137632 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1676037725
transform 1 0 142784 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1676037725
transform 1 0 147936 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1676037725
transform 1 0 153088 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1676037725
transform 1 0 158240 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1676037725
transform 1 0 163392 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1676037725
transform 1 0 168544 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1676037725
transform 1 0 173696 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1676037725
transform 1 0 178848 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1676037725
transform 1 0 184000 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1676037725
transform 1 0 189152 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1676037725
transform 1 0 194304 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1676037725
transform 1 0 199456 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1676037725
transform 1 0 204608 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1676037725
transform 1 0 209760 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1676037725
transform 1 0 214912 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1676037725
transform 1 0 220064 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1676037725
transform 1 0 225216 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1676037725
transform 1 0 230368 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1676037725
transform 1 0 235520 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1676037725
transform 1 0 240672 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1676037725
transform 1 0 245824 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1676037725
transform 1 0 250976 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1676037725
transform 1 0 256128 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1676037725
transform 1 0 261280 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1676037725
transform 1 0 266432 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1676037725
transform 1 0 271584 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1676037725
transform 1 0 276736 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1676037725
transform 1 0 281888 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1676037725
transform 1 0 287040 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1676037725
transform 1 0 292192 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1676037725
transform 1 0 297344 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1676037725
transform 1 0 302496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1676037725
transform 1 0 307648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1676037725
transform 1 0 312800 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1676037725
transform 1 0 317952 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1676037725
transform 1 0 323104 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1676037725
transform 1 0 328256 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1676037725
transform 1 0 333408 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1676037725
transform 1 0 338560 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1676037725
transform 1 0 343712 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1676037725
transform 1 0 348864 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1676037725
transform 1 0 354016 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1676037725
transform 1 0 359168 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1676037725
transform 1 0 364320 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1676037725
transform 1 0 369472 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1676037725
transform 1 0 374624 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1676037725
transform 1 0 379776 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1676037725
transform 1 0 384928 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1676037725
transform 1 0 390080 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1676037725
transform 1 0 395232 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1676037725
transform 1 0 400384 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1676037725
transform 1 0 405536 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1676037725
transform 1 0 410688 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1676037725
transform 1 0 415840 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1676037725
transform 1 0 420992 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1676037725
transform 1 0 426144 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1676037725
transform 1 0 431296 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1676037725
transform 1 0 436448 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1676037725
transform 1 0 441600 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1676037725
transform 1 0 446752 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1676037725
transform 1 0 451904 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1676037725
transform 1 0 457056 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1676037725
transform 1 0 462208 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1676037725
transform 1 0 467360 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1676037725
transform 1 0 472512 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1676037725
transform 1 0 477664 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1676037725
transform 1 0 482816 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1676037725
transform 1 0 487968 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1676037725
transform 1 0 493120 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1676037725
transform 1 0 498272 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1676037725
transform 1 0 503424 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1676037725
transform 1 0 508576 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1676037725
transform 1 0 513728 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1676037725
transform 1 0 518880 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1676037725
transform 1 0 524032 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1676037725
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1676037725
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1676037725
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1676037725
transform 1 0 19136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1676037725
transform 1 0 24288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1676037725
transform 1 0 29440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1676037725
transform 1 0 34592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1676037725
transform 1 0 39744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1676037725
transform 1 0 44896 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1676037725
transform 1 0 50048 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1676037725
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1676037725
transform 1 0 55200 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1676037725
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1676037725
transform 1 0 60352 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1676037725
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1676037725
transform 1 0 65504 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1676037725
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1676037725
transform 1 0 70656 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1676037725
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1676037725
transform 1 0 75808 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1676037725
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1676037725
transform 1 0 80960 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1676037725
transform 1 0 83536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1676037725
transform 1 0 86112 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1676037725
transform 1 0 88688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1676037725
transform 1 0 91264 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1676037725
transform 1 0 93840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1676037725
transform 1 0 96416 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1676037725
transform 1 0 98992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1676037725
transform 1 0 101568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1676037725
transform 1 0 104144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1676037725
transform 1 0 106720 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1676037725
transform 1 0 109296 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1676037725
transform 1 0 111872 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1676037725
transform 1 0 114448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1676037725
transform 1 0 117024 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1676037725
transform 1 0 119600 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1676037725
transform 1 0 122176 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1676037725
transform 1 0 124752 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1676037725
transform 1 0 127328 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1676037725
transform 1 0 129904 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1676037725
transform 1 0 132480 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1676037725
transform 1 0 135056 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1676037725
transform 1 0 137632 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1676037725
transform 1 0 140208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1676037725
transform 1 0 142784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1676037725
transform 1 0 145360 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1676037725
transform 1 0 147936 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1676037725
transform 1 0 150512 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1676037725
transform 1 0 153088 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1676037725
transform 1 0 155664 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1676037725
transform 1 0 158240 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1676037725
transform 1 0 160816 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1676037725
transform 1 0 163392 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1676037725
transform 1 0 165968 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1676037725
transform 1 0 168544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1676037725
transform 1 0 171120 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1676037725
transform 1 0 173696 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1676037725
transform 1 0 176272 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1676037725
transform 1 0 178848 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1676037725
transform 1 0 181424 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1676037725
transform 1 0 184000 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1676037725
transform 1 0 186576 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1676037725
transform 1 0 189152 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1676037725
transform 1 0 191728 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1676037725
transform 1 0 194304 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1676037725
transform 1 0 196880 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1676037725
transform 1 0 199456 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1676037725
transform 1 0 202032 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1676037725
transform 1 0 204608 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1676037725
transform 1 0 207184 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1676037725
transform 1 0 209760 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1676037725
transform 1 0 212336 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1676037725
transform 1 0 214912 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1676037725
transform 1 0 217488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1676037725
transform 1 0 220064 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1676037725
transform 1 0 222640 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1676037725
transform 1 0 225216 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1676037725
transform 1 0 227792 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1676037725
transform 1 0 230368 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1676037725
transform 1 0 232944 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1676037725
transform 1 0 235520 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1676037725
transform 1 0 238096 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1676037725
transform 1 0 240672 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1676037725
transform 1 0 243248 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1676037725
transform 1 0 245824 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1676037725
transform 1 0 248400 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1676037725
transform 1 0 250976 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1676037725
transform 1 0 253552 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1676037725
transform 1 0 256128 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1676037725
transform 1 0 258704 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1676037725
transform 1 0 261280 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1676037725
transform 1 0 263856 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1676037725
transform 1 0 266432 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1676037725
transform 1 0 269008 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1676037725
transform 1 0 271584 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1676037725
transform 1 0 274160 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1676037725
transform 1 0 276736 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1676037725
transform 1 0 279312 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1676037725
transform 1 0 281888 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1676037725
transform 1 0 284464 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1676037725
transform 1 0 287040 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1676037725
transform 1 0 289616 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1676037725
transform 1 0 292192 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1676037725
transform 1 0 294768 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1676037725
transform 1 0 297344 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1676037725
transform 1 0 299920 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1676037725
transform 1 0 302496 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1676037725
transform 1 0 305072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1676037725
transform 1 0 307648 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1676037725
transform 1 0 310224 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1676037725
transform 1 0 312800 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1676037725
transform 1 0 315376 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1676037725
transform 1 0 317952 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1676037725
transform 1 0 320528 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1676037725
transform 1 0 323104 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1676037725
transform 1 0 325680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1676037725
transform 1 0 328256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1676037725
transform 1 0 330832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1676037725
transform 1 0 333408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1676037725
transform 1 0 335984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1676037725
transform 1 0 338560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1676037725
transform 1 0 341136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1676037725
transform 1 0 343712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1676037725
transform 1 0 346288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1676037725
transform 1 0 348864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1676037725
transform 1 0 351440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1676037725
transform 1 0 354016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1676037725
transform 1 0 356592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1676037725
transform 1 0 359168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1676037725
transform 1 0 361744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1676037725
transform 1 0 364320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1676037725
transform 1 0 366896 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1676037725
transform 1 0 369472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1676037725
transform 1 0 372048 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1676037725
transform 1 0 374624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1676037725
transform 1 0 377200 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1676037725
transform 1 0 379776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1676037725
transform 1 0 382352 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1676037725
transform 1 0 384928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1676037725
transform 1 0 387504 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1676037725
transform 1 0 390080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1676037725
transform 1 0 392656 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1676037725
transform 1 0 395232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1676037725
transform 1 0 397808 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1676037725
transform 1 0 400384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1676037725
transform 1 0 402960 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1676037725
transform 1 0 405536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1676037725
transform 1 0 408112 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1676037725
transform 1 0 410688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1676037725
transform 1 0 413264 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1676037725
transform 1 0 415840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1676037725
transform 1 0 418416 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1676037725
transform 1 0 420992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1676037725
transform 1 0 423568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1676037725
transform 1 0 426144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1676037725
transform 1 0 428720 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1676037725
transform 1 0 431296 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1676037725
transform 1 0 433872 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1676037725
transform 1 0 436448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1676037725
transform 1 0 439024 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1676037725
transform 1 0 441600 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1676037725
transform 1 0 444176 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1676037725
transform 1 0 446752 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1676037725
transform 1 0 449328 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1676037725
transform 1 0 451904 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1676037725
transform 1 0 454480 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1676037725
transform 1 0 457056 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1676037725
transform 1 0 459632 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1676037725
transform 1 0 462208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1676037725
transform 1 0 464784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1676037725
transform 1 0 467360 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1676037725
transform 1 0 469936 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1676037725
transform 1 0 472512 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1676037725
transform 1 0 475088 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1676037725
transform 1 0 477664 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1676037725
transform 1 0 480240 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1676037725
transform 1 0 482816 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1676037725
transform 1 0 485392 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1676037725
transform 1 0 487968 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1676037725
transform 1 0 490544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1676037725
transform 1 0 493120 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1676037725
transform 1 0 495696 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1676037725
transform 1 0 498272 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1676037725
transform 1 0 500848 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1676037725
transform 1 0 503424 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1676037725
transform 1 0 506000 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1676037725
transform 1 0 508576 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1676037725
transform 1 0 511152 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1676037725
transform 1 0 513728 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1676037725
transform 1 0 516304 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1676037725
transform 1 0 518880 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1676037725
transform 1 0 521456 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1676037725
transform 1 0 524032 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1676037725
transform 1 0 526608 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _00_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 331568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _01_
timestamp 1676037725
transform -1 0 329544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _02_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 325128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _03_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 324484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _04_
timestamp 1676037725
transform 1 0 323380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _05_
timestamp 1676037725
transform 1 0 319424 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _06_
timestamp 1676037725
transform 1 0 318780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _07_
timestamp 1676037725
transform 1 0 317124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _08_
timestamp 1676037725
transform 1 0 314548 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _09_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 314824 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _10_
timestamp 1676037725
transform -1 0 312892 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _11_
timestamp 1676037725
transform 1 0 310500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _12_
timestamp 1676037725
transform -1 0 311972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _13_
timestamp 1676037725
transform -1 0 309580 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _14_
timestamp 1676037725
transform 1 0 304520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _15_
timestamp 1676037725
transform -1 0 306820 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _16_
timestamp 1676037725
transform -1 0 303324 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _17_
timestamp 1676037725
transform -1 0 301392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _18_
timestamp 1676037725
transform -1 0 301944 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _19_
timestamp 1676037725
transform -1 0 300748 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _20_
timestamp 1676037725
transform -1 0 297620 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _21_
timestamp 1676037725
transform -1 0 298172 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _22_
timestamp 1676037725
transform -1 0 295964 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1676037725
transform 1 0 357328 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _24_
timestamp 1676037725
transform -1 0 357328 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _25_
timestamp 1676037725
transform -1 0 356132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _26_
timestamp 1676037725
transform 1 0 353740 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _27_
timestamp 1676037725
transform -1 0 354660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _28_
timestamp 1676037725
transform -1 0 352544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _29_
timestamp 1676037725
transform 1 0 350244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _30_
timestamp 1676037725
transform -1 0 349876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _31_
timestamp 1676037725
transform -1 0 348588 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1676037725
transform 1 0 346564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _33_
timestamp 1676037725
transform -1 0 345920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _34_
timestamp 1676037725
transform -1 0 344540 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1676037725
transform 1 0 342148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _36_
timestamp 1676037725
transform -1 0 341780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _37_
timestamp 1676037725
transform -1 0 340308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1676037725
transform 1 0 337824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _39_
timestamp 1676037725
transform -1 0 337456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _40_
timestamp 1676037725
transform -1 0 335616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1676037725
transform 1 0 332304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[0\].u_buf
timestamp 1676037725
transform -1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[1\].u_buf
timestamp 1676037725
transform -1 0 20148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[2\].u_buf
timestamp 1676037725
transform -1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[3\].u_buf
timestamp 1676037725
transform -1 0 56212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[4\].u_buf
timestamp 1676037725
transform -1 0 74244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  u_rp\[5\].u_buf
timestamp 1676037725
transform -1 0 92276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  u_rp\[6\].u_buf
timestamp 1676037725
transform -1 0 110308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[7\].u_buf
timestamp 1676037725
transform -1 0 128340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[8\].u_buf
timestamp 1676037725
transform -1 0 146372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[9\].u_buf
timestamp 1676037725
transform -1 0 164404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[10\].u_buf
timestamp 1676037725
transform -1 0 182436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  u_rp\[11\].u_buf
timestamp 1676037725
transform -1 0 200468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  u_rp\[12\].u_buf
timestamp 1676037725
transform -1 0 218500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[13\].u_buf
timestamp 1676037725
transform -1 0 236532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[14\].u_buf
timestamp 1676037725
transform -1 0 254564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[15\].u_buf
timestamp 1676037725
transform -1 0 272596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[16\].u_buf
timestamp 1676037725
transform -1 0 290628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[17\].u_buf
timestamp 1676037725
transform -1 0 308660 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[18\].u_buf
timestamp 1676037725
transform -1 0 326692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[19\].u_buf
timestamp 1676037725
transform -1 0 344724 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[20\].u_buf
timestamp 1676037725
transform -1 0 362756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[21\].u_buf
timestamp 1676037725
transform -1 0 380788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[22\].u_buf
timestamp 1676037725
transform -1 0 398820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[23\].u_buf
timestamp 1676037725
transform -1 0 416852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[24\].u_buf
timestamp 1676037725
transform -1 0 434884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[25\].u_buf
timestamp 1676037725
transform -1 0 452916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[26\].u_buf
timestamp 1676037725
transform -1 0 470948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  wire1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 394312 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire2
timestamp 1676037725
transform 1 0 300196 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire3
timestamp 1676037725
transform 1 0 205436 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire4
timestamp 1676037725
transform 1 0 391000 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire5
timestamp 1676037725
transform 1 0 296332 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire6
timestamp 1676037725
transform 1 0 202308 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 107364 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire8
timestamp 1676037725
transform 1 0 387780 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire9
timestamp 1676037725
transform 1 0 293112 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire10
timestamp 1676037725
transform 1 0 198444 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire11
timestamp 1676037725
transform 1 0 104420 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire12
timestamp 1676037725
transform 1 0 408388 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire13
timestamp 1676037725
transform 1 0 404524 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire14
timestamp 1676037725
transform 1 0 401028 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire15
timestamp 1676037725
transform 1 0 306636 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire16
timestamp 1676037725
transform 1 0 396796 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire17
timestamp 1676037725
transform 1 0 303324 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire18
timestamp 1676037725
transform 1 0 211508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire19
timestamp 1676037725
transform -1 0 118220 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire20
timestamp 1676037725
transform -1 0 213716 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire21
timestamp 1676037725
transform -1 0 311052 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire22
timestamp 1676037725
transform -1 0 119508 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire23
timestamp 1676037725
transform -1 0 214084 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire24
timestamp 1676037725
transform -1 0 309580 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire25
timestamp 1676037725
transform -1 0 118220 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire26
timestamp 1676037725
transform -1 0 213532 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire27
timestamp 1676037725
transform -1 0 308476 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire28
timestamp 1676037725
transform -1 0 118864 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire29
timestamp 1676037725
transform -1 0 212152 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire30
timestamp 1676037725
transform -1 0 308660 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire31
timestamp 1676037725
transform -1 0 118312 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire32
timestamp 1676037725
transform -1 0 212336 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire33
timestamp 1676037725
transform -1 0 307464 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire34
timestamp 1676037725
transform -1 0 117024 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire35
timestamp 1676037725
transform -1 0 210956 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire36
timestamp 1676037725
transform -1 0 306544 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire37
timestamp 1676037725
transform -1 0 116840 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire38
timestamp 1676037725
transform -1 0 211140 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire39
timestamp 1676037725
transform -1 0 307740 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire40
timestamp 1676037725
transform -1 0 115828 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire41
timestamp 1676037725
transform -1 0 209576 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire42
timestamp 1676037725
transform -1 0 306544 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire43
timestamp 1676037725
transform -1 0 114264 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire44
timestamp 1676037725
transform -1 0 209760 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire45
timestamp 1676037725
transform -1 0 305624 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire46
timestamp 1676037725
transform -1 0 115644 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire47
timestamp 1676037725
transform -1 0 208380 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire48
timestamp 1676037725
transform -1 0 305900 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire49
timestamp 1676037725
transform -1 0 115920 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire50
timestamp 1676037725
transform -1 0 210312 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire51
timestamp 1676037725
transform -1 0 304704 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire52
timestamp 1676037725
transform -1 0 114264 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire53
timestamp 1676037725
transform -1 0 209576 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire54
timestamp 1676037725
transform -1 0 304520 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire55
timestamp 1676037725
transform -1 0 125580 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire56
timestamp 1676037725
transform -1 0 220616 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire57
timestamp 1676037725
transform -1 0 125764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire58
timestamp 1676037725
transform -1 0 219880 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  wire59
timestamp 1676037725
transform 1 0 307464 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  wire60
timestamp 1676037725
transform -1 0 125396 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire61
timestamp 1676037725
transform -1 0 219420 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire62
timestamp 1676037725
transform -1 0 124568 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire63
timestamp 1676037725
transform -1 0 219604 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  wire64
timestamp 1676037725
transform 1 0 308292 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  wire65
timestamp 1676037725
transform -1 0 124568 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire66
timestamp 1676037725
transform -1 0 217304 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire67
timestamp 1676037725
transform -1 0 124476 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire68
timestamp 1676037725
transform -1 0 218408 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire69
timestamp 1676037725
transform -1 0 123372 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire70
timestamp 1676037725
transform -1 0 217304 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire71
timestamp 1676037725
transform -1 0 123372 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire72
timestamp 1676037725
transform -1 0 216108 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire73
timestamp 1676037725
transform -1 0 121992 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire74
timestamp 1676037725
transform -1 0 217212 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire75
timestamp 1676037725
transform -1 0 122176 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire76
timestamp 1676037725
transform -1 0 217212 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire77
timestamp 1676037725
transform -1 0 120796 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire78
timestamp 1676037725
transform -1 0 216108 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire79
timestamp 1676037725
transform -1 0 311972 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire80
timestamp 1676037725
transform -1 0 122084 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire81
timestamp 1676037725
transform -1 0 214728 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire82
timestamp 1676037725
transform -1 0 311236 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire83
timestamp 1676037725
transform -1 0 120980 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire84
timestamp 1676037725
transform -1 0 214912 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire85
timestamp 1676037725
transform -1 0 311052 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire86
timestamp 1676037725
transform -1 0 119416 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire87
timestamp 1676037725
transform -1 0 215648 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire88
timestamp 1676037725
transform -1 0 310316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire89
timestamp 1676037725
transform -1 0 120704 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire90
timestamp 1676037725
transform -1 0 213532 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire91
timestamp 1676037725
transform -1 0 309212 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire92
timestamp 1676037725
transform -1 0 119416 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire93
timestamp 1676037725
transform -1 0 214728 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire94
timestamp 1676037725
transform -1 0 309396 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire95
timestamp 1676037725
transform -1 0 259808 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire96
timestamp 1676037725
transform -1 0 353832 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire97
timestamp 1676037725
transform -1 0 448132 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire98
timestamp 1676037725
transform -1 0 223744 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire99
timestamp 1676037725
transform -1 0 317768 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire100
timestamp 1676037725
transform -1 0 412528 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire101
timestamp 1676037725
transform -1 0 205620 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire102
timestamp 1676037725
transform -1 0 299736 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire103
timestamp 1676037725
transform -1 0 394588 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  wire104 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 170292 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  wire105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 265236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  wire106
timestamp 1676037725
transform -1 0 358616 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire107
timestamp 1676037725
transform -1 0 452916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  wire108
timestamp 1676037725
transform -1 0 152260 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  wire109
timestamp 1676037725
transform -1 0 247204 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  wire110
timestamp 1676037725
transform -1 0 340676 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire111
timestamp 1676037725
transform -1 0 435804 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  wire112
timestamp 1676037725
transform -1 0 492568 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire113
timestamp 1676037725
transform -1 0 474720 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  wire114
timestamp 1676037725
transform -1 0 116196 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  wire115
timestamp 1676037725
transform -1 0 211140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  wire116
timestamp 1676037725
transform -1 0 306176 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire117
timestamp 1676037725
transform -1 0 400016 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire118
timestamp 1676037725
transform -1 0 440128 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire119
timestamp 1676037725
transform -1 0 422096 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire120
timestamp 1676037725
transform -1 0 386032 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire121
timestamp 1676037725
transform -1 0 479320 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire122
timestamp 1676037725
transform -1 0 368000 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire123
timestamp 1676037725
transform -1 0 461380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire124
timestamp 1676037725
transform -1 0 331936 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire125
timestamp 1676037725
transform -1 0 425868 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire126
timestamp 1676037725
transform -1 0 313904 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire127
timestamp 1676037725
transform -1 0 407928 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire128
timestamp 1676037725
transform -1 0 277840 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire129
timestamp 1676037725
transform -1 0 371864 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire130
timestamp 1676037725
transform -1 0 466072 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  wire131
timestamp 1676037725
transform -1 0 98164 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  wire132
timestamp 1676037725
transform -1 0 193108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  wire133
timestamp 1676037725
transform -1 0 286672 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire134
timestamp 1676037725
transform -1 0 381984 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire135
timestamp 1676037725
transform 1 0 251620 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire136
timestamp 1676037725
transform 1 0 157228 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire137
timestamp 1676037725
transform 1 0 63204 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire138
timestamp 1676037725
transform 1 0 256404 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire139
timestamp 1676037725
transform 1 0 161184 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire140
timestamp 1676037725
transform 1 0 66792 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire141
timestamp 1676037725
transform -1 0 389620 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  wire142
timestamp 1676037725
transform -1 0 390724 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire143
timestamp 1676037725
transform 1 0 259348 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire144
timestamp 1676037725
transform 1 0 164956 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire145
timestamp 1676037725
transform 1 0 70932 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire146
timestamp 1676037725
transform 1 0 203228 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire147
timestamp 1676037725
transform 1 0 108284 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  wire148
timestamp 1676037725
transform -1 0 393484 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  wire149
timestamp 1676037725
transform -1 0 396060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire150
timestamp 1676037725
transform 1 0 207460 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire151
timestamp 1676037725
transform 1 0 112240 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  wire152
timestamp 1676037725
transform -1 0 397256 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire153
timestamp 1676037725
transform 1 0 211140 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire154
timestamp 1676037725
transform 1 0 116748 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire155
timestamp 1676037725
transform 1 0 215188 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire156
timestamp 1676037725
transform 1 0 121164 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire157
timestamp 1676037725
transform 1 0 220340 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire158
timestamp 1676037725
transform 1 0 125948 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire159
timestamp 1676037725
transform 1 0 225492 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire160
timestamp 1676037725
transform 1 0 130732 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire161
timestamp 1676037725
transform 1 0 36432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire162
timestamp 1676037725
transform 1 0 231288 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire163
timestamp 1676037725
transform 1 0 136620 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire164
timestamp 1676037725
transform 1 0 42596 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire165
timestamp 1676037725
transform 1 0 238372 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire166
timestamp 1676037725
transform 1 0 143244 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire167
timestamp 1676037725
transform 1 0 48852 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire168
timestamp 1676037725
transform 1 0 243524 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire169
timestamp 1676037725
transform 1 0 148764 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire170
timestamp 1676037725
transform 1 0 54372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire171
timestamp 1676037725
transform 1 0 248676 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire172
timestamp 1676037725
transform 1 0 153364 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire173
timestamp 1676037725
transform 1 0 58696 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire174
timestamp 1676037725
transform 1 0 262844 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire175
timestamp 1676037725
transform 1 0 168544 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire176
timestamp 1676037725
transform 1 0 74612 0 1 2176
box -38 -48 866 592
<< labels >>
flabel metal1 s 20066 0 20122 800 0 FreeSans 224 90 0 0 buf_in[0]
port 0 nsew signal input
flabel metal1 s 408482 0 408538 800 0 FreeSans 224 90 0 0 buf_in[10]
port 1 nsew signal input
flabel metal1 s 408210 0 408266 800 0 FreeSans 224 90 0 0 buf_in[11]
port 2 nsew signal input
flabel metal1 s 23330 0 23386 800 0 FreeSans 224 90 0 0 buf_in[12]
port 3 nsew signal input
flabel metal1 s 407666 0 407722 800 0 FreeSans 224 90 0 0 buf_in[13]
port 4 nsew signal input
flabel metal1 s 407394 0 407450 800 0 FreeSans 224 90 0 0 buf_in[14]
port 5 nsew signal input
flabel metal1 s 24146 0 24202 800 0 FreeSans 224 90 0 0 buf_in[15]
port 6 nsew signal input
flabel metal1 s 406850 0 406906 800 0 FreeSans 224 90 0 0 buf_in[16]
port 7 nsew signal input
flabel metal1 s 406578 0 406634 800 0 FreeSans 224 90 0 0 buf_in[17]
port 8 nsew signal input
flabel metal1 s 24962 0 25018 800 0 FreeSans 224 90 0 0 buf_in[18]
port 9 nsew signal input
flabel metal1 s 406034 0 406090 800 0 FreeSans 224 90 0 0 buf_in[19]
port 10 nsew signal input
flabel metal1 s 410930 0 410986 800 0 FreeSans 224 90 0 0 buf_in[1]
port 11 nsew signal input
flabel metal1 s 405762 0 405818 800 0 FreeSans 224 90 0 0 buf_in[20]
port 12 nsew signal input
flabel metal1 s 25778 0 25834 800 0 FreeSans 224 90 0 0 buf_in[21]
port 13 nsew signal input
flabel metal1 s 405218 0 405274 800 0 FreeSans 224 90 0 0 buf_in[22]
port 14 nsew signal input
flabel metal1 s 404946 0 405002 800 0 FreeSans 224 90 0 0 buf_in[23]
port 15 nsew signal input
flabel metal1 s 26594 0 26650 800 0 FreeSans 224 90 0 0 buf_in[24]
port 16 nsew signal input
flabel metal1 s 404402 0 404458 800 0 FreeSans 224 90 0 0 buf_in[25]
port 17 nsew signal input
flabel metal1 s 404130 0 404186 800 0 FreeSans 224 90 0 0 buf_in[26]
port 18 nsew signal input
flabel metal1 s 27410 0 27466 800 0 FreeSans 224 90 0 0 buf_in[27]
port 19 nsew signal input
flabel metal1 s 403586 0 403642 800 0 FreeSans 224 90 0 0 buf_in[28]
port 20 nsew signal input
flabel metal1 s 403314 0 403370 800 0 FreeSans 224 90 0 0 buf_in[29]
port 21 nsew signal input
flabel metal1 s 410658 0 410714 800 0 FreeSans 224 90 0 0 buf_in[2]
port 22 nsew signal input
flabel metal1 s 28226 0 28282 800 0 FreeSans 224 90 0 0 buf_in[30]
port 23 nsew signal input
flabel metal1 s 402770 0 402826 800 0 FreeSans 224 90 0 0 buf_in[31]
port 24 nsew signal input
flabel metal1 s 402498 0 402554 800 0 FreeSans 224 90 0 0 buf_in[32]
port 25 nsew signal input
flabel metal1 s 29042 0 29098 800 0 FreeSans 224 90 0 0 buf_in[33]
port 26 nsew signal input
flabel metal1 s 401954 0 402010 800 0 FreeSans 224 90 0 0 buf_in[34]
port 27 nsew signal input
flabel metal1 s 401682 0 401738 800 0 FreeSans 224 90 0 0 buf_in[35]
port 28 nsew signal input
flabel metal1 s 29858 0 29914 800 0 FreeSans 224 90 0 0 buf_in[36]
port 29 nsew signal input
flabel metal1 s 401138 0 401194 800 0 FreeSans 224 90 0 0 buf_in[37]
port 30 nsew signal input
flabel metal1 s 400866 0 400922 800 0 FreeSans 224 90 0 0 buf_in[38]
port 31 nsew signal input
flabel metal1 s 30674 0 30730 800 0 FreeSans 224 90 0 0 buf_in[39]
port 32 nsew signal input
flabel metal1 s 20882 0 20938 800 0 FreeSans 224 90 0 0 buf_in[3]
port 33 nsew signal input
flabel metal1 s 400322 0 400378 800 0 FreeSans 224 90 0 0 buf_in[40]
port 34 nsew signal input
flabel metal1 s 400050 0 400106 800 0 FreeSans 224 90 0 0 buf_in[41]
port 35 nsew signal input
flabel metal1 s 410114 0 410170 800 0 FreeSans 224 90 0 0 buf_in[4]
port 36 nsew signal input
flabel metal1 s 409842 0 409898 800 0 FreeSans 224 90 0 0 buf_in[5]
port 37 nsew signal input
flabel metal1 s 21698 0 21754 800 0 FreeSans 224 90 0 0 buf_in[6]
port 38 nsew signal input
flabel metal1 s 409298 0 409354 800 0 FreeSans 224 90 0 0 buf_in[7]
port 39 nsew signal input
flabel metal1 s 409026 0 409082 800 0 FreeSans 224 90 0 0 buf_in[8]
port 40 nsew signal input
flabel metal1 s 22514 0 22570 800 0 FreeSans 224 90 0 0 buf_in[9]
port 41 nsew signal input
flabel metal1 s 411202 0 411258 800 0 FreeSans 224 90 0 0 buf_out[0]
port 42 nsew signal tristate
flabel metal1 s 22786 0 22842 800 0 FreeSans 224 90 0 0 buf_out[10]
port 43 nsew signal tristate
flabel metal1 s 23058 0 23114 800 0 FreeSans 224 90 0 0 buf_out[11]
port 44 nsew signal tristate
flabel metal1 s 407938 0 407994 800 0 FreeSans 224 90 0 0 buf_out[12]
port 45 nsew signal tristate
flabel metal1 s 23602 0 23658 800 0 FreeSans 224 90 0 0 buf_out[13]
port 46 nsew signal tristate
flabel metal1 s 23874 0 23930 800 0 FreeSans 224 90 0 0 buf_out[14]
port 47 nsew signal tristate
flabel metal1 s 407122 0 407178 800 0 FreeSans 224 90 0 0 buf_out[15]
port 48 nsew signal tristate
flabel metal1 s 24418 0 24474 800 0 FreeSans 224 90 0 0 buf_out[16]
port 49 nsew signal tristate
flabel metal1 s 24690 0 24746 800 0 FreeSans 224 90 0 0 buf_out[17]
port 50 nsew signal tristate
flabel metal1 s 406306 0 406362 800 0 FreeSans 224 90 0 0 buf_out[18]
port 51 nsew signal tristate
flabel metal1 s 25234 0 25290 800 0 FreeSans 224 90 0 0 buf_out[19]
port 52 nsew signal tristate
flabel metal1 s 20338 0 20394 800 0 FreeSans 224 90 0 0 buf_out[1]
port 53 nsew signal tristate
flabel metal1 s 25506 0 25562 800 0 FreeSans 224 90 0 0 buf_out[20]
port 54 nsew signal tristate
flabel metal1 s 405490 0 405546 800 0 FreeSans 224 90 0 0 buf_out[21]
port 55 nsew signal tristate
flabel metal1 s 26050 0 26106 800 0 FreeSans 224 90 0 0 buf_out[22]
port 56 nsew signal tristate
flabel metal1 s 26322 0 26378 800 0 FreeSans 224 90 0 0 buf_out[23]
port 57 nsew signal tristate
flabel metal1 s 404674 0 404730 800 0 FreeSans 224 90 0 0 buf_out[24]
port 58 nsew signal tristate
flabel metal1 s 26866 0 26922 800 0 FreeSans 224 90 0 0 buf_out[25]
port 59 nsew signal tristate
flabel metal1 s 27138 0 27194 800 0 FreeSans 224 90 0 0 buf_out[26]
port 60 nsew signal tristate
flabel metal1 s 403858 0 403914 800 0 FreeSans 224 90 0 0 buf_out[27]
port 61 nsew signal tristate
flabel metal1 s 27682 0 27738 800 0 FreeSans 224 90 0 0 buf_out[28]
port 62 nsew signal tristate
flabel metal1 s 27954 0 28010 800 0 FreeSans 224 90 0 0 buf_out[29]
port 63 nsew signal tristate
flabel metal1 s 20610 0 20666 800 0 FreeSans 224 90 0 0 buf_out[2]
port 64 nsew signal tristate
flabel metal1 s 403042 0 403098 800 0 FreeSans 224 90 0 0 buf_out[30]
port 65 nsew signal tristate
flabel metal1 s 28498 0 28554 800 0 FreeSans 224 90 0 0 buf_out[31]
port 66 nsew signal tristate
flabel metal1 s 28770 0 28826 800 0 FreeSans 224 90 0 0 buf_out[32]
port 67 nsew signal tristate
flabel metal1 s 402226 0 402282 800 0 FreeSans 224 90 0 0 buf_out[33]
port 68 nsew signal tristate
flabel metal1 s 29314 0 29370 800 0 FreeSans 224 90 0 0 buf_out[34]
port 69 nsew signal tristate
flabel metal1 s 29586 0 29642 800 0 FreeSans 224 90 0 0 buf_out[35]
port 70 nsew signal tristate
flabel metal1 s 401410 0 401466 800 0 FreeSans 224 90 0 0 buf_out[36]
port 71 nsew signal tristate
flabel metal1 s 30130 0 30186 800 0 FreeSans 224 90 0 0 buf_out[37]
port 72 nsew signal tristate
flabel metal1 s 30402 0 30458 800 0 FreeSans 224 90 0 0 buf_out[38]
port 73 nsew signal tristate
flabel metal1 s 400594 0 400650 800 0 FreeSans 224 90 0 0 buf_out[39]
port 74 nsew signal tristate
flabel metal1 s 410386 0 410442 800 0 FreeSans 224 90 0 0 buf_out[3]
port 75 nsew signal tristate
flabel metal1 s 30946 0 31002 800 0 FreeSans 224 90 0 0 buf_out[40]
port 76 nsew signal tristate
flabel metal1 s 31218 0 31274 800 0 FreeSans 224 90 0 0 buf_out[41]
port 77 nsew signal tristate
flabel metal1 s 21154 0 21210 800 0 FreeSans 224 90 0 0 buf_out[4]
port 78 nsew signal tristate
flabel metal1 s 21426 0 21482 800 0 FreeSans 224 90 0 0 buf_out[5]
port 79 nsew signal tristate
flabel metal1 s 409570 0 409626 800 0 FreeSans 224 90 0 0 buf_out[6]
port 80 nsew signal tristate
flabel metal1 s 21970 0 22026 800 0 FreeSans 224 90 0 0 buf_out[7]
port 81 nsew signal tristate
flabel metal1 s 22242 0 22298 800 0 FreeSans 224 90 0 0 buf_out[8]
port 82 nsew signal tristate
flabel metal1 s 408754 0 408810 800 0 FreeSans 224 90 0 0 buf_out[9]
port 83 nsew signal tristate
flabel metal1 s 480018 0 480074 800 0 FreeSans 224 90 0 0 ch_in[0]
port 84 nsew signal input
flabel metal1 s 490898 0 490954 800 0 FreeSans 224 90 0 0 ch_in[10]
port 85 nsew signal input
flabel metal1 s 187074 9200 187130 10000 0 FreeSans 224 90 0 0 ch_in[11]
port 86 nsew signal input
flabel metal1 s 493074 0 493130 800 0 FreeSans 224 90 0 0 ch_in[12]
port 87 nsew signal input
flabel metal1 s 494162 0 494218 800 0 FreeSans 224 90 0 0 ch_in[13]
port 88 nsew signal input
flabel metal1 s 238074 9200 238130 10000 0 FreeSans 224 90 0 0 ch_in[14]
port 89 nsew signal input
flabel metal1 s 496338 0 496394 800 0 FreeSans 224 90 0 0 ch_in[15]
port 90 nsew signal input
flabel metal1 s 497426 0 497482 800 0 FreeSans 224 90 0 0 ch_in[16]
port 91 nsew signal input
flabel metal1 s 289074 9200 289130 10000 0 FreeSans 224 90 0 0 ch_in[17]
port 92 nsew signal input
flabel metal1 s 499602 0 499658 800 0 FreeSans 224 90 0 0 ch_in[18]
port 93 nsew signal input
flabel metal1 s 500690 0 500746 800 0 FreeSans 224 90 0 0 ch_in[19]
port 94 nsew signal input
flabel metal1 s 481106 0 481162 800 0 FreeSans 224 90 0 0 ch_in[1]
port 95 nsew signal input
flabel metal1 s 340074 9200 340130 10000 0 FreeSans 224 90 0 0 ch_in[20]
port 96 nsew signal input
flabel metal1 s 502866 0 502922 800 0 FreeSans 224 90 0 0 ch_in[21]
port 97 nsew signal input
flabel metal1 s 503954 0 504010 800 0 FreeSans 224 90 0 0 ch_in[22]
port 98 nsew signal input
flabel metal1 s 391074 9200 391130 10000 0 FreeSans 224 90 0 0 ch_in[23]
port 99 nsew signal input
flabel metal1 s 506130 0 506186 800 0 FreeSans 224 90 0 0 ch_in[24]
port 100 nsew signal input
flabel metal1 s 507218 0 507274 800 0 FreeSans 224 90 0 0 ch_in[25]
port 101 nsew signal input
flabel metal1 s 442074 9200 442130 10000 0 FreeSans 224 90 0 0 ch_in[26]
port 102 nsew signal input
flabel metal1 s 34074 9200 34130 10000 0 FreeSans 224 90 0 0 ch_in[2]
port 103 nsew signal input
flabel metal1 s 483282 0 483338 800 0 FreeSans 224 90 0 0 ch_in[3]
port 104 nsew signal input
flabel metal1 s 484370 0 484426 800 0 FreeSans 224 90 0 0 ch_in[4]
port 105 nsew signal input
flabel metal1 s 85074 9200 85130 10000 0 FreeSans 224 90 0 0 ch_in[5]
port 106 nsew signal input
flabel metal1 s 486546 0 486602 800 0 FreeSans 224 90 0 0 ch_in[6]
port 107 nsew signal input
flabel metal1 s 487634 0 487690 800 0 FreeSans 224 90 0 0 ch_in[7]
port 108 nsew signal input
flabel metal1 s 136074 9200 136130 10000 0 FreeSans 224 90 0 0 ch_in[8]
port 109 nsew signal input
flabel metal1 s 489810 0 489866 800 0 FreeSans 224 90 0 0 ch_in[9]
port 110 nsew signal input
flabel metal1 s 74 9200 130 10000 0 FreeSans 224 90 0 0 ch_out[0]
port 111 nsew signal tristate
flabel metal1 s 170074 9200 170130 10000 0 FreeSans 224 90 0 0 ch_out[10]
port 112 nsew signal tristate
flabel metal1 s 491986 0 492042 800 0 FreeSans 224 90 0 0 ch_out[11]
port 113 nsew signal tristate
flabel metal1 s 204074 9200 204130 10000 0 FreeSans 224 90 0 0 ch_out[12]
port 114 nsew signal tristate
flabel metal1 s 221074 9200 221130 10000 0 FreeSans 224 90 0 0 ch_out[13]
port 115 nsew signal tristate
flabel metal1 s 495250 0 495306 800 0 FreeSans 224 90 0 0 ch_out[14]
port 116 nsew signal tristate
flabel metal1 s 255074 9200 255130 10000 0 FreeSans 224 90 0 0 ch_out[15]
port 117 nsew signal tristate
flabel metal1 s 272074 9200 272130 10000 0 FreeSans 224 90 0 0 ch_out[16]
port 118 nsew signal tristate
flabel metal1 s 498514 0 498570 800 0 FreeSans 224 90 0 0 ch_out[17]
port 119 nsew signal tristate
flabel metal1 s 306074 9200 306130 10000 0 FreeSans 224 90 0 0 ch_out[18]
port 120 nsew signal tristate
flabel metal1 s 323074 9200 323130 10000 0 FreeSans 224 90 0 0 ch_out[19]
port 121 nsew signal tristate
flabel metal1 s 17074 9200 17130 10000 0 FreeSans 224 90 0 0 ch_out[1]
port 122 nsew signal tristate
flabel metal1 s 501778 0 501834 800 0 FreeSans 224 90 0 0 ch_out[20]
port 123 nsew signal tristate
flabel metal1 s 357074 9200 357130 10000 0 FreeSans 224 90 0 0 ch_out[21]
port 124 nsew signal tristate
flabel metal1 s 374074 9200 374130 10000 0 FreeSans 224 90 0 0 ch_out[22]
port 125 nsew signal tristate
flabel metal1 s 505042 0 505098 800 0 FreeSans 224 90 0 0 ch_out[23]
port 126 nsew signal tristate
flabel metal1 s 408074 9200 408130 10000 0 FreeSans 224 90 0 0 ch_out[24]
port 127 nsew signal tristate
flabel metal1 s 425074 9200 425130 10000 0 FreeSans 224 90 0 0 ch_out[25]
port 128 nsew signal tristate
flabel metal1 s 508306 0 508362 800 0 FreeSans 224 90 0 0 ch_out[26]
port 129 nsew signal tristate
flabel metal1 s 482194 0 482250 800 0 FreeSans 224 90 0 0 ch_out[2]
port 130 nsew signal tristate
flabel metal1 s 51074 9200 51130 10000 0 FreeSans 224 90 0 0 ch_out[3]
port 131 nsew signal tristate
flabel metal1 s 68074 9200 68130 10000 0 FreeSans 224 90 0 0 ch_out[4]
port 132 nsew signal tristate
flabel metal1 s 485458 0 485514 800 0 FreeSans 224 90 0 0 ch_out[5]
port 133 nsew signal tristate
flabel metal1 s 102074 9200 102130 10000 0 FreeSans 224 90 0 0 ch_out[6]
port 134 nsew signal tristate
flabel metal1 s 119074 9200 119130 10000 0 FreeSans 224 90 0 0 ch_out[7]
port 135 nsew signal tristate
flabel metal1 s 488722 0 488778 800 0 FreeSans 224 90 0 0 ch_out[8]
port 136 nsew signal tristate
flabel metal1 s 153074 9200 153130 10000 0 FreeSans 224 90 0 0 ch_out[9]
port 137 nsew signal tristate
flabel metal2 s -416 656 -96 9136 0 FreeSans 1792 90 0 0 vccd1
port 138 nsew power bidirectional
flabel metal3 s -416 656 530336 976 0 FreeSans 1920 0 0 0 vccd1
port 138 nsew power bidirectional
flabel metal3 s -416 8816 530336 9136 0 FreeSans 1920 0 0 0 vccd1
port 138 nsew power bidirectional
flabel metal2 s 530016 656 530336 9136 0 FreeSans 1792 90 0 0 vccd1
port 138 nsew power bidirectional
flabel metal2 s 66908 -4 67228 9796 0 FreeSans 1792 90 0 0 vccd1
port 138 nsew power bidirectional
flabel metal2 s 198836 -4 199156 9796 0 FreeSans 1792 90 0 0 vccd1
port 138 nsew power bidirectional
flabel metal2 s 330764 -4 331084 9796 0 FreeSans 1792 90 0 0 vccd1
port 138 nsew power bidirectional
flabel metal2 s 462692 -4 463012 9796 0 FreeSans 1792 90 0 0 vccd1
port 138 nsew power bidirectional
flabel metal3 s -1076 2695 530996 3015 0 FreeSans 1920 0 0 0 vccd1
port 138 nsew power bidirectional
flabel metal3 s -1076 4054 530996 4374 0 FreeSans 1920 0 0 0 vccd1
port 138 nsew power bidirectional
flabel metal3 s -1076 5413 530996 5733 0 FreeSans 1920 0 0 0 vccd1
port 138 nsew power bidirectional
flabel metal3 s -1076 6772 530996 7092 0 FreeSans 1920 0 0 0 vccd1
port 138 nsew power bidirectional
flabel metal2 s -1076 -4 -756 9796 0 FreeSans 1792 90 0 0 vssd1
port 139 nsew ground bidirectional
flabel metal3 s -1076 -4 530996 316 0 FreeSans 1920 0 0 0 vssd1
port 139 nsew ground bidirectional
flabel metal3 s -1076 9476 530996 9796 0 FreeSans 1920 0 0 0 vssd1
port 139 nsew ground bidirectional
flabel metal2 s 530676 -4 530996 9796 0 FreeSans 1792 90 0 0 vssd1
port 139 nsew ground bidirectional
flabel metal2 s 67568 -4 67888 9796 0 FreeSans 1792 90 0 0 vssd1
port 139 nsew ground bidirectional
flabel metal2 s 199496 -4 199816 9796 0 FreeSans 1792 90 0 0 vssd1
port 139 nsew ground bidirectional
flabel metal2 s 331424 -4 331744 9796 0 FreeSans 1792 90 0 0 vssd1
port 139 nsew ground bidirectional
flabel metal2 s 463352 -4 463672 9796 0 FreeSans 1792 90 0 0 vssd1
port 139 nsew ground bidirectional
flabel metal3 s -1076 3355 530996 3675 0 FreeSans 1920 0 0 0 vssd1
port 139 nsew ground bidirectional
flabel metal3 s -1076 4714 530996 5034 0 FreeSans 1920 0 0 0 vssd1
port 139 nsew ground bidirectional
flabel metal3 s -1076 6073 530996 6393 0 FreeSans 1920 0 0 0 vssd1
port 139 nsew ground bidirectional
flabel metal3 s -1076 7432 530996 7752 0 FreeSans 1920 0 0 0 vssd1
port 139 nsew ground bidirectional
rlabel metal1 264960 7072 264960 7072 0 vccd1
rlabel metal1 264960 7616 264960 7616 0 vssd1
rlabel metal1 20155 782 20155 782 0 buf_in[0]
rlabel metal2 346702 2312 346702 2312 0 buf_in[10]
rlabel metal2 348266 3332 348266 3332 0 buf_in[11]
rlabel metal1 40802 4522 40802 4522 0 buf_in[12]
rlabel metal2 342102 2686 342102 2686 0 buf_in[13]
rlabel metal2 353326 3876 353326 3876 0 buf_in[14]
rlabel metal1 42090 2312 42090 2312 0 buf_in[15]
rlabel metal2 337318 1224 337318 1224 0 buf_in[16]
rlabel metal2 336398 2992 336398 2992 0 buf_in[17]
rlabel metal2 48346 2040 48346 2040 0 buf_in[18]
rlabel metal1 331430 2958 331430 2958 0 buf_in[19]
rlabel metal2 358202 2074 358202 2074 0 buf_in[1]
rlabel metal1 329728 2414 329728 2414 0 buf_in[20]
rlabel metal2 41998 2108 41998 2108 0 buf_in[21]
rlabel metal1 324760 2822 324760 2822 0 buf_in[22]
rlabel metal1 404908 782 404908 782 0 buf_in[23]
rlabel metal1 26687 782 26687 782 0 buf_in[24]
rlabel metal1 404356 782 404356 782 0 buf_in[25]
rlabel metal1 404080 782 404080 782 0 buf_in[26]
rlabel metal2 126086 2074 126086 2074 0 buf_in[27]
rlabel metal2 399970 187 399970 187 0 buf_in[28]
rlabel metal2 350566 4250 350566 4250 0 buf_in[29]
rlabel metal2 356086 1428 356086 1428 0 buf_in[2]
rlabel metal1 28320 782 28320 782 0 buf_in[30]
rlabel metal1 393300 782 393300 782 0 buf_in[31]
rlabel metal2 309442 3230 309442 3230 0 buf_in[32]
rlabel metal1 116380 4114 116380 4114 0 buf_in[33]
rlabel metal1 307556 4454 307556 4454 0 buf_in[34]
rlabel metal1 401771 782 401771 782 0 buf_in[35]
rlabel metal2 112378 1700 112378 1700 0 buf_in[36]
rlabel metal1 397302 2346 397302 2346 0 buf_in[37]
rlabel metal1 400837 782 400837 782 0 buf_in[38]
rlabel metal2 108422 1802 108422 1802 0 buf_in[39]
rlabel metal1 20973 782 20973 782 0 buf_in[3]
rlabel metal1 393622 2822 393622 2822 0 buf_in[40]
rlabel metal2 390494 2108 390494 2108 0 buf_in[41]
rlabel metal1 410060 782 410060 782 0 buf_in[4]
rlabel metal2 352406 1360 352406 1360 0 buf_in[5]
rlabel metal1 21788 782 21788 782 0 buf_in[6]
rlabel metal2 349738 1326 349738 1326 0 buf_in[7]
rlabel metal2 348450 1292 348450 1292 0 buf_in[8]
rlabel metal2 62606 2142 62606 2142 0 buf_in[9]
rlabel metal1 411164 782 411164 782 0 buf_out[0]
rlabel metal2 116334 3672 116334 3672 0 buf_out[10]
rlabel metal2 117622 2040 117622 2040 0 buf_out[11]
rlabel metal2 342378 4046 342378 4046 0 buf_out[12]
rlabel metal2 118174 2584 118174 2584 0 buf_out[13]
rlabel metal2 117346 2142 117346 2142 0 buf_out[14]
rlabel metal2 338054 4012 338054 4012 0 buf_out[15]
rlabel metal1 24535 782 24535 782 0 buf_out[16]
rlabel metal2 117530 1802 117530 1802 0 buf_out[17]
rlabel metal2 332534 3978 332534 3978 0 buf_out[18]
rlabel metal1 25353 782 25353 782 0 buf_out[19]
rlabel metal1 20431 782 20431 782 0 buf_out[1]
rlabel metal1 25629 782 25629 782 0 buf_out[20]
rlabel metal1 405451 782 405451 782 0 buf_out[21]
rlabel metal2 118726 1292 118726 1292 0 buf_out[22]
rlabel metal1 26457 782 26457 782 0 buf_out[23]
rlabel metal1 404632 782 404632 782 0 buf_out[24]
rlabel metal2 31878 1139 31878 1139 0 buf_out[25]
rlabel metal2 120198 1258 120198 1258 0 buf_out[26]
rlabel metal1 403804 782 403804 782 0 buf_out[27]
rlabel metal1 27777 782 27777 782 0 buf_out[28]
rlabel metal2 121486 1394 121486 1394 0 buf_out[29]
rlabel metal1 20593 782 20593 782 0 buf_out[2]
rlabel metal2 310730 5644 310730 5644 0 buf_out[30]
rlabel via2 28658 459 28658 459 0 buf_out[31]
rlabel metal2 122866 1632 122866 1632 0 buf_out[32]
rlabel metal2 304750 4760 304750 4760 0 buf_out[33]
rlabel metal2 31786 442 31786 442 0 buf_out[34]
rlabel metal1 29700 782 29700 782 0 buf_out[35]
rlabel metal2 308522 4930 308522 4930 0 buf_out[36]
rlabel metal2 123878 1564 123878 1564 0 buf_out[37]
rlabel metal2 36478 748 36478 748 0 buf_out[38]
rlabel metal2 307694 2193 307694 2193 0 buf_out[39]
rlabel metal2 353970 3434 353970 3434 0 buf_out[3]
rlabel metal1 31065 782 31065 782 0 buf_out[40]
rlabel metal2 125258 1224 125258 1224 0 buf_out[41]
rlabel metal1 21247 782 21247 782 0 buf_out[4]
rlabel metal1 21521 782 21521 782 0 buf_out[5]
rlabel metal2 350474 2992 350474 2992 0 buf_out[6]
rlabel metal1 21912 510 21912 510 0 buf_out[7]
rlabel metal2 116150 3298 116150 3298 0 buf_out[8]
rlabel metal2 346794 1224 346794 1224 0 buf_out[9]
rlabel metal2 382766 2890 382766 2890 0 ch_in[0]
rlabel metal2 466578 1972 466578 1972 0 ch_in[10]
rlabel metal2 200238 4284 200238 4284 0 ch_in[11]
rlabel metal2 408526 2720 408526 2720 0 ch_in[12]
rlabel metal2 426558 2142 426558 2142 0 ch_in[13]
rlabel metal2 254058 4590 254058 4590 0 ch_in[14]
rlabel metal2 461886 1904 461886 1904 0 ch_in[15]
rlabel metal1 497046 782 497046 782 0 ch_in[16]
rlabel metal1 289301 9214 289301 9214 0 ch_in[17]
rlabel metal2 422602 2822 422602 2822 0 ch_in[18]
rlabel metal2 488566 1564 488566 1564 0 ch_in[19]
rlabel metal1 399970 2822 399970 2822 0 ch_in[1]
rlabel metal2 362250 4624 362250 4624 0 ch_in[20]
rlabel metal1 502623 782 502623 782 0 ch_in[21]
rlabel metal1 503578 782 503578 782 0 ch_in[22]
rlabel metal2 416346 4658 416346 4658 0 ch_in[23]
rlabel metal1 505773 782 505773 782 0 ch_in[24]
rlabel metal1 507189 782 507189 782 0 ch_in[25]
rlabel metal2 470442 4522 470442 4522 0 ch_in[26]
rlabel metal2 37674 4828 37674 4828 0 ch_in[2]
rlabel metal2 435758 1870 435758 1870 0 ch_in[3]
rlabel metal1 453146 3026 453146 3026 0 ch_in[4]
rlabel metal2 92046 4624 92046 4624 0 ch_in[5]
rlabel metal1 486190 782 486190 782 0 ch_in[6]
rlabel metal1 487279 782 487279 782 0 ch_in[7]
rlabel metal1 136351 9214 136351 9214 0 ch_in[8]
rlabel metal2 448638 2074 448638 2074 0 ch_in[9]
rlabel metal1 996 9214 996 9214 0 ch_out[0]
rlabel metal2 179446 4386 179446 4386 0 ch_out[10]
rlabel metal1 491664 782 491664 782 0 ch_out[11]
rlabel metal1 218132 2278 218132 2278 0 ch_out[12]
rlabel metal2 236302 4216 236302 4216 0 ch_out[13]
rlabel metal1 494907 714 494907 714 0 ch_out[14]
rlabel metal1 272090 2278 272090 2278 0 ch_out[15]
rlabel metal1 289386 2278 289386 2278 0 ch_out[16]
rlabel metal2 411470 952 411470 952 0 ch_out[17]
rlabel metal1 306208 8942 306208 8942 0 ch_out[18]
rlabel metal1 344494 2312 344494 2312 0 ch_out[19]
rlabel metal2 19918 4726 19918 4726 0 ch_out[1]
rlabel metal1 411378 714 411378 714 0 ch_out[20]
rlabel metal2 380558 4420 380558 4420 0 ch_out[21]
rlabel metal1 374715 9214 374715 9214 0 ch_out[22]
rlabel metal1 505050 782 505050 782 0 ch_out[23]
rlabel metal1 408273 8942 408273 8942 0 ch_out[24]
rlabel metal2 442842 5508 442842 5508 0 ch_out[25]
rlabel metal1 508293 782 508293 782 0 ch_out[26]
rlabel metal2 388470 3298 388470 3298 0 ch_out[2]
rlabel metal1 53130 6834 53130 6834 0 ch_out[3]
rlabel metal2 74014 4726 74014 4726 0 ch_out[4]
rlabel metal2 391690 1632 391690 1632 0 ch_out[5]
rlabel metal1 102187 9214 102187 9214 0 ch_out[6]
rlabel metal1 127512 2278 127512 2278 0 ch_out[7]
rlabel metal1 488697 782 488697 782 0 ch_out[8]
rlabel via1 153111 8942 153111 8942 0 ch_out[9]
rlabel metal2 146142 1428 146142 1428 0 net1
rlabel metal2 199410 1666 199410 1666 0 net10
rlabel metal2 411838 4726 411838 4726 0 net100
rlabel metal2 110814 3842 110814 3842 0 net101
rlabel metal1 206172 2822 206172 2822 0 net102
rlabel metal2 299598 1700 299598 1700 0 net103
rlabel metal2 74658 2108 74658 2108 0 net104
rlabel metal2 170798 1326 170798 1326 0 net105
rlabel metal2 265742 1530 265742 1530 0 net106
rlabel metal2 359582 2754 359582 2754 0 net107
rlabel metal2 63618 3876 63618 3876 0 net108
rlabel metal2 152214 1428 152214 1428 0 net109
rlabel metal2 116150 1224 116150 1224 0 net11
rlabel metal2 247158 1360 247158 1360 0 net110
rlabel metal2 390586 1513 390586 1513 0 net111
rlabel metal1 412620 1462 412620 1462 0 net112
rlabel metal1 380834 2414 380834 2414 0 net113
rlabel metal1 20378 2414 20378 2414 0 net114
rlabel metal1 117024 2414 117024 2414 0 net115
rlabel metal1 211094 2380 211094 2380 0 net116
rlabel metal2 389206 1564 389206 1564 0 net117
rlabel metal2 346242 1870 346242 1870 0 net118
rlabel metal2 421406 3978 421406 3978 0 net119
rlabel metal2 362526 5168 362526 5168 0 net12
rlabel metal1 290582 2448 290582 2448 0 net120
rlabel metal2 386538 2176 386538 2176 0 net121
rlabel metal2 273102 3298 273102 3298 0 net122
rlabel metal1 367862 2448 367862 2448 0 net123
rlabel metal2 237038 1666 237038 1666 0 net124
rlabel metal1 332718 2822 332718 2822 0 net125
rlabel metal2 218454 1326 218454 1326 0 net126
rlabel metal2 407238 4930 407238 4930 0 net127
rlabel metal2 277150 1734 277150 1734 0 net128
rlabel metal2 349830 1156 349830 1156 0 net129
rlabel metal2 308430 5474 308430 5474 0 net13
rlabel via2 372462 2363 372462 2363 0 net130
rlabel metal2 2622 1972 2622 1972 0 net131
rlabel metal2 98670 3298 98670 3298 0 net132
rlabel metal2 193614 1394 193614 1394 0 net133
rlabel metal2 287454 3468 287454 3468 0 net134
rlabel metal1 255898 2312 255898 2312 0 net135
rlabel metal2 157918 1598 157918 1598 0 net136
rlabel metal2 63526 3604 63526 3604 0 net137
rlabel metal2 257094 1530 257094 1530 0 net138
rlabel metal2 255806 1734 255806 1734 0 net139
rlabel metal2 254334 1564 254334 1564 0 net14
rlabel metal2 120106 1598 120106 1598 0 net140
rlabel metal2 295826 1428 295826 1428 0 net141
rlabel metal2 298678 4318 298678 4318 0 net142
rlabel metal1 352038 3162 352038 3162 0 net143
rlabel metal2 165554 1564 165554 1564 0 net144
rlabel metal2 74566 2550 74566 2550 0 net145
rlabel metal1 211646 4216 211646 4216 0 net146
rlabel metal2 108974 2210 108974 2210 0 net147
rlabel metal2 351946 4964 351946 4964 0 net148
rlabel metal1 302013 2414 302013 2414 0 net149
rlabel metal2 332626 1054 332626 1054 0 net15
rlabel metal2 211554 4522 211554 4522 0 net150
rlabel metal2 112930 2006 112930 2006 0 net151
rlabel metal1 303324 3026 303324 3026 0 net152
rlabel metal2 304198 4250 304198 4250 0 net153
rlabel metal1 117438 4012 117438 4012 0 net154
rlabel metal1 310500 4114 310500 4114 0 net155
rlabel metal2 215234 2380 215234 2380 0 net156
rlabel metal2 221030 3536 221030 3536 0 net157
rlabel metal2 214498 4828 214498 4828 0 net158
rlabel metal2 226182 2210 226182 2210 0 net159
rlabel metal2 211554 2142 211554 2142 0 net16
rlabel metal2 131422 3570 131422 3570 0 net160
rlabel metal2 130226 2125 130226 2125 0 net161
rlabel metal2 231978 2176 231978 2176 0 net162
rlabel metal2 137310 3740 137310 3740 0 net163
rlabel metal2 42918 2142 42918 2142 0 net164
rlabel metal2 332350 3774 332350 3774 0 net165
rlabel metal2 237774 3502 237774 3502 0 net166
rlabel metal1 143290 2414 143290 2414 0 net167
rlabel metal2 244214 2108 244214 2108 0 net168
rlabel metal1 149362 2516 149362 2516 0 net169
rlabel metal2 396934 2125 396934 2125 0 net17
rlabel via2 148258 2533 148258 2533 0 net170
rlabel metal1 249366 2482 249366 2482 0 net171
rlabel metal2 154054 2142 154054 2142 0 net172
rlabel metal2 152766 1904 152766 1904 0 net173
rlabel metal1 349922 2924 349922 2924 0 net174
rlabel metal2 169234 4420 169234 4420 0 net175
rlabel metal2 75302 2108 75302 2108 0 net176
rlabel metal2 211830 2550 211830 2550 0 net18
rlabel metal2 335294 2142 335294 2142 0 net19
rlabel metal2 300794 2295 300794 2295 0 net2
rlabel metal2 118082 2618 118082 2618 0 net20
rlabel metal2 213578 2703 213578 2703 0 net21
rlabel metal2 337226 2142 337226 2142 0 net22
rlabel metal2 213394 4862 213394 4862 0 net23
rlabel metal2 213946 2788 213946 2788 0 net24
rlabel metal1 309212 4454 309212 4454 0 net25
rlabel metal2 117898 3740 117898 3740 0 net26
rlabel metal2 212842 4930 212842 4930 0 net27
rlabel metal1 308660 4998 308660 4998 0 net28
rlabel metal2 211462 1802 211462 1802 0 net29
rlabel metal2 206126 1938 206126 1938 0 net3
rlabel metal1 212612 3026 212612 3026 0 net30
rlabel metal1 307418 3468 307418 3468 0 net31
rlabel metal1 118174 3536 118174 3536 0 net32
rlabel metal2 212198 2652 212198 2652 0 net33
rlabel metal2 306498 4012 306498 4012 0 net34
rlabel metal1 116886 3094 116886 3094 0 net35
rlabel metal2 210818 1972 210818 1972 0 net36
rlabel metal1 307786 3026 307786 3026 0 net37
rlabel metal2 116702 3706 116702 3706 0 net38
rlabel metal1 211002 3468 211002 3468 0 net39
rlabel metal1 92230 2380 92230 2380 0 net4
rlabel metal1 306590 4454 306590 4454 0 net40
rlabel metal2 115690 2312 115690 2312 0 net41
rlabel metal2 209438 4318 209438 4318 0 net42
rlabel metal2 352314 1938 352314 1938 0 net43
rlabel metal1 114172 2414 114172 2414 0 net44
rlabel metal2 209622 4352 209622 4352 0 net45
rlabel metal2 354430 1904 354430 1904 0 net46
rlabel metal1 115506 3536 115506 3536 0 net47
rlabel metal2 208426 4726 208426 4726 0 net48
rlabel metal2 304842 5066 304842 5066 0 net49
rlabel metal2 391138 2465 391138 2465 0 net5
rlabel metal2 116058 4046 116058 4046 0 net50
rlabel metal1 210174 4046 210174 4046 0 net51
rlabel metal2 304382 2924 304382 2924 0 net52
rlabel metal1 115644 3706 115644 3706 0 net53
rlabel metal2 209070 4964 209070 4964 0 net54
rlabel metal2 295458 3706 295458 3706 0 net55
rlabel metal1 125534 2380 125534 2380 0 net56
rlabel metal1 249274 2414 249274 2414 0 net57
rlabel metal2 126270 4556 126270 4556 0 net58
rlabel metal2 306590 3570 306590 3570 0 net59
rlabel metal1 296516 2414 296516 2414 0 net6
rlabel metal2 300242 5202 300242 5202 0 net60
rlabel metal2 125902 5440 125902 5440 0 net61
rlabel metal1 301484 2618 301484 2618 0 net62
rlabel metal1 124476 2414 124476 2414 0 net63
rlabel metal2 307786 3706 307786 3706 0 net64
rlabel metal1 296700 2924 296700 2924 0 net65
rlabel metal2 216614 2040 216614 2040 0 net66
rlabel metal1 306590 2890 306590 2890 0 net67
rlabel metal2 125166 5542 125166 5542 0 net68
rlabel metal1 217902 3026 217902 3026 0 net69
rlabel via2 107686 2397 107686 2397 0 net7
rlabel metal1 123372 2414 123372 2414 0 net70
rlabel metal1 216338 2414 216338 2414 0 net71
rlabel metal2 215418 2227 215418 2227 0 net72
rlabel metal2 308522 3298 308522 3298 0 net73
rlabel metal1 122130 2414 122130 2414 0 net74
rlabel metal1 314364 2618 314364 2618 0 net75
rlabel metal2 122590 3281 122590 3281 0 net76
rlabel metal1 312294 3026 312294 3026 0 net77
rlabel metal2 212566 3434 212566 3434 0 net78
rlabel metal1 311650 2924 311650 2924 0 net79
rlabel metal1 104236 2414 104236 2414 0 net8
rlabel metal2 311190 3332 311190 3332 0 net80
rlabel metal2 214038 2295 214038 2295 0 net81
rlabel metal2 214314 4437 214314 4437 0 net82
rlabel metal1 311006 3060 311006 3060 0 net83
rlabel metal1 210358 3128 210358 3128 0 net84
rlabel metal2 310730 3400 310730 3400 0 net85
rlabel metal1 310270 3536 310270 3536 0 net86
rlabel metal1 119278 2448 119278 2448 0 net87
rlabel metal1 309580 3570 309580 3570 0 net88
rlabel metal2 309718 3774 309718 3774 0 net89
rlabel metal1 387550 2414 387550 2414 0 net9
rlabel metal2 212842 1904 212842 1904 0 net90
rlabel metal1 308890 4012 308890 4012 0 net91
rlabel metal1 309764 3502 309764 3502 0 net92
rlabel metal2 214038 3162 214038 3162 0 net93
rlabel metal1 214590 3468 214590 3468 0 net94
rlabel metal2 164358 3196 164358 3196 0 net95
rlabel metal2 353326 2159 353326 2159 0 net96
rlabel metal2 353694 2618 353694 2618 0 net97
rlabel metal2 128846 2142 128846 2142 0 net98
rlabel metal2 224250 2193 224250 2193 0 net99
<< properties >>
string FIXED_BBOX 0 0 530000 10000
<< end >>
