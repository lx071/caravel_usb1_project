// This is the unpowered netlist.
module bus_rep_north (buf_in,
    buf_out,
    ch_in,
    ch_out);
 input [41:0] buf_in;
 output [41:0] buf_out;
 input [26:0] ch_in;
 output [26:0] ch_out;

 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA__00__A (.DIODE(buf_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__01__A (.DIODE(buf_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__02__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__03__A (.DIODE(buf_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__04__A (.DIODE(buf_in[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA__05__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__06__A (.DIODE(buf_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__07__A (.DIODE(buf_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__08__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__09__A (.DIODE(buf_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__10__A (.DIODE(buf_in[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA__11__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__12__A (.DIODE(buf_in[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA__13__A (.DIODE(buf_in[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA__14__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__15__A (.DIODE(buf_in[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA__16__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__17__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__18__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__19__A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__20__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__21__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__22__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__23__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__24__A (.DIODE(buf_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__25__A (.DIODE(buf_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__26__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__27__A (.DIODE(buf_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__28__A (.DIODE(buf_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__29__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__30__A (.DIODE(buf_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__31__A (.DIODE(buf_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__32__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__33__A (.DIODE(buf_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__34__A (.DIODE(buf_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA__35__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__36__A (.DIODE(buf_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA__37__A (.DIODE(buf_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA__38__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__39__A (.DIODE(buf_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__40__A (.DIODE(buf_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__41__A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[0].u_buf_A  (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[10].u_buf_A  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[11].u_buf_A  (.DIODE(ch_in[11]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[12].u_buf_A  (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[13].u_buf_A  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[14].u_buf_A  (.DIODE(ch_in[14]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[15].u_buf_A  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[16].u_buf_A  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[17].u_buf_A  (.DIODE(ch_in[17]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[18].u_buf_A  (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[19].u_buf_A  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[1].u_buf_A  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[20].u_buf_A  (.DIODE(ch_in[20]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[21].u_buf_A  (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[22].u_buf_A  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[23].u_buf_A  (.DIODE(ch_in[23]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[24].u_buf_A  (.DIODE(ch_in[24]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[25].u_buf_A  (.DIODE(ch_in[25]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[26].u_buf_A  (.DIODE(ch_in[26]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[2].u_buf_A  (.DIODE(ch_in[2]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[3].u_buf_A  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[4].u_buf_A  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[5].u_buf_A  (.DIODE(ch_in[5]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[6].u_buf_A  (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[7].u_buf_A  (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[8].u_buf_A  (.DIODE(ch_in[8]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[9].u_buf_A  (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire100_A (.DIODE(ch_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire101_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire102_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire103_A (.DIODE(ch_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire104_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire105_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire106_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire107_A (.DIODE(ch_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire108_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire109_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire10_A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire110_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire111_A (.DIODE(ch_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire112_A (.DIODE(ch_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire113_A (.DIODE(ch_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire114_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire115_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire116_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire117_A (.DIODE(ch_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire118_A (.DIODE(ch_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire119_A (.DIODE(ch_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire11_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire120_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire121_A (.DIODE(ch_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire122_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire123_A (.DIODE(ch_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire124_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire125_A (.DIODE(ch_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire126_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire127_A (.DIODE(ch_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire128_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire129_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire12_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire130_A (.DIODE(ch_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire131_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire132_A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire133_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire134_A (.DIODE(ch_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire135_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire136_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire137_A (.DIODE(buf_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire138_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire139_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire13_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire140_A (.DIODE(buf_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire141_A (.DIODE(buf_in[41]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire142_A (.DIODE(buf_in[40]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire143_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire144_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire145_A (.DIODE(buf_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire146_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire147_A (.DIODE(buf_in[39]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire148_A (.DIODE(buf_in[38]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire149_A (.DIODE(buf_in[37]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire14_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire150_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire151_A (.DIODE(buf_in[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire152_A (.DIODE(buf_in[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire153_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire154_A (.DIODE(buf_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire155_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire156_A (.DIODE(buf_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire157_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire158_A (.DIODE(buf_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire159_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire15_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire160_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire161_A (.DIODE(buf_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire162_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire163_A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire164_A (.DIODE(buf_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire165_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire166_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire167_A (.DIODE(buf_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire168_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire169_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire16_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire170_A (.DIODE(buf_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire171_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire172_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire173_A (.DIODE(buf_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire174_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire175_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire176_A (.DIODE(buf_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire17_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire19_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire20_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire21_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire22_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire23_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire24_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire25_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire26_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire27_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire28_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire29_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire30_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire31_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire32_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire33_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire34_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire35_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire36_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire37_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire38_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire39_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire3_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire40_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire41_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire42_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire43_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire44_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire45_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire46_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire47_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire48_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire49_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire4_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire50_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire51_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire52_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire53_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire54_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire55_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire56_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire57_A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire58_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire5_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire60_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire61_A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire62_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire63_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire65_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire66_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire67_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire68_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire69_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire6_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire70_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire71_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire72_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire73_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire74_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire75_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire76_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire77_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire78_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire80_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire81_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire83_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire84_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire86_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire87_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire89_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire8_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire90_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire91_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire92_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire93_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire94_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire95_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire96_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire97_A (.DIODE(ch_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire98_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire99_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire9_A (.DIODE(net10));
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1566 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1957 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1971 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2087 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2420 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2700 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2732 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2816 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2871 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2997 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3008 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3703 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3723 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3759 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3807 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3815 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3843 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3863 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3876 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3988 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4715 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4859 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4911 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4985 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5003 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5047 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5054 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1260 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1303 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1316 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1525 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1545 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1557 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1565 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1575 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1587 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1599 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1611 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1625 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1657 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1669 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1761 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1775 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1781 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1813 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1816 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2177 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2182 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2196 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2208 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2223 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2229 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2235 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2238 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2252 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2258 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2268 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2281 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2294 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2297 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2301 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2311 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2324 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2337 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2350 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2353 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2357 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2360 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2373 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2386 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2392 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2398 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2406 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2657 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2669 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2677 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2701 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2723 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2735 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2743 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2751 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2763 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2775 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2787 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2799 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2812 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2818 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2842 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2854 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3193 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3207 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3219 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3223 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3229 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3235 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3243 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3246 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3249 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3257 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3264 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3270 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3278 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3298 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3305 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3313 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3323 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3333 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3343 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3359 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3361 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3369 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3379 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3395 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3403 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3411 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3415 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3421 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3433 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3438 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3444 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3458 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3464 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3505 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3508 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3516 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3520 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3526 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3583 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3585 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3592 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3598 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3604 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3616 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3628 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3641 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3653 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3658 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3664 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3676 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3682 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3687 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3693 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3697 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3701 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3707 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3719 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3733 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3739 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3751 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3757 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3769 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3779 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3793 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3799 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3807 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3809 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3817 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3822 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3826 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3829 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3843 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3855 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3861 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3865 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3871 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3876 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3882 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3894 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3906 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3918 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3927 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3939 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3963 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4113 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4129 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4213 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_4235 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_4241 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_4247 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4255 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4257 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_4265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4273 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_4283 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4291 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_4295 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4299 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4306 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4313 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4317 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_4325 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_4333 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4338 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4344 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4347 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_4359 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4423 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4429 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4441 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4465 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4493 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4515 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_4527 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4549 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4573 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4585 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4591 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4593 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4605 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4629 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4641 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4647 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4649 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4661 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4685 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4697 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4703 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_4705 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4713 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_4717 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4739 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_4751 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4759 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4761 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4773 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4797 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4809 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4815 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4817 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4829 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4853 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4865 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4871 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4873 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4885 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_4897 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_4911 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_4917 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_4925 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4929 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4941 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4965 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4977 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4983 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4985 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4997 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5021 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_5033 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5039 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5041 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5053 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5077 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_5089 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5095 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_5097 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5103 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5115 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5127 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5139 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5151 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5189 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_5201 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5207 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5233 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5245 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_5257 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5263 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5265 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5301 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_5313 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5319 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5345 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5357 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_5369 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5375 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5389 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5413 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_5425 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5431 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5433 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5445 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5457 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5469 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_5481 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5487 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5489 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5501 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5513 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5525 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_5537 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5543 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5545 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5557 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5569 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5581 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_5593 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5599 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5601 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5613 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5625 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5637 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_5649 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5655 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5657 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5669 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5681 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5693 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_5705 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5711 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5713 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_5725 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1300 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1328 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2237 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2249 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2253 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2266 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2269 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2273 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2283 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2296 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2309 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2322 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2336 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2349 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2362 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2375 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2379 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2385 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2397 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3009 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3065 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3089 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3201 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3233 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3245 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3259 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3271 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3275 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3277 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3281 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3287 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3300 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3310 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3320 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3330 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3333 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3341 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3351 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3361 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3371 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3377 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3383 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3387 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3393 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3405 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3429 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3625 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3649 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3761 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3849 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_3861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3872 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_3884 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4097 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4129 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4185 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_4267 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4271 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_4274 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_4280 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4285 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4301 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4507 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4563 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4565 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4601 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4613 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4619 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4621 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4633 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4657 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4669 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4675 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4677 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4689 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4713 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4725 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4731 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4733 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4745 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4781 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4787 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4789 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4801 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4825 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4837 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4843 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4845 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4857 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4893 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4899 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4901 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4913 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4937 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4949 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4955 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4957 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4969 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4993 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5011 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5013 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5025 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5049 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5061 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5067 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5069 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5081 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5105 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5117 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5123 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5125 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5137 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5161 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5173 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5179 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5181 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5193 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5217 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5229 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5235 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5237 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5249 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5261 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5273 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5285 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5291 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5293 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5305 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5317 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5329 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5341 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5347 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5349 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5361 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5373 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5385 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5397 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5403 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5405 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5417 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5429 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5441 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5453 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5459 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5461 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5473 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5485 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5497 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5509 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5515 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5517 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5529 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5541 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5553 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5565 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5571 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5573 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5585 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5597 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5609 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5621 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5627 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5629 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5641 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5653 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5665 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5677 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5683 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5685 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5697 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5709 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5721 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1296 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1302 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2255 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2261 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2274 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2282 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2292 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_2297 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2302 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2315 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2332 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_2349 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2353 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2357 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2361 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2364 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2372 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2375 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2387 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2399 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3273 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3293 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3296 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3302 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3305 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3309 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3313 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3320 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3326 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3334 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3342 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3349 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3355 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3359 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3361 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3367 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3901 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4461 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4479 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4493 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4517 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4529 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4549 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4573 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4585 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4591 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4593 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4605 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4629 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4641 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4647 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4649 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4661 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4685 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4697 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4703 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4705 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4717 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4741 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4753 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4759 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4761 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4773 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4797 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4809 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4815 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4817 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4829 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4853 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4865 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4871 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4873 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4885 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4909 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4921 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4927 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4929 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4941 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4965 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4977 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4983 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4985 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4997 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5021 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5033 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5039 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5041 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5053 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5077 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5089 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5095 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5097 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5109 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5133 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5145 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5151 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5153 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5165 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5189 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5201 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5207 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5209 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5221 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5233 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5245 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5257 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5263 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5265 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5277 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5289 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5301 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5313 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5319 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5321 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5333 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5345 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5357 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5369 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5375 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5377 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5389 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5401 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5413 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5425 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5431 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5433 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5445 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5457 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5469 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5481 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5487 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5489 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5501 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5513 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5525 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5537 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5543 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5545 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5557 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5569 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5581 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5593 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5599 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5601 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5613 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5625 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5637 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5649 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5655 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5657 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5669 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5681 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5693 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5705 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5711 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5713 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_5725 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1254 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1288 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1302 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1321 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2267 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2269 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2273 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2276 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2280 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2283 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2295 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2298 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2304 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2310 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2316 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_2322 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2331 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_2334 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2342 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2345 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2357 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_2369 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3009 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3065 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3089 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3201 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3289 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_3301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3312 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3318 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3324 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3330 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3333 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3343 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3349 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3355 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3375 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3625 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3649 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3761 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3885 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4097 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4185 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4507 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4563 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4565 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4601 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4613 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4619 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4621 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4633 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4657 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4669 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4675 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4677 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4689 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4713 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4725 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4731 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4733 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4745 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4781 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4787 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4789 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4801 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4825 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4837 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4843 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4845 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4857 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4893 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4899 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4901 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4913 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4937 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4949 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4955 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4957 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4969 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4993 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5011 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5013 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5025 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5049 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5061 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5067 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5069 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5081 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5105 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5117 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5123 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5125 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5137 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5161 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5173 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5179 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5181 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5193 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5217 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5229 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5235 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5237 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5249 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5261 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5273 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5285 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5291 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5293 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5305 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5317 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5329 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5341 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5347 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5349 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5361 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5373 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5385 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5397 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5403 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5405 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5417 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5429 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5441 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5453 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5459 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5461 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5473 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5485 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5497 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5509 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5515 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5517 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5529 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5541 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5553 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5565 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5571 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5573 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5585 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5597 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5609 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5621 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5627 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5629 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5641 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5653 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5665 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5677 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5683 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5685 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5697 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5709 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5721 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1260 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2265 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2277 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2283 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2297 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2311 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2315 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2318 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2324 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2330 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2336 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2339 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3303 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_3305 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_3313 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3318 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3324 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3332 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3338 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3342 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3345 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3901 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4461 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4479 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4493 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4517 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4529 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4549 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4573 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4585 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4591 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4593 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4605 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4629 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4641 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4647 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4649 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4661 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4685 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4697 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4703 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4705 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4717 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4741 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4753 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4759 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4761 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4773 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4797 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4809 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4815 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4817 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4829 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4853 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4865 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4871 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4873 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4885 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4909 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4921 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4927 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4929 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4941 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4965 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4977 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4983 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4985 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4997 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5021 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5033 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5039 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5041 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5053 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5077 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5089 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5095 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5097 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5109 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5133 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5145 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5151 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5153 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5165 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5189 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5201 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5207 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5209 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5221 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5233 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5245 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5257 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5263 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5265 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5277 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5289 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5301 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5313 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5319 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5321 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5333 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5345 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5357 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5369 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5375 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5377 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5389 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5401 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5413 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5425 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5431 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5433 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5445 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5457 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5469 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5481 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5487 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5489 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5501 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5513 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5525 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5537 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5543 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5545 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5557 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5569 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5581 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5593 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5599 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5601 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5613 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5625 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5637 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5649 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5655 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5657 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5669 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5681 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5693 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5705 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5711 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5713 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_5725 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3009 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3065 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3089 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3201 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3325 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3625 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3649 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3761 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3885 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4097 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4185 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4507 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4563 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4565 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4601 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4613 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4619 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4621 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4633 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4657 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4669 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4675 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4677 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4689 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4713 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4725 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4731 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4733 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4745 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4781 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4787 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4789 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4801 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4825 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4837 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4843 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4845 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4857 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4893 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4899 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4901 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4913 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4937 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4949 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4955 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4957 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4969 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4993 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5011 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5013 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5025 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5049 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5061 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5067 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5069 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5081 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5105 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5117 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5123 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5125 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5137 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5161 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5173 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5179 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5181 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5193 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5217 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5229 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5235 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5237 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5249 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5261 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5273 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5285 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5291 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5293 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5305 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5317 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5329 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5341 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5347 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5349 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5361 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5373 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5385 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5397 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5403 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5405 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5417 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5429 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5441 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5453 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5459 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5461 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5473 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5485 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5497 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5509 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5515 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5517 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5529 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5541 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5553 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5565 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5571 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5573 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5585 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5597 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5609 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5621 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5627 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5629 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5641 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5653 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5665 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5677 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5683 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5685 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5697 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5709 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5721 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3341 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3901 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4461 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4479 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4493 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4517 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4529 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4549 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4573 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4585 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4591 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4593 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4605 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4629 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4641 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4647 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4649 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4661 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4685 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4697 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4703 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4705 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4717 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4741 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4753 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4759 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4761 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4773 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4797 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4809 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4815 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4817 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4829 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4853 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4865 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4871 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4873 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4885 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4909 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4921 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4927 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4929 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4941 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4965 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4977 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4983 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4985 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4997 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5021 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5033 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5039 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5041 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5053 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5077 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5089 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5095 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5097 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5109 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5133 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5145 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5151 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5153 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5165 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5177 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5189 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5201 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5207 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5209 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5221 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5233 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5245 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5257 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5263 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5265 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5277 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5289 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5301 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5313 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5319 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5321 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5333 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5345 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5357 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5369 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5375 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5377 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5389 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5401 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5413 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5425 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5431 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5433 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5445 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5457 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5469 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5481 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5487 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5489 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5501 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5513 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5525 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5537 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5543 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5545 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5557 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5569 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5581 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5593 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5599 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5601 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5613 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5625 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5637 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5649 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5655 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5657 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5669 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5681 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5693 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5705 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5711 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5713 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_5725 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3009 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3065 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3089 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3201 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3325 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3625 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3649 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3761 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3885 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4097 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4129 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4185 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4507 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4563 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4565 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4601 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4613 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4619 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4621 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4633 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4657 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4669 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4675 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4677 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4689 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4713 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4725 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4731 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4733 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4745 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4781 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4787 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4789 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4801 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4825 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4837 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4843 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4845 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4857 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4893 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4899 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4901 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4913 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4937 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4949 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4955 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4957 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4969 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4993 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5011 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5013 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5025 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5049 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5061 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5067 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5069 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5081 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5093 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5105 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5117 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5123 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5125 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5137 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5161 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5173 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5179 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5181 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5193 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5217 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5229 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5235 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5237 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5249 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5261 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5273 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5285 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5291 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5293 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5305 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5317 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5329 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5341 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5347 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5349 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5361 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5373 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5385 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5397 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5403 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5405 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5417 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5429 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5441 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5453 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5459 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5461 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5473 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5485 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5497 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5509 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5515 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5517 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5529 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5541 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5553 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5565 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5571 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5573 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5585 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5597 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5609 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5621 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5627 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5629 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5641 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5653 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5665 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5677 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5683 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5685 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5697 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5709 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5721 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1369 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1649 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1929 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2209 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2489 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2689 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2769 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2785 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3009 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3037 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3049 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3065 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3093 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3121 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3149 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3177 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3233 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3261 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3289 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3317 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3329 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3345 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3373 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3401 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3429 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3457 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3513 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3541 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3569 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3597 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3609 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3625 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3653 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3681 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3709 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3737 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3793 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3821 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3849 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3877 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3889 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3905 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3933 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3961 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3989 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4017 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4073 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4101 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4129 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4157 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4169 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4185 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4213 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4241 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4269 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4297 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4353 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4381 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4409 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4437 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4449 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4465 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4493 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4521 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4549 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4565 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4577 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4589 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4593 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4605 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4621 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4633 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4645 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4649 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4661 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4677 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4689 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4701 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4705 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4717 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4729 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4733 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4745 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4757 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4761 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4773 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4789 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4801 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4813 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4817 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4829 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4845 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4857 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4869 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4873 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4885 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4901 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4913 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4925 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4929 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4941 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4957 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4969 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4981 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4985 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4997 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5009 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5013 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5025 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5037 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5041 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5053 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5069 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5081 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5093 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5097 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5109 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5137 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5149 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5153 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5165 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5177 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5193 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5205 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5209 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5221 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5233 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5249 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5261 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5265 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5277 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5289 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5293 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5305 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5317 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5321 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5333 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5345 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5361 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5373 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5377 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5389 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5401 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5417 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5429 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5433 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5445 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5457 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5473 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5485 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5489 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5501 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5513 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5529 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5541 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5545 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5557 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5569 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5585 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5597 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5601 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5613 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5625 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5641 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5653 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5657 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5669 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5681 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_5709 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5713 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_5725 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_993 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__clkbuf_2 _00_ (.A(buf_in[19]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 _01_ (.A(buf_in[20]),
    .X(net89));
 sky130_fd_sc_hd__buf_2 _02_ (.A(net162),
    .X(buf_out[21]));
 sky130_fd_sc_hd__clkbuf_1 _03_ (.A(buf_in[22]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 _04_ (.A(buf_in[23]),
    .X(net83));
 sky130_fd_sc_hd__buf_2 _05_ (.A(net159),
    .X(buf_out[24]));
 sky130_fd_sc_hd__clkbuf_1 _06_ (.A(buf_in[25]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _07_ (.A(buf_in[26]),
    .X(net77));
 sky130_fd_sc_hd__buf_2 _08_ (.A(net157),
    .X(buf_out[27]));
 sky130_fd_sc_hd__clkbuf_4 _09_ (.A(buf_in[28]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_4 _10_ (.A(buf_in[29]),
    .X(net73));
 sky130_fd_sc_hd__buf_2 _11_ (.A(net155),
    .X(buf_out[30]));
 sky130_fd_sc_hd__clkbuf_4 _12_ (.A(buf_in[31]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_4 _13_ (.A(buf_in[32]),
    .X(net69));
 sky130_fd_sc_hd__buf_2 _14_ (.A(net153),
    .X(buf_out[33]));
 sky130_fd_sc_hd__clkbuf_4 _15_ (.A(buf_in[34]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 _16_ (.A(net152),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 _17_ (.A(net150),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 _18_ (.A(net149),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 _19_ (.A(net148),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 _20_ (.A(net146),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 _21_ (.A(net142),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_4 _22_ (.A(net141),
    .X(net55));
 sky130_fd_sc_hd__buf_2 _23_ (.A(net174),
    .X(buf_out[0]));
 sky130_fd_sc_hd__buf_2 _24_ (.A(buf_in[1]),
    .X(net52));
 sky130_fd_sc_hd__buf_2 _25_ (.A(buf_in[2]),
    .X(net49));
 sky130_fd_sc_hd__buf_2 _26_ (.A(net143),
    .X(buf_out[3]));
 sky130_fd_sc_hd__clkbuf_2 _27_ (.A(buf_in[4]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 _28_ (.A(buf_in[5]),
    .X(net43));
 sky130_fd_sc_hd__buf_2 _29_ (.A(net138),
    .X(buf_out[6]));
 sky130_fd_sc_hd__clkbuf_2 _30_ (.A(buf_in[7]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 _31_ (.A(buf_in[8]),
    .X(net37));
 sky130_fd_sc_hd__buf_2 _32_ (.A(net135),
    .X(buf_out[9]));
 sky130_fd_sc_hd__clkbuf_2 _33_ (.A(buf_in[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 _34_ (.A(buf_in[11]),
    .X(net31));
 sky130_fd_sc_hd__buf_2 _35_ (.A(net171),
    .X(buf_out[12]));
 sky130_fd_sc_hd__clkbuf_2 _36_ (.A(buf_in[13]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 _37_ (.A(buf_in[14]),
    .X(net25));
 sky130_fd_sc_hd__buf_2 _38_ (.A(net168),
    .X(buf_out[15]));
 sky130_fd_sc_hd__clkbuf_2 _39_ (.A(buf_in[16]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 _40_ (.A(buf_in[17]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 _41_ (.A(net165),
    .X(buf_out[18]));
 sky130_fd_sc_hd__buf_2 \u_rp[0].u_buf  (.A(net131),
    .X(ch_out[0]));
 sky130_fd_sc_hd__buf_2 \u_rp[10].u_buf  (.A(net128),
    .X(ch_out[10]));
 sky130_fd_sc_hd__clkbuf_1 \u_rp[11].u_buf  (.A(ch_in[11]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 \u_rp[12].u_buf  (.A(net126),
    .X(ch_out[12]));
 sky130_fd_sc_hd__buf_2 \u_rp[13].u_buf  (.A(net124),
    .X(ch_out[13]));
 sky130_fd_sc_hd__buf_2 \u_rp[14].u_buf  (.A(ch_in[14]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 \u_rp[15].u_buf  (.A(net122),
    .X(ch_out[15]));
 sky130_fd_sc_hd__buf_2 \u_rp[16].u_buf  (.A(net120),
    .X(ch_out[16]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[17].u_buf  (.A(ch_in[17]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 \u_rp[18].u_buf  (.A(net119),
    .X(ch_out[18]));
 sky130_fd_sc_hd__buf_2 \u_rp[19].u_buf  (.A(net118),
    .X(ch_out[19]));
 sky130_fd_sc_hd__buf_2 \u_rp[1].u_buf  (.A(net114),
    .X(ch_out[1]));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[20].u_buf  (.A(ch_in[20]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 \u_rp[21].u_buf  (.A(net113),
    .X(ch_out[21]));
 sky130_fd_sc_hd__buf_2 \u_rp[22].u_buf  (.A(net112),
    .X(ch_out[22]));
 sky130_fd_sc_hd__buf_2 \u_rp[23].u_buf  (.A(ch_in[23]),
    .X(ch_out[23]));
 sky130_fd_sc_hd__buf_2 \u_rp[24].u_buf  (.A(ch_in[24]),
    .X(ch_out[24]));
 sky130_fd_sc_hd__buf_2 \u_rp[25].u_buf  (.A(ch_in[25]),
    .X(ch_out[25]));
 sky130_fd_sc_hd__buf_2 \u_rp[26].u_buf  (.A(ch_in[26]),
    .X(ch_out[26]));
 sky130_fd_sc_hd__buf_2 \u_rp[2].u_buf  (.A(ch_in[2]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 \u_rp[3].u_buf  (.A(net108),
    .X(ch_out[3]));
 sky130_fd_sc_hd__buf_2 \u_rp[4].u_buf  (.A(net104),
    .X(ch_out[4]));
 sky130_fd_sc_hd__clkbuf_1 \u_rp[5].u_buf  (.A(ch_in[5]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 \u_rp[6].u_buf  (.A(net101),
    .X(ch_out[6]));
 sky130_fd_sc_hd__buf_2 \u_rp[7].u_buf  (.A(net98),
    .X(ch_out[7]));
 sky130_fd_sc_hd__buf_2 \u_rp[8].u_buf  (.A(ch_in[8]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 \u_rp[9].u_buf  (.A(net95),
    .X(ch_out[9]));
 sky130_fd_sc_hd__buf_6 wire1 (.A(net2),
    .X(ch_out[8]));
 sky130_fd_sc_hd__buf_6 wire10 (.A(net11),
    .X(net10));
 sky130_fd_sc_hd__buf_6 wire100 (.A(ch_in[7]),
    .X(net100));
 sky130_fd_sc_hd__buf_6 wire101 (.A(net102),
    .X(net101));
 sky130_fd_sc_hd__buf_6 wire102 (.A(net103),
    .X(net102));
 sky130_fd_sc_hd__buf_6 wire103 (.A(ch_in[6]),
    .X(net103));
 sky130_fd_sc_hd__buf_12 wire104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__buf_8 wire105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__buf_6 wire106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__buf_4 wire107 (.A(ch_in[4]),
    .X(net107));
 sky130_fd_sc_hd__buf_12 wire108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__buf_8 wire109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__buf_6 wire11 (.A(net8),
    .X(net11));
 sky130_fd_sc_hd__buf_6 wire110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__buf_4 wire111 (.A(ch_in[3]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_4 wire112 (.A(ch_in[22]),
    .X(net112));
 sky130_fd_sc_hd__buf_4 wire113 (.A(ch_in[21]),
    .X(net113));
 sky130_fd_sc_hd__buf_12 wire114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__buf_8 wire115 (.A(net116),
    .X(net115));
 sky130_fd_sc_hd__buf_6 wire116 (.A(net117),
    .X(net116));
 sky130_fd_sc_hd__buf_6 wire117 (.A(ch_in[1]),
    .X(net117));
 sky130_fd_sc_hd__buf_6 wire118 (.A(ch_in[19]),
    .X(net118));
 sky130_fd_sc_hd__buf_6 wire119 (.A(ch_in[18]),
    .X(net119));
 sky130_fd_sc_hd__buf_4 wire12 (.A(net12),
    .X(ch_out[20]));
 sky130_fd_sc_hd__buf_6 wire120 (.A(net121),
    .X(net120));
 sky130_fd_sc_hd__buf_4 wire121 (.A(ch_in[16]),
    .X(net121));
 sky130_fd_sc_hd__buf_6 wire122 (.A(net123),
    .X(net122));
 sky130_fd_sc_hd__buf_4 wire123 (.A(ch_in[15]),
    .X(net123));
 sky130_fd_sc_hd__buf_6 wire124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__buf_6 wire125 (.A(ch_in[13]),
    .X(net125));
 sky130_fd_sc_hd__buf_6 wire126 (.A(net127),
    .X(net126));
 sky130_fd_sc_hd__buf_6 wire127 (.A(ch_in[12]),
    .X(net127));
 sky130_fd_sc_hd__buf_6 wire128 (.A(net129),
    .X(net128));
 sky130_fd_sc_hd__buf_6 wire129 (.A(net130),
    .X(net129));
 sky130_fd_sc_hd__buf_6 wire13 (.A(net13),
    .X(ch_out[17]));
 sky130_fd_sc_hd__buf_4 wire130 (.A(ch_in[10]),
    .X(net130));
 sky130_fd_sc_hd__buf_12 wire131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__buf_8 wire132 (.A(net133),
    .X(net132));
 sky130_fd_sc_hd__buf_6 wire133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__buf_6 wire134 (.A(ch_in[0]),
    .X(net134));
 sky130_fd_sc_hd__buf_6 wire135 (.A(net136),
    .X(net135));
 sky130_fd_sc_hd__buf_6 wire136 (.A(net137),
    .X(net136));
 sky130_fd_sc_hd__buf_4 wire137 (.A(buf_in[9]),
    .X(net137));
 sky130_fd_sc_hd__buf_6 wire138 (.A(net139),
    .X(net138));
 sky130_fd_sc_hd__buf_6 wire139 (.A(net140),
    .X(net139));
 sky130_fd_sc_hd__buf_6 wire14 (.A(net15),
    .X(ch_out[14]));
 sky130_fd_sc_hd__buf_4 wire140 (.A(buf_in[6]),
    .X(net140));
 sky130_fd_sc_hd__buf_4 wire141 (.A(buf_in[41]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_4 wire142 (.A(buf_in[40]),
    .X(net142));
 sky130_fd_sc_hd__buf_6 wire143 (.A(net144),
    .X(net143));
 sky130_fd_sc_hd__buf_6 wire144 (.A(net145),
    .X(net144));
 sky130_fd_sc_hd__buf_6 wire145 (.A(buf_in[3]),
    .X(net145));
 sky130_fd_sc_hd__buf_6 wire146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__buf_6 wire147 (.A(buf_in[39]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 wire148 (.A(buf_in[38]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_4 wire149 (.A(buf_in[37]),
    .X(net149));
 sky130_fd_sc_hd__buf_6 wire15 (.A(net14),
    .X(net15));
 sky130_fd_sc_hd__buf_6 wire150 (.A(net151),
    .X(net150));
 sky130_fd_sc_hd__buf_6 wire151 (.A(buf_in[36]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_4 wire152 (.A(buf_in[35]),
    .X(net152));
 sky130_fd_sc_hd__buf_6 wire153 (.A(net154),
    .X(net153));
 sky130_fd_sc_hd__buf_6 wire154 (.A(buf_in[33]),
    .X(net154));
 sky130_fd_sc_hd__buf_6 wire155 (.A(net156),
    .X(net155));
 sky130_fd_sc_hd__buf_6 wire156 (.A(buf_in[30]),
    .X(net156));
 sky130_fd_sc_hd__buf_6 wire157 (.A(net158),
    .X(net157));
 sky130_fd_sc_hd__buf_6 wire158 (.A(buf_in[27]),
    .X(net158));
 sky130_fd_sc_hd__buf_6 wire159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__buf_6 wire16 (.A(net17),
    .X(ch_out[11]));
 sky130_fd_sc_hd__buf_6 wire160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__buf_4 wire161 (.A(buf_in[24]),
    .X(net161));
 sky130_fd_sc_hd__buf_6 wire162 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__buf_6 wire163 (.A(net164),
    .X(net163));
 sky130_fd_sc_hd__buf_4 wire164 (.A(buf_in[21]),
    .X(net164));
 sky130_fd_sc_hd__buf_6 wire165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__buf_6 wire166 (.A(net167),
    .X(net166));
 sky130_fd_sc_hd__buf_4 wire167 (.A(buf_in[18]),
    .X(net167));
 sky130_fd_sc_hd__buf_6 wire168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__buf_6 wire169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__buf_6 wire17 (.A(net18),
    .X(net17));
 sky130_fd_sc_hd__buf_4 wire170 (.A(buf_in[15]),
    .X(net170));
 sky130_fd_sc_hd__buf_6 wire171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__buf_6 wire172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__buf_4 wire173 (.A(buf_in[12]),
    .X(net173));
 sky130_fd_sc_hd__buf_6 wire174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__buf_6 wire175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__buf_6 wire176 (.A(buf_in[0]),
    .X(net176));
 sky130_fd_sc_hd__buf_4 wire18 (.A(net16),
    .X(net18));
 sky130_fd_sc_hd__buf_6 wire19 (.A(net20),
    .X(buf_out[17]));
 sky130_fd_sc_hd__buf_6 wire2 (.A(net3),
    .X(net2));
 sky130_fd_sc_hd__buf_6 wire20 (.A(net21),
    .X(net20));
 sky130_fd_sc_hd__buf_4 wire21 (.A(net19),
    .X(net21));
 sky130_fd_sc_hd__buf_6 wire22 (.A(net23),
    .X(buf_out[16]));
 sky130_fd_sc_hd__buf_6 wire23 (.A(net24),
    .X(net23));
 sky130_fd_sc_hd__buf_4 wire24 (.A(net22),
    .X(net24));
 sky130_fd_sc_hd__buf_6 wire25 (.A(net26),
    .X(buf_out[14]));
 sky130_fd_sc_hd__buf_6 wire26 (.A(net27),
    .X(net26));
 sky130_fd_sc_hd__buf_4 wire27 (.A(net25),
    .X(net27));
 sky130_fd_sc_hd__buf_6 wire28 (.A(net29),
    .X(buf_out[13]));
 sky130_fd_sc_hd__buf_6 wire29 (.A(net30),
    .X(net29));
 sky130_fd_sc_hd__buf_6 wire3 (.A(net1),
    .X(net3));
 sky130_fd_sc_hd__buf_4 wire30 (.A(net28),
    .X(net30));
 sky130_fd_sc_hd__buf_6 wire31 (.A(net32),
    .X(buf_out[11]));
 sky130_fd_sc_hd__buf_6 wire32 (.A(net33),
    .X(net32));
 sky130_fd_sc_hd__buf_4 wire33 (.A(net31),
    .X(net33));
 sky130_fd_sc_hd__buf_6 wire34 (.A(net35),
    .X(buf_out[10]));
 sky130_fd_sc_hd__buf_6 wire35 (.A(net36),
    .X(net35));
 sky130_fd_sc_hd__buf_4 wire36 (.A(net34),
    .X(net36));
 sky130_fd_sc_hd__buf_6 wire37 (.A(net38),
    .X(buf_out[8]));
 sky130_fd_sc_hd__buf_6 wire38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__buf_4 wire39 (.A(net37),
    .X(net39));
 sky130_fd_sc_hd__buf_6 wire4 (.A(net5),
    .X(ch_out[5]));
 sky130_fd_sc_hd__buf_6 wire40 (.A(net41),
    .X(buf_out[7]));
 sky130_fd_sc_hd__buf_6 wire41 (.A(net42),
    .X(net41));
 sky130_fd_sc_hd__buf_4 wire42 (.A(net40),
    .X(net42));
 sky130_fd_sc_hd__buf_6 wire43 (.A(net44),
    .X(buf_out[5]));
 sky130_fd_sc_hd__buf_6 wire44 (.A(net45),
    .X(net44));
 sky130_fd_sc_hd__buf_4 wire45 (.A(net43),
    .X(net45));
 sky130_fd_sc_hd__buf_6 wire46 (.A(net47),
    .X(buf_out[4]));
 sky130_fd_sc_hd__buf_6 wire47 (.A(net48),
    .X(net47));
 sky130_fd_sc_hd__buf_4 wire48 (.A(net46),
    .X(net48));
 sky130_fd_sc_hd__buf_6 wire49 (.A(net50),
    .X(buf_out[2]));
 sky130_fd_sc_hd__buf_6 wire5 (.A(net6),
    .X(net5));
 sky130_fd_sc_hd__buf_6 wire50 (.A(net51),
    .X(net50));
 sky130_fd_sc_hd__buf_6 wire51 (.A(net49),
    .X(net51));
 sky130_fd_sc_hd__buf_6 wire52 (.A(net53),
    .X(buf_out[1]));
 sky130_fd_sc_hd__buf_6 wire53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__buf_6 wire54 (.A(net52),
    .X(net54));
 sky130_fd_sc_hd__buf_4 wire55 (.A(net56),
    .X(buf_out[41]));
 sky130_fd_sc_hd__buf_6 wire56 (.A(net55),
    .X(net56));
 sky130_fd_sc_hd__buf_4 wire57 (.A(net58),
    .X(buf_out[40]));
 sky130_fd_sc_hd__buf_6 wire58 (.A(net57),
    .X(net58));
 sky130_fd_sc_hd__buf_2 wire59 (.A(net59),
    .X(buf_out[39]));
 sky130_fd_sc_hd__buf_6 wire6 (.A(net7),
    .X(net6));
 sky130_fd_sc_hd__buf_4 wire60 (.A(net61),
    .X(buf_out[38]));
 sky130_fd_sc_hd__buf_6 wire61 (.A(net60),
    .X(net61));
 sky130_fd_sc_hd__buf_6 wire62 (.A(net63),
    .X(buf_out[37]));
 sky130_fd_sc_hd__buf_6 wire63 (.A(net62),
    .X(net63));
 sky130_fd_sc_hd__buf_2 wire64 (.A(net64),
    .X(buf_out[36]));
 sky130_fd_sc_hd__buf_6 wire65 (.A(net66),
    .X(buf_out[35]));
 sky130_fd_sc_hd__buf_6 wire66 (.A(net65),
    .X(net66));
 sky130_fd_sc_hd__buf_6 wire67 (.A(net68),
    .X(buf_out[34]));
 sky130_fd_sc_hd__buf_6 wire68 (.A(net67),
    .X(net68));
 sky130_fd_sc_hd__buf_6 wire69 (.A(net70),
    .X(buf_out[32]));
 sky130_fd_sc_hd__buf_4 wire7 (.A(net4),
    .X(net7));
 sky130_fd_sc_hd__buf_6 wire70 (.A(net69),
    .X(net70));
 sky130_fd_sc_hd__buf_6 wire71 (.A(net72),
    .X(buf_out[31]));
 sky130_fd_sc_hd__buf_6 wire72 (.A(net71),
    .X(net72));
 sky130_fd_sc_hd__buf_6 wire73 (.A(net74),
    .X(buf_out[29]));
 sky130_fd_sc_hd__buf_6 wire74 (.A(net73),
    .X(net74));
 sky130_fd_sc_hd__buf_6 wire75 (.A(net76),
    .X(buf_out[28]));
 sky130_fd_sc_hd__buf_6 wire76 (.A(net75),
    .X(net76));
 sky130_fd_sc_hd__buf_6 wire77 (.A(net78),
    .X(buf_out[26]));
 sky130_fd_sc_hd__buf_6 wire78 (.A(net79),
    .X(net78));
 sky130_fd_sc_hd__buf_4 wire79 (.A(net77),
    .X(net79));
 sky130_fd_sc_hd__buf_6 wire8 (.A(net9),
    .X(ch_out[2]));
 sky130_fd_sc_hd__buf_6 wire80 (.A(net81),
    .X(buf_out[25]));
 sky130_fd_sc_hd__buf_6 wire81 (.A(net82),
    .X(net81));
 sky130_fd_sc_hd__buf_4 wire82 (.A(net80),
    .X(net82));
 sky130_fd_sc_hd__buf_6 wire83 (.A(net84),
    .X(buf_out[23]));
 sky130_fd_sc_hd__buf_6 wire84 (.A(net85),
    .X(net84));
 sky130_fd_sc_hd__buf_4 wire85 (.A(net83),
    .X(net85));
 sky130_fd_sc_hd__buf_6 wire86 (.A(net87),
    .X(buf_out[22]));
 sky130_fd_sc_hd__buf_6 wire87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__buf_4 wire88 (.A(net86),
    .X(net88));
 sky130_fd_sc_hd__buf_6 wire89 (.A(net90),
    .X(buf_out[20]));
 sky130_fd_sc_hd__buf_6 wire9 (.A(net10),
    .X(net9));
 sky130_fd_sc_hd__buf_6 wire90 (.A(net91),
    .X(net90));
 sky130_fd_sc_hd__buf_4 wire91 (.A(net89),
    .X(net91));
 sky130_fd_sc_hd__buf_6 wire92 (.A(net93),
    .X(buf_out[19]));
 sky130_fd_sc_hd__buf_6 wire93 (.A(net94),
    .X(net93));
 sky130_fd_sc_hd__buf_4 wire94 (.A(net92),
    .X(net94));
 sky130_fd_sc_hd__buf_6 wire95 (.A(net96),
    .X(net95));
 sky130_fd_sc_hd__buf_6 wire96 (.A(net97),
    .X(net96));
 sky130_fd_sc_hd__buf_4 wire97 (.A(ch_in[9]),
    .X(net97));
 sky130_fd_sc_hd__buf_6 wire98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__buf_6 wire99 (.A(net100),
    .X(net99));
endmodule

