magic
tech sky130A
magscale 1 2
timestamp 1698825822
<< obsli1 >>
rect 1104 2159 528816 9809
<< metal1 >>
rect 200062 11200 200118 12000
rect 200606 11200 200662 12000
rect 201150 11200 201206 12000
rect 201694 11200 201750 12000
rect 202238 11200 202294 12000
rect 202782 11200 202838 12000
rect 203326 11200 203382 12000
rect 203870 11200 203926 12000
rect 204414 11200 204470 12000
rect 204958 11200 205014 12000
rect 205502 11200 205558 12000
rect 206046 11200 206102 12000
rect 206590 11200 206646 12000
rect 207134 11200 207190 12000
rect 207678 11200 207734 12000
rect 208222 11200 208278 12000
rect 208766 11200 208822 12000
rect 209310 11200 209366 12000
rect 209854 11200 209910 12000
rect 210398 11200 210454 12000
rect 210942 11200 210998 12000
rect 211486 11200 211542 12000
rect 212030 11200 212086 12000
rect 212574 11200 212630 12000
rect 213118 11200 213174 12000
rect 213662 11200 213718 12000
rect 214206 11200 214262 12000
rect 214750 11200 214806 12000
rect 215294 11200 215350 12000
rect 215838 11200 215894 12000
rect 216382 11200 216438 12000
rect 216926 11200 216982 12000
rect 217470 11200 217526 12000
rect 218014 11200 218070 12000
rect 218558 11200 218614 12000
rect 219102 11200 219158 12000
rect 219646 11200 219702 12000
rect 220190 11200 220246 12000
rect 220734 11200 220790 12000
rect 221278 11200 221334 12000
rect 221822 11200 221878 12000
rect 222366 11200 222422 12000
rect 222910 11200 222966 12000
rect 223454 11200 223510 12000
rect 223998 11200 224054 12000
rect 224542 11200 224598 12000
rect 225086 11200 225142 12000
rect 225630 11200 225686 12000
rect 226174 11200 226230 12000
rect 226718 11200 226774 12000
rect 227262 11200 227318 12000
rect 227806 11200 227862 12000
rect 228350 11200 228406 12000
rect 228894 11200 228950 12000
rect 229438 11200 229494 12000
rect 229982 11200 230038 12000
rect 230526 11200 230582 12000
rect 231070 11200 231126 12000
rect 231614 11200 231670 12000
rect 232158 11200 232214 12000
rect 232702 11200 232758 12000
rect 233246 11200 233302 12000
rect 233790 11200 233846 12000
rect 234334 11200 234390 12000
rect 234878 11200 234934 12000
rect 235422 11200 235478 12000
rect 235966 11200 236022 12000
rect 236510 11200 236566 12000
rect 237054 11200 237110 12000
rect 237598 11200 237654 12000
rect 238142 11200 238198 12000
rect 238686 11200 238742 12000
rect 239230 11200 239286 12000
rect 239774 11200 239830 12000
rect 240318 11200 240374 12000
rect 240862 11200 240918 12000
rect 241406 11200 241462 12000
rect 241950 11200 242006 12000
rect 242494 11200 242550 12000
rect 243038 11200 243094 12000
rect 243582 11200 243638 12000
rect 244126 11172 244182 12000
rect 244670 11200 244726 12000
rect 245214 11200 245270 12000
rect 245758 11200 245814 12000
rect 246302 11200 246358 12000
rect 246846 11200 246902 12000
rect 247390 11200 247446 12000
rect 247934 11200 247990 12000
rect 248478 11200 248534 12000
rect 249022 11200 249078 12000
rect 249566 11200 249622 12000
rect 250110 11200 250166 12000
rect 250654 11200 250710 12000
rect 251198 11200 251254 12000
rect 251742 11200 251798 12000
rect 252286 11200 252342 12000
rect 252830 11200 252886 12000
rect 253374 11200 253430 12000
rect 253918 11200 253974 12000
rect 254462 11200 254518 12000
rect 255006 11200 255062 12000
rect 255550 11200 255606 12000
rect 256094 11200 256150 12000
rect 256638 11200 256694 12000
rect 257182 11200 257238 12000
rect 360066 11200 360122 12000
rect 360610 11200 360666 12000
rect 361154 11200 361210 12000
rect 361698 11200 361754 12000
rect 362242 11200 362298 12000
rect 362786 11200 362842 12000
rect 363330 11200 363386 12000
rect 363874 11200 363930 12000
rect 364418 11200 364474 12000
rect 364962 11200 365018 12000
rect 365506 11200 365562 12000
rect 366050 11200 366106 12000
rect 366594 11200 366650 12000
rect 367138 11200 367194 12000
rect 367682 11200 367738 12000
rect 368226 11200 368282 12000
rect 368770 11200 368826 12000
rect 369314 11200 369370 12000
rect 369858 11200 369914 12000
rect 370402 11200 370458 12000
rect 370946 11200 371002 12000
rect 371490 11200 371546 12000
rect 372034 11200 372090 12000
rect 372578 11200 372634 12000
rect 373122 11200 373178 12000
rect 373666 11200 373722 12000
rect 374210 11200 374266 12000
rect 374754 11200 374810 12000
rect 375298 11200 375354 12000
rect 375842 11200 375898 12000
rect 376386 11200 376442 12000
rect 376930 11200 376986 12000
rect 377474 11200 377530 12000
rect 378018 11200 378074 12000
rect 378562 11200 378618 12000
rect 379106 11200 379162 12000
rect 379650 11200 379706 12000
rect 380194 11200 380250 12000
rect 380738 11200 380794 12000
rect 381282 11200 381338 12000
rect 381826 11200 381882 12000
rect 382370 11200 382426 12000
rect 382914 11200 382970 12000
rect 383458 11200 383514 12000
rect 384002 11200 384058 12000
rect 384546 11172 384602 12000
rect 385090 11200 385146 12000
rect 385634 11200 385690 12000
rect 386178 11200 386234 12000
rect 386722 11200 386778 12000
rect 387266 11200 387322 12000
rect 387810 11200 387866 12000
rect 388354 11200 388410 12000
rect 388898 11200 388954 12000
rect 389442 11200 389498 12000
rect 389986 11200 390042 12000
rect 390530 11200 390586 12000
rect 391074 11200 391130 12000
rect 391618 11200 391674 12000
rect 392162 11200 392218 12000
rect 392706 11200 392762 12000
rect 393250 11200 393306 12000
rect 393794 11200 393850 12000
rect 394338 11200 394394 12000
rect 394882 11200 394938 12000
rect 395426 11200 395482 12000
rect 395970 11200 396026 12000
rect 396514 11200 396570 12000
rect 397058 11172 397114 12000
rect 397602 11200 397658 12000
rect 398146 11200 398202 12000
rect 398690 11200 398746 12000
rect 399234 11200 399290 12000
rect 399778 11200 399834 12000
rect 400322 11200 400378 12000
rect 400866 11200 400922 12000
rect 401410 11200 401466 12000
rect 401954 11200 402010 12000
rect 402498 11200 402554 12000
rect 403042 11200 403098 12000
rect 403586 11200 403642 12000
rect 404130 11200 404186 12000
rect 440034 11200 440090 12000
rect 440306 11200 440362 12000
rect 440578 11200 440634 12000
rect 440850 11200 440906 12000
rect 441122 11200 441178 12000
rect 441394 11200 441450 12000
rect 441666 11200 441722 12000
rect 441938 11200 441994 12000
rect 442210 11200 442266 12000
rect 442482 11200 442538 12000
rect 442754 11172 442810 12000
rect 443026 11200 443082 12000
rect 443298 11200 443354 12000
rect 443570 11200 443626 12000
rect 443842 11200 443898 12000
rect 444114 11200 444170 12000
rect 444386 11200 444442 12000
rect 444658 11200 444714 12000
rect 444930 11200 444986 12000
rect 445202 11200 445258 12000
rect 445474 11200 445530 12000
rect 445746 11200 445802 12000
rect 446018 11200 446074 12000
rect 446290 11200 446346 12000
rect 446562 11200 446618 12000
rect 446834 11200 446890 12000
rect 447106 11172 447162 12000
rect 447378 11200 447434 12000
rect 447650 11200 447706 12000
rect 447922 11200 447978 12000
rect 448194 11200 448250 12000
rect 448466 11200 448522 12000
rect 480018 11200 480074 12000
rect 480290 11172 480346 12000
rect 480562 11200 480618 12000
rect 480834 11200 480890 12000
rect 481106 11200 481162 12000
rect 481378 11200 481434 12000
rect 481650 11200 481706 12000
rect 481922 11200 481978 12000
rect 482194 11200 482250 12000
rect 482466 11200 482522 12000
rect 482738 11200 482794 12000
rect 483010 11172 483066 12000
rect 483282 11200 483338 12000
rect 483554 11200 483610 12000
rect 483826 11200 483882 12000
rect 484098 11200 484154 12000
rect 484370 11200 484426 12000
rect 484642 11200 484698 12000
rect 484914 11200 484970 12000
rect 485186 11200 485242 12000
rect 485458 11200 485514 12000
rect 485730 11200 485786 12000
rect 486002 11200 486058 12000
rect 486274 11200 486330 12000
rect 486546 11200 486602 12000
rect 486818 11200 486874 12000
rect 487090 11200 487146 12000
rect 487362 11200 487418 12000
rect 487634 11200 487690 12000
rect 487906 11200 487962 12000
rect 488178 11200 488234 12000
rect 488450 11200 488506 12000
rect 488722 11200 488778 12000
rect 74 0 130 800
rect 1162 0 1218 800
rect 2250 0 2306 800
rect 3338 0 3394 800
rect 4426 0 4482 800
rect 5514 0 5570 800
rect 6602 0 6658 800
rect 7690 0 7746 800
rect 8778 0 8834 800
rect 9866 0 9922 800
rect 10954 0 11010 800
rect 12042 0 12098 800
rect 13130 0 13186 800
rect 14218 0 14274 800
rect 15306 0 15362 800
rect 16394 0 16450 800
rect 17482 0 17538 800
rect 18570 0 18626 800
rect 19658 0 19714 800
rect 20746 0 20802 800
rect 21834 0 21890 800
rect 22922 0 22978 800
rect 24010 0 24066 800
rect 25098 0 25154 800
rect 26186 0 26242 800
rect 27274 0 27330 800
rect 28362 0 28418 800
rect 29450 0 29506 800
rect 30538 0 30594 800
rect 31626 0 31682 800
rect 32714 0 32770 800
rect 33802 0 33858 800
rect 34890 0 34946 800
rect 35978 0 36034 800
rect 37066 0 37122 800
rect 38154 0 38210 800
rect 39242 0 39298 800
rect 40330 0 40386 800
rect 41418 0 41474 800
rect 42506 0 42562 800
rect 43594 0 43650 800
rect 44682 0 44738 800
rect 45770 0 45826 800
rect 46858 0 46914 800
rect 47946 0 48002 800
rect 49034 0 49090 800
rect 50122 0 50178 800
rect 51210 0 51266 800
rect 52298 0 52354 800
rect 53386 0 53442 800
rect 54474 0 54530 800
rect 55562 0 55618 800
rect 56650 0 56706 800
rect 57738 0 57794 800
rect 58826 0 58882 800
rect 59914 0 59970 800
rect 61002 0 61058 800
rect 62090 0 62146 800
rect 63178 0 63234 800
rect 64266 0 64322 800
rect 65354 0 65410 800
rect 66442 0 66498 800
rect 67530 0 67586 800
rect 68618 0 68674 800
rect 69706 0 69762 800
rect 70794 0 70850 800
rect 71882 0 71938 800
rect 72970 0 73026 800
rect 74058 0 74114 800
rect 75146 0 75202 800
rect 76234 0 76290 800
rect 77322 0 77378 800
rect 78410 0 78466 800
rect 79498 0 79554 800
rect 80586 0 80642 800
rect 81674 0 81730 800
rect 82762 0 82818 800
rect 83850 0 83906 800
rect 84938 0 84994 800
rect 86026 0 86082 800
rect 87114 0 87170 800
rect 88202 0 88258 800
rect 89290 0 89346 800
rect 90378 0 90434 800
rect 91466 0 91522 800
rect 92554 0 92610 800
rect 93642 0 93698 800
rect 94730 0 94786 800
rect 95818 0 95874 800
rect 96906 0 96962 800
rect 97994 0 98050 800
rect 99082 0 99138 800
rect 100170 0 100226 800
rect 101258 0 101314 800
rect 102346 0 102402 800
rect 103434 0 103490 800
rect 104522 0 104578 800
rect 105610 0 105666 800
rect 106698 0 106754 800
rect 107786 0 107842 800
rect 108874 0 108930 800
rect 109962 0 110018 800
rect 111050 0 111106 800
rect 112138 0 112194 800
rect 113226 0 113282 800
rect 114314 0 114370 800
rect 120026 0 120082 800
rect 122202 0 122258 800
rect 124378 0 124434 800
rect 126554 0 126610 800
rect 128730 0 128786 800
rect 130906 0 130962 800
rect 133082 0 133138 800
rect 135258 0 135314 800
rect 137434 0 137490 800
rect 139610 0 139666 800
rect 141786 0 141842 800
rect 143962 0 144018 800
rect 146138 0 146194 800
rect 148314 0 148370 800
rect 150490 0 150546 800
rect 152666 0 152722 800
rect 154842 0 154898 800
rect 157018 0 157074 800
rect 159194 0 159250 800
rect 161370 0 161426 800
rect 162050 0 162106 800
rect 164226 0 164282 800
rect 166402 0 166458 800
rect 168578 0 168634 800
rect 170754 0 170810 800
rect 172930 0 172986 800
rect 175106 0 175162 800
rect 177282 0 177338 800
rect 179458 0 179514 800
rect 181634 0 181690 800
rect 183810 0 183866 800
rect 185986 0 186042 800
rect 188162 0 188218 800
rect 190338 0 190394 800
rect 192514 0 192570 800
rect 194690 0 194746 800
rect 220054 0 220110 800
rect 222230 0 222286 800
rect 224406 0 224462 800
rect 226582 0 226638 800
rect 228758 0 228814 800
rect 230934 0 230990 800
rect 233110 0 233166 800
rect 235286 0 235342 800
rect 237462 0 237518 800
rect 239638 0 239694 800
rect 241814 0 241870 800
rect 243990 0 244046 800
rect 246166 0 246222 800
rect 248342 0 248398 800
rect 250518 0 250574 800
rect 252694 0 252750 800
rect 254870 0 254926 800
rect 257046 0 257102 800
rect 259222 0 259278 800
rect 261398 0 261454 800
rect 263574 0 263630 800
rect 265750 0 265806 800
rect 267926 0 267982 800
rect 270102 0 270158 800
rect 272278 0 272334 800
rect 274454 0 274510 800
rect 276630 0 276686 800
rect 278806 0 278862 800
rect 280982 0 281038 800
rect 283158 0 283214 800
rect 285334 0 285390 800
rect 287510 0 287566 800
rect 289686 0 289742 800
rect 291862 0 291918 800
rect 294038 0 294094 800
rect 296214 0 296270 800
rect 298390 0 298446 800
rect 300566 0 300622 800
rect 302742 0 302798 800
rect 304918 0 304974 800
rect 307094 0 307150 800
rect 309270 0 309326 800
rect 311446 0 311502 800
rect 313622 0 313678 800
rect 315798 0 315854 800
rect 317974 0 318030 800
rect 360066 0 360122 800
rect 362242 0 362298 800
rect 364418 0 364474 800
rect 366594 0 366650 800
rect 368770 0 368826 800
rect 370946 0 371002 800
rect 373122 0 373178 800
rect 375298 0 375354 800
rect 377474 0 377530 800
rect 379650 0 379706 800
rect 381826 0 381882 800
rect 384002 0 384058 800
rect 386178 0 386234 800
rect 388354 0 388410 800
rect 390530 0 390586 800
rect 392706 0 392762 800
rect 394882 0 394938 800
rect 397058 0 397114 800
rect 399234 0 399290 800
rect 401410 0 401466 800
rect 403586 0 403642 800
rect 405762 0 405818 800
rect 407938 0 407994 800
rect 410114 0 410170 800
rect 412290 0 412346 800
rect 414466 0 414522 800
rect 416642 0 416698 800
rect 418818 0 418874 800
rect 420994 0 421050 800
rect 423170 0 423226 800
rect 425346 0 425402 800
rect 427522 0 427578 800
rect 429698 0 429754 800
rect 431874 0 431930 800
rect 434050 0 434106 800
rect 436226 0 436282 800
rect 438402 0 438458 800
rect 440578 0 440634 800
rect 442754 0 442810 800
rect 444930 0 444986 800
rect 447106 0 447162 800
rect 449282 0 449338 800
rect 451458 0 451514 800
rect 453634 0 453690 800
rect 455810 0 455866 800
rect 457986 0 458042 800
rect 460162 0 460218 800
rect 462338 0 462394 800
rect 464514 0 464570 800
rect 466690 0 466746 800
rect 468866 0 468922 800
rect 471042 0 471098 800
rect 473218 0 473274 800
rect 475394 0 475450 800
rect 477570 0 477626 800
rect 479746 0 479802 800
rect 481922 0 481978 800
rect 484098 0 484154 800
rect 486274 0 486330 800
rect 488450 0 488506 800
rect 490626 0 490682 800
rect 492802 0 492858 800
rect 494978 0 495034 800
rect 497154 0 497210 800
rect 499330 0 499386 800
<< obsm1 >>
rect 130 11144 200006 11960
rect 200174 11144 200550 11960
rect 200718 11144 201094 11960
rect 201262 11144 201638 11960
rect 201806 11144 202182 11960
rect 202350 11144 202726 11960
rect 202894 11144 203270 11960
rect 203438 11144 203814 11960
rect 203982 11144 204358 11960
rect 204526 11144 204902 11960
rect 205070 11144 205446 11960
rect 205614 11144 205990 11960
rect 206158 11144 206534 11960
rect 206702 11144 207078 11960
rect 207246 11144 207622 11960
rect 207790 11144 208166 11960
rect 208334 11144 208710 11960
rect 208878 11144 209254 11960
rect 209422 11144 209798 11960
rect 209966 11144 210342 11960
rect 210510 11144 210886 11960
rect 211054 11144 211430 11960
rect 211598 11144 211974 11960
rect 212142 11144 212518 11960
rect 212686 11144 213062 11960
rect 213230 11144 213606 11960
rect 213774 11144 214150 11960
rect 214318 11144 214694 11960
rect 214862 11144 215238 11960
rect 215406 11144 215782 11960
rect 215950 11144 216326 11960
rect 216494 11144 216870 11960
rect 217038 11144 217414 11960
rect 217582 11144 217958 11960
rect 218126 11144 218502 11960
rect 218670 11144 219046 11960
rect 219214 11144 219590 11960
rect 219758 11144 220134 11960
rect 220302 11144 220678 11960
rect 220846 11144 221222 11960
rect 221390 11144 221766 11960
rect 221934 11144 222310 11960
rect 222478 11144 222854 11960
rect 223022 11144 223398 11960
rect 223566 11144 223942 11960
rect 224110 11144 224486 11960
rect 224654 11144 225030 11960
rect 225198 11144 225574 11960
rect 225742 11144 226118 11960
rect 226286 11144 226662 11960
rect 226830 11144 227206 11960
rect 227374 11144 227750 11960
rect 227918 11144 228294 11960
rect 228462 11144 228838 11960
rect 229006 11144 229382 11960
rect 229550 11144 229926 11960
rect 230094 11144 230470 11960
rect 230638 11144 231014 11960
rect 231182 11144 231558 11960
rect 231726 11144 232102 11960
rect 232270 11144 232646 11960
rect 232814 11144 233190 11960
rect 233358 11144 233734 11960
rect 233902 11144 234278 11960
rect 234446 11144 234822 11960
rect 234990 11144 235366 11960
rect 235534 11144 235910 11960
rect 236078 11144 236454 11960
rect 236622 11144 236998 11960
rect 237166 11144 237542 11960
rect 237710 11144 238086 11960
rect 238254 11144 238630 11960
rect 238798 11144 239174 11960
rect 239342 11144 239718 11960
rect 239886 11144 240262 11960
rect 240430 11144 240806 11960
rect 240974 11144 241350 11960
rect 241518 11144 241894 11960
rect 242062 11144 242438 11960
rect 242606 11144 242982 11960
rect 243150 11144 243526 11960
rect 243694 11144 244070 11960
rect 130 11116 244070 11144
rect 244238 11144 244614 11960
rect 244782 11144 245158 11960
rect 245326 11144 245702 11960
rect 245870 11144 246246 11960
rect 246414 11144 246790 11960
rect 246958 11144 247334 11960
rect 247502 11144 247878 11960
rect 248046 11144 248422 11960
rect 248590 11144 248966 11960
rect 249134 11144 249510 11960
rect 249678 11144 250054 11960
rect 250222 11144 250598 11960
rect 250766 11144 251142 11960
rect 251310 11144 251686 11960
rect 251854 11144 252230 11960
rect 252398 11144 252774 11960
rect 252942 11144 253318 11960
rect 253486 11144 253862 11960
rect 254030 11144 254406 11960
rect 254574 11144 254950 11960
rect 255118 11144 255494 11960
rect 255662 11144 256038 11960
rect 256206 11144 256582 11960
rect 256750 11144 257126 11960
rect 257294 11144 360010 11960
rect 360178 11144 360554 11960
rect 360722 11144 361098 11960
rect 361266 11144 361642 11960
rect 361810 11144 362186 11960
rect 362354 11144 362730 11960
rect 362898 11144 363274 11960
rect 363442 11144 363818 11960
rect 363986 11144 364362 11960
rect 364530 11144 364906 11960
rect 365074 11144 365450 11960
rect 365618 11144 365994 11960
rect 366162 11144 366538 11960
rect 366706 11144 367082 11960
rect 367250 11144 367626 11960
rect 367794 11144 368170 11960
rect 368338 11144 368714 11960
rect 368882 11144 369258 11960
rect 369426 11144 369802 11960
rect 369970 11144 370346 11960
rect 370514 11144 370890 11960
rect 371058 11144 371434 11960
rect 371602 11144 371978 11960
rect 372146 11144 372522 11960
rect 372690 11144 373066 11960
rect 373234 11144 373610 11960
rect 373778 11144 374154 11960
rect 374322 11144 374698 11960
rect 374866 11144 375242 11960
rect 375410 11144 375786 11960
rect 375954 11144 376330 11960
rect 376498 11144 376874 11960
rect 377042 11144 377418 11960
rect 377586 11144 377962 11960
rect 378130 11144 378506 11960
rect 378674 11144 379050 11960
rect 379218 11144 379594 11960
rect 379762 11144 380138 11960
rect 380306 11144 380682 11960
rect 380850 11144 381226 11960
rect 381394 11144 381770 11960
rect 381938 11144 382314 11960
rect 382482 11144 382858 11960
rect 383026 11144 383402 11960
rect 383570 11144 383946 11960
rect 384114 11144 384490 11960
rect 244238 11116 384490 11144
rect 384658 11144 385034 11960
rect 385202 11144 385578 11960
rect 385746 11144 386122 11960
rect 386290 11144 386666 11960
rect 386834 11144 387210 11960
rect 387378 11144 387754 11960
rect 387922 11144 388298 11960
rect 388466 11144 388842 11960
rect 389010 11144 389386 11960
rect 389554 11144 389930 11960
rect 390098 11144 390474 11960
rect 390642 11144 391018 11960
rect 391186 11144 391562 11960
rect 391730 11144 392106 11960
rect 392274 11144 392650 11960
rect 392818 11144 393194 11960
rect 393362 11144 393738 11960
rect 393906 11144 394282 11960
rect 394450 11144 394826 11960
rect 394994 11144 395370 11960
rect 395538 11144 395914 11960
rect 396082 11144 396458 11960
rect 396626 11144 397002 11960
rect 384658 11116 397002 11144
rect 397170 11144 397546 11960
rect 397714 11144 398090 11960
rect 398258 11144 398634 11960
rect 398802 11144 399178 11960
rect 399346 11144 399722 11960
rect 399890 11144 400266 11960
rect 400434 11144 400810 11960
rect 400978 11144 401354 11960
rect 401522 11144 401898 11960
rect 402066 11144 402442 11960
rect 402610 11144 402986 11960
rect 403154 11144 403530 11960
rect 403698 11144 404074 11960
rect 404242 11144 439978 11960
rect 440146 11144 440250 11960
rect 440418 11144 440522 11960
rect 440690 11144 440794 11960
rect 440962 11144 441066 11960
rect 441234 11144 441338 11960
rect 441506 11144 441610 11960
rect 441778 11144 441882 11960
rect 442050 11144 442154 11960
rect 442322 11144 442426 11960
rect 442594 11144 442698 11960
rect 397170 11116 442698 11144
rect 442866 11144 442970 11960
rect 443138 11144 443242 11960
rect 443410 11144 443514 11960
rect 443682 11144 443786 11960
rect 443954 11144 444058 11960
rect 444226 11144 444330 11960
rect 444498 11144 444602 11960
rect 444770 11144 444874 11960
rect 445042 11144 445146 11960
rect 445314 11144 445418 11960
rect 445586 11144 445690 11960
rect 445858 11144 445962 11960
rect 446130 11144 446234 11960
rect 446402 11144 446506 11960
rect 446674 11144 446778 11960
rect 446946 11144 447050 11960
rect 442866 11116 447050 11144
rect 447218 11144 447322 11960
rect 447490 11144 447594 11960
rect 447762 11144 447866 11960
rect 448034 11144 448138 11960
rect 448306 11144 448410 11960
rect 448578 11144 479962 11960
rect 480130 11144 480234 11960
rect 447218 11116 480234 11144
rect 480402 11144 480506 11960
rect 480674 11144 480778 11960
rect 480946 11144 481050 11960
rect 481218 11144 481322 11960
rect 481490 11144 481594 11960
rect 481762 11144 481866 11960
rect 482034 11144 482138 11960
rect 482306 11144 482410 11960
rect 482578 11144 482682 11960
rect 482850 11144 482954 11960
rect 480402 11116 482954 11144
rect 483122 11144 483226 11960
rect 483394 11144 483498 11960
rect 483666 11144 483770 11960
rect 483938 11144 484042 11960
rect 484210 11144 484314 11960
rect 484482 11144 484586 11960
rect 484754 11144 484858 11960
rect 485026 11144 485130 11960
rect 485298 11144 485402 11960
rect 485570 11144 485674 11960
rect 485842 11144 485946 11960
rect 486114 11144 486218 11960
rect 486386 11144 486490 11960
rect 486658 11144 486762 11960
rect 486930 11144 487034 11960
rect 487202 11144 487306 11960
rect 487474 11144 487578 11960
rect 487746 11144 487850 11960
rect 488018 11144 488122 11960
rect 488290 11144 488394 11960
rect 488562 11144 488666 11960
rect 488834 11144 528816 11960
rect 483122 11116 528816 11144
rect 130 856 528816 11116
rect 186 8 1106 856
rect 1274 8 2194 856
rect 2362 8 3282 856
rect 3450 8 4370 856
rect 4538 8 5458 856
rect 5626 8 6546 856
rect 6714 8 7634 856
rect 7802 8 8722 856
rect 8890 8 9810 856
rect 9978 8 10898 856
rect 11066 8 11986 856
rect 12154 8 13074 856
rect 13242 8 14162 856
rect 14330 8 15250 856
rect 15418 8 16338 856
rect 16506 8 17426 856
rect 17594 8 18514 856
rect 18682 8 19602 856
rect 19770 8 20690 856
rect 20858 8 21778 856
rect 21946 8 22866 856
rect 23034 8 23954 856
rect 24122 8 25042 856
rect 25210 8 26130 856
rect 26298 8 27218 856
rect 27386 8 28306 856
rect 28474 8 29394 856
rect 29562 8 30482 856
rect 30650 8 31570 856
rect 31738 8 32658 856
rect 32826 8 33746 856
rect 33914 8 34834 856
rect 35002 8 35922 856
rect 36090 8 37010 856
rect 37178 8 38098 856
rect 38266 8 39186 856
rect 39354 8 40274 856
rect 40442 8 41362 856
rect 41530 8 42450 856
rect 42618 8 43538 856
rect 43706 8 44626 856
rect 44794 8 45714 856
rect 45882 8 46802 856
rect 46970 8 47890 856
rect 48058 8 48978 856
rect 49146 8 50066 856
rect 50234 8 51154 856
rect 51322 8 52242 856
rect 52410 8 53330 856
rect 53498 8 54418 856
rect 54586 8 55506 856
rect 55674 8 56594 856
rect 56762 8 57682 856
rect 57850 8 58770 856
rect 58938 8 59858 856
rect 60026 8 60946 856
rect 61114 8 62034 856
rect 62202 8 63122 856
rect 63290 8 64210 856
rect 64378 8 65298 856
rect 65466 8 66386 856
rect 66554 8 67474 856
rect 67642 8 68562 856
rect 68730 8 69650 856
rect 69818 8 70738 856
rect 70906 8 71826 856
rect 71994 8 72914 856
rect 73082 8 74002 856
rect 74170 8 75090 856
rect 75258 8 76178 856
rect 76346 8 77266 856
rect 77434 8 78354 856
rect 78522 8 79442 856
rect 79610 8 80530 856
rect 80698 8 81618 856
rect 81786 8 82706 856
rect 82874 8 83794 856
rect 83962 8 84882 856
rect 85050 8 85970 856
rect 86138 8 87058 856
rect 87226 8 88146 856
rect 88314 8 89234 856
rect 89402 8 90322 856
rect 90490 8 91410 856
rect 91578 8 92498 856
rect 92666 8 93586 856
rect 93754 8 94674 856
rect 94842 8 95762 856
rect 95930 8 96850 856
rect 97018 8 97938 856
rect 98106 8 99026 856
rect 99194 8 100114 856
rect 100282 8 101202 856
rect 101370 8 102290 856
rect 102458 8 103378 856
rect 103546 8 104466 856
rect 104634 8 105554 856
rect 105722 8 106642 856
rect 106810 8 107730 856
rect 107898 8 108818 856
rect 108986 8 109906 856
rect 110074 8 110994 856
rect 111162 8 112082 856
rect 112250 8 113170 856
rect 113338 8 114258 856
rect 114426 8 119970 856
rect 120138 8 122146 856
rect 122314 8 124322 856
rect 124490 8 126498 856
rect 126666 8 128674 856
rect 128842 8 130850 856
rect 131018 8 133026 856
rect 133194 8 135202 856
rect 135370 8 137378 856
rect 137546 8 139554 856
rect 139722 8 141730 856
rect 141898 8 143906 856
rect 144074 8 146082 856
rect 146250 8 148258 856
rect 148426 8 150434 856
rect 150602 8 152610 856
rect 152778 8 154786 856
rect 154954 8 156962 856
rect 157130 8 159138 856
rect 159306 8 161314 856
rect 161482 8 161994 856
rect 162162 8 164170 856
rect 164338 8 166346 856
rect 166514 8 168522 856
rect 168690 8 170698 856
rect 170866 8 172874 856
rect 173042 8 175050 856
rect 175218 8 177226 856
rect 177394 8 179402 856
rect 179570 8 181578 856
rect 181746 8 183754 856
rect 183922 8 185930 856
rect 186098 8 188106 856
rect 188274 8 190282 856
rect 190450 8 192458 856
rect 192626 8 194634 856
rect 194802 8 219998 856
rect 220166 8 222174 856
rect 222342 8 224350 856
rect 224518 8 226526 856
rect 226694 8 228702 856
rect 228870 8 230878 856
rect 231046 8 233054 856
rect 233222 8 235230 856
rect 235398 8 237406 856
rect 237574 8 239582 856
rect 239750 8 241758 856
rect 241926 8 243934 856
rect 244102 8 246110 856
rect 246278 8 248286 856
rect 248454 8 250462 856
rect 250630 8 252638 856
rect 252806 8 254814 856
rect 254982 8 256990 856
rect 257158 8 259166 856
rect 259334 8 261342 856
rect 261510 8 263518 856
rect 263686 8 265694 856
rect 265862 8 267870 856
rect 268038 8 270046 856
rect 270214 8 272222 856
rect 272390 8 274398 856
rect 274566 8 276574 856
rect 276742 8 278750 856
rect 278918 8 280926 856
rect 281094 8 283102 856
rect 283270 8 285278 856
rect 285446 8 287454 856
rect 287622 8 289630 856
rect 289798 8 291806 856
rect 291974 8 293982 856
rect 294150 8 296158 856
rect 296326 8 298334 856
rect 298502 8 300510 856
rect 300678 8 302686 856
rect 302854 8 304862 856
rect 305030 8 307038 856
rect 307206 8 309214 856
rect 309382 8 311390 856
rect 311558 8 313566 856
rect 313734 8 315742 856
rect 315910 8 317918 856
rect 318086 8 360010 856
rect 360178 8 362186 856
rect 362354 8 364362 856
rect 364530 8 366538 856
rect 366706 8 368714 856
rect 368882 8 370890 856
rect 371058 8 373066 856
rect 373234 8 375242 856
rect 375410 8 377418 856
rect 377586 8 379594 856
rect 379762 8 381770 856
rect 381938 8 383946 856
rect 384114 8 386122 856
rect 386290 8 388298 856
rect 388466 8 390474 856
rect 390642 8 392650 856
rect 392818 8 394826 856
rect 394994 8 397002 856
rect 397170 8 399178 856
rect 399346 8 401354 856
rect 401522 8 403530 856
rect 403698 8 405706 856
rect 405874 8 407882 856
rect 408050 8 410058 856
rect 410226 8 412234 856
rect 412402 8 414410 856
rect 414578 8 416586 856
rect 416754 8 418762 856
rect 418930 8 420938 856
rect 421106 8 423114 856
rect 423282 8 425290 856
rect 425458 8 427466 856
rect 427634 8 429642 856
rect 429810 8 431818 856
rect 431986 8 433994 856
rect 434162 8 436170 856
rect 436338 8 438346 856
rect 438514 8 440522 856
rect 440690 8 442698 856
rect 442866 8 444874 856
rect 445042 8 447050 856
rect 447218 8 449226 856
rect 449394 8 451402 856
rect 451570 8 453578 856
rect 453746 8 455754 856
rect 455922 8 457930 856
rect 458098 8 460106 856
rect 460274 8 462282 856
rect 462450 8 464458 856
rect 464626 8 466634 856
rect 466802 8 468810 856
rect 468978 8 470986 856
rect 471154 8 473162 856
rect 473330 8 475338 856
rect 475506 8 477514 856
rect 477682 8 479690 856
rect 479858 8 481866 856
rect 482034 8 484042 856
rect 484210 8 486218 856
rect 486386 8 488394 856
rect 488562 8 490570 856
rect 490738 8 492746 856
rect 492914 8 494922 856
rect 495090 8 497098 856
rect 497266 8 499274 856
rect 499442 8 528816 856
<< metal2 >>
rect -1076 -4 -756 11972
rect -416 656 -96 11312
rect 66908 -4 67228 11972
rect 67568 -4 67888 11972
rect 198836 -4 199156 11972
rect 199496 -4 199816 11972
rect 330764 -4 331084 11972
rect 331424 -4 331744 11972
rect 462692 -4 463012 11972
rect 463352 -4 463672 11972
rect 530016 656 530336 11312
rect 530676 -4 530996 11972
<< obsm2 >>
rect 848 2 66852 11966
rect 67284 2 67512 11966
rect 67944 2 198780 11966
rect 199212 2 199440 11966
rect 199872 2 330708 11966
rect 331140 2 331368 11966
rect 331800 2 462636 11966
rect 463068 2 463296 11966
rect 463728 2 514260 11966
<< metal3 >>
rect -1076 11652 530996 11972
rect -416 10992 530336 11312
rect -1076 9340 530996 9660
rect -1076 8680 530996 9000
rect -1076 7436 530996 7756
rect -1076 6776 530996 7096
rect -1076 5532 530996 5852
rect -1076 4872 530996 5192
rect -1076 3628 530996 3948
rect -1076 2968 530996 3288
rect -416 656 530336 976
rect -1076 -4 530996 316
<< obsm3 >>
rect 28349 11392 394023 11525
rect 28349 9740 394023 10912
rect 28349 9080 394023 9260
rect 28349 7836 394023 8600
rect 28349 7176 394023 7356
rect 28349 5932 394023 6696
rect 28349 5272 394023 5452
rect 28349 4028 394023 4792
rect 28349 3368 394023 3548
rect 28349 1056 394023 2888
rect 28349 443 394023 576
<< labels >>
rlabel metal1 s 74 0 130 800 6 ch_in[0]
port 1 nsew signal input
rlabel metal1 s 108874 0 108930 800 6 ch_in[100]
port 2 nsew signal input
rlabel metal1 s 109962 0 110018 800 6 ch_in[101]
port 3 nsew signal input
rlabel metal1 s 255550 11200 255606 12000 6 ch_in[102]
port 4 nsew signal input
rlabel metal1 s 112138 0 112194 800 6 ch_in[103]
port 5 nsew signal input
rlabel metal1 s 113226 0 113282 800 6 ch_in[104]
port 6 nsew signal input
rlabel metal1 s 257182 11200 257238 12000 6 ch_in[105]
port 7 nsew signal input
rlabel metal1 s 120026 0 120082 800 6 ch_in[106]
port 8 nsew signal input
rlabel metal1 s 360610 11200 360666 12000 6 ch_in[107]
port 9 nsew signal input
rlabel metal1 s 124378 0 124434 800 6 ch_in[108]
port 10 nsew signal input
rlabel metal1 s 361698 11200 361754 12000 6 ch_in[109]
port 11 nsew signal input
rlabel metal1 s 10954 0 11010 800 6 ch_in[10]
port 12 nsew signal input
rlabel metal1 s 128730 0 128786 800 6 ch_in[110]
port 13 nsew signal input
rlabel metal1 s 362786 11200 362842 12000 6 ch_in[111]
port 14 nsew signal input
rlabel metal1 s 133082 0 133138 800 6 ch_in[112]
port 15 nsew signal input
rlabel metal1 s 363874 11200 363930 12000 6 ch_in[113]
port 16 nsew signal input
rlabel metal1 s 137434 0 137490 800 6 ch_in[114]
port 17 nsew signal input
rlabel metal1 s 364962 11200 365018 12000 6 ch_in[115]
port 18 nsew signal input
rlabel metal1 s 141786 0 141842 800 6 ch_in[116]
port 19 nsew signal input
rlabel metal1 s 366050 11200 366106 12000 6 ch_in[117]
port 20 nsew signal input
rlabel metal1 s 146138 0 146194 800 6 ch_in[118]
port 21 nsew signal input
rlabel metal1 s 367138 11200 367194 12000 6 ch_in[119]
port 22 nsew signal input
rlabel metal1 s 12042 0 12098 800 6 ch_in[11]
port 23 nsew signal input
rlabel metal1 s 150490 0 150546 800 6 ch_in[120]
port 24 nsew signal input
rlabel metal1 s 368226 11200 368282 12000 6 ch_in[121]
port 25 nsew signal input
rlabel metal1 s 154842 0 154898 800 6 ch_in[122]
port 26 nsew signal input
rlabel metal1 s 369314 11200 369370 12000 6 ch_in[123]
port 27 nsew signal input
rlabel metal1 s 159194 0 159250 800 6 ch_in[124]
port 28 nsew signal input
rlabel metal1 s 370402 11200 370458 12000 6 ch_in[125]
port 29 nsew signal input
rlabel metal1 s 162050 0 162106 800 6 ch_in[126]
port 30 nsew signal input
rlabel metal1 s 371490 11200 371546 12000 6 ch_in[127]
port 31 nsew signal input
rlabel metal1 s 166402 0 166458 800 6 ch_in[128]
port 32 nsew signal input
rlabel metal1 s 372578 11200 372634 12000 6 ch_in[129]
port 33 nsew signal input
rlabel metal1 s 206590 11200 206646 12000 6 ch_in[12]
port 34 nsew signal input
rlabel metal1 s 170754 0 170810 800 6 ch_in[130]
port 35 nsew signal input
rlabel metal1 s 373666 11200 373722 12000 6 ch_in[131]
port 36 nsew signal input
rlabel metal1 s 175106 0 175162 800 6 ch_in[132]
port 37 nsew signal input
rlabel metal1 s 374754 11200 374810 12000 6 ch_in[133]
port 38 nsew signal input
rlabel metal1 s 179458 0 179514 800 6 ch_in[134]
port 39 nsew signal input
rlabel metal1 s 375842 11200 375898 12000 6 ch_in[135]
port 40 nsew signal input
rlabel metal1 s 183810 0 183866 800 6 ch_in[136]
port 41 nsew signal input
rlabel metal1 s 376930 11200 376986 12000 6 ch_in[137]
port 42 nsew signal input
rlabel metal1 s 188162 0 188218 800 6 ch_in[138]
port 43 nsew signal input
rlabel metal1 s 378018 11200 378074 12000 6 ch_in[139]
port 44 nsew signal input
rlabel metal1 s 14218 0 14274 800 6 ch_in[13]
port 45 nsew signal input
rlabel metal1 s 192514 0 192570 800 6 ch_in[140]
port 46 nsew signal input
rlabel metal1 s 379106 11200 379162 12000 6 ch_in[141]
port 47 nsew signal input
rlabel metal1 s 379650 11200 379706 12000 6 ch_in[142]
port 48 nsew signal input
rlabel metal1 s 380194 11200 380250 12000 6 ch_in[143]
port 49 nsew signal input
rlabel metal1 s 380738 11200 380794 12000 6 ch_in[144]
port 50 nsew signal input
rlabel metal1 s 381282 11200 381338 12000 6 ch_in[145]
port 51 nsew signal input
rlabel metal1 s 381826 11200 381882 12000 6 ch_in[146]
port 52 nsew signal input
rlabel metal1 s 382370 11200 382426 12000 6 ch_in[147]
port 53 nsew signal input
rlabel metal1 s 382914 11200 382970 12000 6 ch_in[148]
port 54 nsew signal input
rlabel metal1 s 383458 11200 383514 12000 6 ch_in[149]
port 55 nsew signal input
rlabel metal1 s 15306 0 15362 800 6 ch_in[14]
port 56 nsew signal input
rlabel metal1 s 384002 11200 384058 12000 6 ch_in[150]
port 57 nsew signal input
rlabel metal1 s 384546 11172 384602 12000 6 ch_in[151]
port 58 nsew signal input
rlabel metal1 s 385090 11200 385146 12000 6 ch_in[152]
port 59 nsew signal input
rlabel metal1 s 385634 11200 385690 12000 6 ch_in[153]
port 60 nsew signal input
rlabel metal1 s 386178 11200 386234 12000 6 ch_in[154]
port 61 nsew signal input
rlabel metal1 s 386722 11200 386778 12000 6 ch_in[155]
port 62 nsew signal input
rlabel metal1 s 387266 11200 387322 12000 6 ch_in[156]
port 63 nsew signal input
rlabel metal1 s 387810 11200 387866 12000 6 ch_in[157]
port 64 nsew signal input
rlabel metal1 s 388354 11200 388410 12000 6 ch_in[158]
port 65 nsew signal input
rlabel metal1 s 388898 11200 388954 12000 6 ch_in[159]
port 66 nsew signal input
rlabel metal1 s 16394 0 16450 800 6 ch_in[15]
port 67 nsew signal input
rlabel metal1 s 389442 11200 389498 12000 6 ch_in[160]
port 68 nsew signal input
rlabel metal1 s 389986 11200 390042 12000 6 ch_in[161]
port 69 nsew signal input
rlabel metal1 s 390530 11200 390586 12000 6 ch_in[162]
port 70 nsew signal input
rlabel metal1 s 391074 11200 391130 12000 6 ch_in[163]
port 71 nsew signal input
rlabel metal1 s 391618 11200 391674 12000 6 ch_in[164]
port 72 nsew signal input
rlabel metal1 s 392162 11200 392218 12000 6 ch_in[165]
port 73 nsew signal input
rlabel metal1 s 392706 11200 392762 12000 6 ch_in[166]
port 74 nsew signal input
rlabel metal1 s 393250 11200 393306 12000 6 ch_in[167]
port 75 nsew signal input
rlabel metal1 s 393794 11200 393850 12000 6 ch_in[168]
port 76 nsew signal input
rlabel metal1 s 394338 11200 394394 12000 6 ch_in[169]
port 77 nsew signal input
rlabel metal1 s 208766 11200 208822 12000 6 ch_in[16]
port 78 nsew signal input
rlabel metal1 s 394882 11200 394938 12000 6 ch_in[170]
port 79 nsew signal input
rlabel metal1 s 395426 11200 395482 12000 6 ch_in[171]
port 80 nsew signal input
rlabel metal1 s 395970 11200 396026 12000 6 ch_in[172]
port 81 nsew signal input
rlabel metal1 s 396514 11200 396570 12000 6 ch_in[173]
port 82 nsew signal input
rlabel metal1 s 397058 11172 397114 12000 6 ch_in[174]
port 83 nsew signal input
rlabel metal1 s 397602 11200 397658 12000 6 ch_in[175]
port 84 nsew signal input
rlabel metal1 s 398146 11200 398202 12000 6 ch_in[176]
port 85 nsew signal input
rlabel metal1 s 398690 11200 398746 12000 6 ch_in[177]
port 86 nsew signal input
rlabel metal1 s 399234 11200 399290 12000 6 ch_in[178]
port 87 nsew signal input
rlabel metal1 s 399778 11200 399834 12000 6 ch_in[179]
port 88 nsew signal input
rlabel metal1 s 18570 0 18626 800 6 ch_in[17]
port 89 nsew signal input
rlabel metal1 s 400322 11200 400378 12000 6 ch_in[180]
port 90 nsew signal input
rlabel metal1 s 400866 11200 400922 12000 6 ch_in[181]
port 91 nsew signal input
rlabel metal1 s 401410 11200 401466 12000 6 ch_in[182]
port 92 nsew signal input
rlabel metal1 s 401954 11200 402010 12000 6 ch_in[183]
port 93 nsew signal input
rlabel metal1 s 402498 11200 402554 12000 6 ch_in[184]
port 94 nsew signal input
rlabel metal1 s 403042 11200 403098 12000 6 ch_in[185]
port 95 nsew signal input
rlabel metal1 s 403586 11200 403642 12000 6 ch_in[186]
port 96 nsew signal input
rlabel metal1 s 404130 11200 404186 12000 6 ch_in[187]
port 97 nsew signal input
rlabel metal1 s 440034 11200 440090 12000 6 ch_in[188]
port 98 nsew signal input
rlabel metal1 s 440306 11200 440362 12000 6 ch_in[189]
port 99 nsew signal input
rlabel metal1 s 19658 0 19714 800 6 ch_in[18]
port 100 nsew signal input
rlabel metal1 s 440578 11200 440634 12000 6 ch_in[190]
port 101 nsew signal input
rlabel metal1 s 440850 11200 440906 12000 6 ch_in[191]
port 102 nsew signal input
rlabel metal1 s 441122 11200 441178 12000 6 ch_in[192]
port 103 nsew signal input
rlabel metal1 s 441394 11200 441450 12000 6 ch_in[193]
port 104 nsew signal input
rlabel metal1 s 441666 11200 441722 12000 6 ch_in[194]
port 105 nsew signal input
rlabel metal1 s 441938 11200 441994 12000 6 ch_in[195]
port 106 nsew signal input
rlabel metal1 s 442210 11200 442266 12000 6 ch_in[196]
port 107 nsew signal input
rlabel metal1 s 442482 11200 442538 12000 6 ch_in[197]
port 108 nsew signal input
rlabel metal1 s 442754 11172 442810 12000 6 ch_in[198]
port 109 nsew signal input
rlabel metal1 s 443026 11200 443082 12000 6 ch_in[199]
port 110 nsew signal input
rlabel metal1 s 20746 0 20802 800 6 ch_in[19]
port 111 nsew signal input
rlabel metal1 s 1162 0 1218 800 6 ch_in[1]
port 112 nsew signal input
rlabel metal1 s 443298 11200 443354 12000 6 ch_in[200]
port 113 nsew signal input
rlabel metal1 s 443570 11200 443626 12000 6 ch_in[201]
port 114 nsew signal input
rlabel metal1 s 443842 11200 443898 12000 6 ch_in[202]
port 115 nsew signal input
rlabel metal1 s 444114 11200 444170 12000 6 ch_in[203]
port 116 nsew signal input
rlabel metal1 s 444386 11200 444442 12000 6 ch_in[204]
port 117 nsew signal input
rlabel metal1 s 444658 11200 444714 12000 6 ch_in[205]
port 118 nsew signal input
rlabel metal1 s 444930 11200 444986 12000 6 ch_in[206]
port 119 nsew signal input
rlabel metal1 s 445202 11200 445258 12000 6 ch_in[207]
port 120 nsew signal input
rlabel metal1 s 445474 11200 445530 12000 6 ch_in[208]
port 121 nsew signal input
rlabel metal1 s 445746 11200 445802 12000 6 ch_in[209]
port 122 nsew signal input
rlabel metal1 s 210942 11200 210998 12000 6 ch_in[20]
port 123 nsew signal input
rlabel metal1 s 446018 11200 446074 12000 6 ch_in[210]
port 124 nsew signal input
rlabel metal1 s 446290 11200 446346 12000 6 ch_in[211]
port 125 nsew signal input
rlabel metal1 s 446562 11200 446618 12000 6 ch_in[212]
port 126 nsew signal input
rlabel metal1 s 446834 11200 446890 12000 6 ch_in[213]
port 127 nsew signal input
rlabel metal1 s 447106 11172 447162 12000 6 ch_in[214]
port 128 nsew signal input
rlabel metal1 s 447378 11200 447434 12000 6 ch_in[215]
port 129 nsew signal input
rlabel metal1 s 447650 11200 447706 12000 6 ch_in[216]
port 130 nsew signal input
rlabel metal1 s 447922 11200 447978 12000 6 ch_in[217]
port 131 nsew signal input
rlabel metal1 s 448194 11200 448250 12000 6 ch_in[218]
port 132 nsew signal input
rlabel metal1 s 448466 11200 448522 12000 6 ch_in[219]
port 133 nsew signal input
rlabel metal1 s 22922 0 22978 800 6 ch_in[21]
port 134 nsew signal input
rlabel metal1 s 480018 11200 480074 12000 6 ch_in[220]
port 135 nsew signal input
rlabel metal1 s 480290 11172 480346 12000 6 ch_in[221]
port 136 nsew signal input
rlabel metal1 s 480562 11200 480618 12000 6 ch_in[222]
port 137 nsew signal input
rlabel metal1 s 480834 11200 480890 12000 6 ch_in[223]
port 138 nsew signal input
rlabel metal1 s 481106 11200 481162 12000 6 ch_in[224]
port 139 nsew signal input
rlabel metal1 s 481378 11200 481434 12000 6 ch_in[225]
port 140 nsew signal input
rlabel metal1 s 481650 11200 481706 12000 6 ch_in[226]
port 141 nsew signal input
rlabel metal1 s 481922 11200 481978 12000 6 ch_in[227]
port 142 nsew signal input
rlabel metal1 s 482194 11200 482250 12000 6 ch_in[228]
port 143 nsew signal input
rlabel metal1 s 482466 11200 482522 12000 6 ch_in[229]
port 144 nsew signal input
rlabel metal1 s 24010 0 24066 800 6 ch_in[22]
port 145 nsew signal input
rlabel metal1 s 482738 11200 482794 12000 6 ch_in[230]
port 146 nsew signal input
rlabel metal1 s 483010 11172 483066 12000 6 ch_in[231]
port 147 nsew signal input
rlabel metal1 s 483282 11200 483338 12000 6 ch_in[232]
port 148 nsew signal input
rlabel metal1 s 483554 11200 483610 12000 6 ch_in[233]
port 149 nsew signal input
rlabel metal1 s 483826 11200 483882 12000 6 ch_in[234]
port 150 nsew signal input
rlabel metal1 s 484098 11200 484154 12000 6 ch_in[235]
port 151 nsew signal input
rlabel metal1 s 484370 11200 484426 12000 6 ch_in[236]
port 152 nsew signal input
rlabel metal1 s 484642 11200 484698 12000 6 ch_in[237]
port 153 nsew signal input
rlabel metal1 s 484914 11200 484970 12000 6 ch_in[238]
port 154 nsew signal input
rlabel metal1 s 485186 11200 485242 12000 6 ch_in[239]
port 155 nsew signal input
rlabel metal1 s 25098 0 25154 800 6 ch_in[23]
port 156 nsew signal input
rlabel metal1 s 485458 11200 485514 12000 6 ch_in[240]
port 157 nsew signal input
rlabel metal1 s 485730 11200 485786 12000 6 ch_in[241]
port 158 nsew signal input
rlabel metal1 s 486002 11200 486058 12000 6 ch_in[242]
port 159 nsew signal input
rlabel metal1 s 486274 11200 486330 12000 6 ch_in[243]
port 160 nsew signal input
rlabel metal1 s 486546 11200 486602 12000 6 ch_in[244]
port 161 nsew signal input
rlabel metal1 s 486818 11200 486874 12000 6 ch_in[245]
port 162 nsew signal input
rlabel metal1 s 487090 11200 487146 12000 6 ch_in[246]
port 163 nsew signal input
rlabel metal1 s 487362 11200 487418 12000 6 ch_in[247]
port 164 nsew signal input
rlabel metal1 s 487634 11200 487690 12000 6 ch_in[248]
port 165 nsew signal input
rlabel metal1 s 487906 11200 487962 12000 6 ch_in[249]
port 166 nsew signal input
rlabel metal1 s 213118 11200 213174 12000 6 ch_in[24]
port 167 nsew signal input
rlabel metal1 s 488178 11200 488234 12000 6 ch_in[250]
port 168 nsew signal input
rlabel metal1 s 488450 11200 488506 12000 6 ch_in[251]
port 169 nsew signal input
rlabel metal1 s 499330 0 499386 800 6 ch_in[252]
port 170 nsew signal input
rlabel metal1 s 27274 0 27330 800 6 ch_in[25]
port 171 nsew signal input
rlabel metal1 s 28362 0 28418 800 6 ch_in[26]
port 172 nsew signal input
rlabel metal1 s 214750 11200 214806 12000 6 ch_in[27]
port 173 nsew signal input
rlabel metal1 s 30538 0 30594 800 6 ch_in[28]
port 174 nsew signal input
rlabel metal1 s 31626 0 31682 800 6 ch_in[29]
port 175 nsew signal input
rlabel metal1 s 201150 11200 201206 12000 6 ch_in[2]
port 176 nsew signal input
rlabel metal1 s 216382 11200 216438 12000 6 ch_in[30]
port 177 nsew signal input
rlabel metal1 s 33802 0 33858 800 6 ch_in[31]
port 178 nsew signal input
rlabel metal1 s 34890 0 34946 800 6 ch_in[32]
port 179 nsew signal input
rlabel metal1 s 218014 11200 218070 12000 6 ch_in[33]
port 180 nsew signal input
rlabel metal1 s 37066 0 37122 800 6 ch_in[34]
port 181 nsew signal input
rlabel metal1 s 38154 0 38210 800 6 ch_in[35]
port 182 nsew signal input
rlabel metal1 s 219646 11200 219702 12000 6 ch_in[36]
port 183 nsew signal input
rlabel metal1 s 40330 0 40386 800 6 ch_in[37]
port 184 nsew signal input
rlabel metal1 s 41418 0 41474 800 6 ch_in[38]
port 185 nsew signal input
rlabel metal1 s 221278 11200 221334 12000 6 ch_in[39]
port 186 nsew signal input
rlabel metal1 s 3338 0 3394 800 6 ch_in[3]
port 187 nsew signal input
rlabel metal1 s 43594 0 43650 800 6 ch_in[40]
port 188 nsew signal input
rlabel metal1 s 44682 0 44738 800 6 ch_in[41]
port 189 nsew signal input
rlabel metal1 s 222910 11200 222966 12000 6 ch_in[42]
port 190 nsew signal input
rlabel metal1 s 46858 0 46914 800 6 ch_in[43]
port 191 nsew signal input
rlabel metal1 s 47946 0 48002 800 6 ch_in[44]
port 192 nsew signal input
rlabel metal1 s 224542 11200 224598 12000 6 ch_in[45]
port 193 nsew signal input
rlabel metal1 s 50122 0 50178 800 6 ch_in[46]
port 194 nsew signal input
rlabel metal1 s 51210 0 51266 800 6 ch_in[47]
port 195 nsew signal input
rlabel metal1 s 226174 11200 226230 12000 6 ch_in[48]
port 196 nsew signal input
rlabel metal1 s 53386 0 53442 800 6 ch_in[49]
port 197 nsew signal input
rlabel metal1 s 4426 0 4482 800 6 ch_in[4]
port 198 nsew signal input
rlabel metal1 s 54474 0 54530 800 6 ch_in[50]
port 199 nsew signal input
rlabel metal1 s 227806 11200 227862 12000 6 ch_in[51]
port 200 nsew signal input
rlabel metal1 s 56650 0 56706 800 6 ch_in[52]
port 201 nsew signal input
rlabel metal1 s 57738 0 57794 800 6 ch_in[53]
port 202 nsew signal input
rlabel metal1 s 229438 11200 229494 12000 6 ch_in[54]
port 203 nsew signal input
rlabel metal1 s 59914 0 59970 800 6 ch_in[55]
port 204 nsew signal input
rlabel metal1 s 61002 0 61058 800 6 ch_in[56]
port 205 nsew signal input
rlabel metal1 s 231070 11200 231126 12000 6 ch_in[57]
port 206 nsew signal input
rlabel metal1 s 63178 0 63234 800 6 ch_in[58]
port 207 nsew signal input
rlabel metal1 s 64266 0 64322 800 6 ch_in[59]
port 208 nsew signal input
rlabel metal1 s 5514 0 5570 800 6 ch_in[5]
port 209 nsew signal input
rlabel metal1 s 232702 11200 232758 12000 6 ch_in[60]
port 210 nsew signal input
rlabel metal1 s 66442 0 66498 800 6 ch_in[61]
port 211 nsew signal input
rlabel metal1 s 67530 0 67586 800 6 ch_in[62]
port 212 nsew signal input
rlabel metal1 s 234334 11200 234390 12000 6 ch_in[63]
port 213 nsew signal input
rlabel metal1 s 69706 0 69762 800 6 ch_in[64]
port 214 nsew signal input
rlabel metal1 s 70794 0 70850 800 6 ch_in[65]
port 215 nsew signal input
rlabel metal1 s 235966 11200 236022 12000 6 ch_in[66]
port 216 nsew signal input
rlabel metal1 s 72970 0 73026 800 6 ch_in[67]
port 217 nsew signal input
rlabel metal1 s 74058 0 74114 800 6 ch_in[68]
port 218 nsew signal input
rlabel metal1 s 237598 11200 237654 12000 6 ch_in[69]
port 219 nsew signal input
rlabel metal1 s 6602 0 6658 800 6 ch_in[6]
port 220 nsew signal input
rlabel metal1 s 76234 0 76290 800 6 ch_in[70]
port 221 nsew signal input
rlabel metal1 s 77322 0 77378 800 6 ch_in[71]
port 222 nsew signal input
rlabel metal1 s 239230 11200 239286 12000 6 ch_in[72]
port 223 nsew signal input
rlabel metal1 s 79498 0 79554 800 6 ch_in[73]
port 224 nsew signal input
rlabel metal1 s 80586 0 80642 800 6 ch_in[74]
port 225 nsew signal input
rlabel metal1 s 240862 11200 240918 12000 6 ch_in[75]
port 226 nsew signal input
rlabel metal1 s 82762 0 82818 800 6 ch_in[76]
port 227 nsew signal input
rlabel metal1 s 83850 0 83906 800 6 ch_in[77]
port 228 nsew signal input
rlabel metal1 s 242494 11200 242550 12000 6 ch_in[78]
port 229 nsew signal input
rlabel metal1 s 86026 0 86082 800 6 ch_in[79]
port 230 nsew signal input
rlabel metal1 s 7690 0 7746 800 6 ch_in[7]
port 231 nsew signal input
rlabel metal1 s 87114 0 87170 800 6 ch_in[80]
port 232 nsew signal input
rlabel metal1 s 244126 11172 244182 12000 6 ch_in[81]
port 233 nsew signal input
rlabel metal1 s 89290 0 89346 800 6 ch_in[82]
port 234 nsew signal input
rlabel metal1 s 90378 0 90434 800 6 ch_in[83]
port 235 nsew signal input
rlabel metal1 s 245758 11200 245814 12000 6 ch_in[84]
port 236 nsew signal input
rlabel metal1 s 92554 0 92610 800 6 ch_in[85]
port 237 nsew signal input
rlabel metal1 s 93642 0 93698 800 6 ch_in[86]
port 238 nsew signal input
rlabel metal1 s 247390 11200 247446 12000 6 ch_in[87]
port 239 nsew signal input
rlabel metal1 s 95818 0 95874 800 6 ch_in[88]
port 240 nsew signal input
rlabel metal1 s 96906 0 96962 800 6 ch_in[89]
port 241 nsew signal input
rlabel metal1 s 204414 11200 204470 12000 6 ch_in[8]
port 242 nsew signal input
rlabel metal1 s 249022 11200 249078 12000 6 ch_in[90]
port 243 nsew signal input
rlabel metal1 s 99082 0 99138 800 6 ch_in[91]
port 244 nsew signal input
rlabel metal1 s 100170 0 100226 800 6 ch_in[92]
port 245 nsew signal input
rlabel metal1 s 250654 11200 250710 12000 6 ch_in[93]
port 246 nsew signal input
rlabel metal1 s 102346 0 102402 800 6 ch_in[94]
port 247 nsew signal input
rlabel metal1 s 103434 0 103490 800 6 ch_in[95]
port 248 nsew signal input
rlabel metal1 s 252286 11200 252342 12000 6 ch_in[96]
port 249 nsew signal input
rlabel metal1 s 105610 0 105666 800 6 ch_in[97]
port 250 nsew signal input
rlabel metal1 s 106698 0 106754 800 6 ch_in[98]
port 251 nsew signal input
rlabel metal1 s 253918 11200 253974 12000 6 ch_in[99]
port 252 nsew signal input
rlabel metal1 s 9866 0 9922 800 6 ch_in[9]
port 253 nsew signal input
rlabel metal1 s 200062 11200 200118 12000 6 ch_out[0]
port 254 nsew signal output
rlabel metal1 s 254462 11200 254518 12000 6 ch_out[100]
port 255 nsew signal output
rlabel metal1 s 255006 11200 255062 12000 6 ch_out[101]
port 256 nsew signal output
rlabel metal1 s 111050 0 111106 800 6 ch_out[102]
port 257 nsew signal output
rlabel metal1 s 256094 11200 256150 12000 6 ch_out[103]
port 258 nsew signal output
rlabel metal1 s 256638 11200 256694 12000 6 ch_out[104]
port 259 nsew signal output
rlabel metal1 s 114314 0 114370 800 6 ch_out[105]
port 260 nsew signal output
rlabel metal1 s 360066 11200 360122 12000 6 ch_out[106]
port 261 nsew signal output
rlabel metal1 s 122202 0 122258 800 6 ch_out[107]
port 262 nsew signal output
rlabel metal1 s 361154 11200 361210 12000 6 ch_out[108]
port 263 nsew signal output
rlabel metal1 s 126554 0 126610 800 6 ch_out[109]
port 264 nsew signal output
rlabel metal1 s 205502 11200 205558 12000 6 ch_out[10]
port 265 nsew signal output
rlabel metal1 s 362242 11200 362298 12000 6 ch_out[110]
port 266 nsew signal output
rlabel metal1 s 130906 0 130962 800 6 ch_out[111]
port 267 nsew signal output
rlabel metal1 s 363330 11200 363386 12000 6 ch_out[112]
port 268 nsew signal output
rlabel metal1 s 135258 0 135314 800 6 ch_out[113]
port 269 nsew signal output
rlabel metal1 s 364418 11200 364474 12000 6 ch_out[114]
port 270 nsew signal output
rlabel metal1 s 139610 0 139666 800 6 ch_out[115]
port 271 nsew signal output
rlabel metal1 s 365506 11200 365562 12000 6 ch_out[116]
port 272 nsew signal output
rlabel metal1 s 143962 0 144018 800 6 ch_out[117]
port 273 nsew signal output
rlabel metal1 s 366594 11200 366650 12000 6 ch_out[118]
port 274 nsew signal output
rlabel metal1 s 148314 0 148370 800 6 ch_out[119]
port 275 nsew signal output
rlabel metal1 s 206046 11200 206102 12000 6 ch_out[11]
port 276 nsew signal output
rlabel metal1 s 367682 11200 367738 12000 6 ch_out[120]
port 277 nsew signal output
rlabel metal1 s 152666 0 152722 800 6 ch_out[121]
port 278 nsew signal output
rlabel metal1 s 368770 11200 368826 12000 6 ch_out[122]
port 279 nsew signal output
rlabel metal1 s 157018 0 157074 800 6 ch_out[123]
port 280 nsew signal output
rlabel metal1 s 369858 11200 369914 12000 6 ch_out[124]
port 281 nsew signal output
rlabel metal1 s 161370 0 161426 800 6 ch_out[125]
port 282 nsew signal output
rlabel metal1 s 370946 11200 371002 12000 6 ch_out[126]
port 283 nsew signal output
rlabel metal1 s 164226 0 164282 800 6 ch_out[127]
port 284 nsew signal output
rlabel metal1 s 372034 11200 372090 12000 6 ch_out[128]
port 285 nsew signal output
rlabel metal1 s 168578 0 168634 800 6 ch_out[129]
port 286 nsew signal output
rlabel metal1 s 13130 0 13186 800 6 ch_out[12]
port 287 nsew signal output
rlabel metal1 s 373122 11200 373178 12000 6 ch_out[130]
port 288 nsew signal output
rlabel metal1 s 172930 0 172986 800 6 ch_out[131]
port 289 nsew signal output
rlabel metal1 s 374210 11200 374266 12000 6 ch_out[132]
port 290 nsew signal output
rlabel metal1 s 177282 0 177338 800 6 ch_out[133]
port 291 nsew signal output
rlabel metal1 s 375298 11200 375354 12000 6 ch_out[134]
port 292 nsew signal output
rlabel metal1 s 181634 0 181690 800 6 ch_out[135]
port 293 nsew signal output
rlabel metal1 s 376386 11200 376442 12000 6 ch_out[136]
port 294 nsew signal output
rlabel metal1 s 185986 0 186042 800 6 ch_out[137]
port 295 nsew signal output
rlabel metal1 s 377474 11200 377530 12000 6 ch_out[138]
port 296 nsew signal output
rlabel metal1 s 190338 0 190394 800 6 ch_out[139]
port 297 nsew signal output
rlabel metal1 s 207134 11200 207190 12000 6 ch_out[13]
port 298 nsew signal output
rlabel metal1 s 378562 11200 378618 12000 6 ch_out[140]
port 299 nsew signal output
rlabel metal1 s 194690 0 194746 800 6 ch_out[141]
port 300 nsew signal output
rlabel metal1 s 220054 0 220110 800 6 ch_out[142]
port 301 nsew signal output
rlabel metal1 s 222230 0 222286 800 6 ch_out[143]
port 302 nsew signal output
rlabel metal1 s 224406 0 224462 800 6 ch_out[144]
port 303 nsew signal output
rlabel metal1 s 226582 0 226638 800 6 ch_out[145]
port 304 nsew signal output
rlabel metal1 s 228758 0 228814 800 6 ch_out[146]
port 305 nsew signal output
rlabel metal1 s 230934 0 230990 800 6 ch_out[147]
port 306 nsew signal output
rlabel metal1 s 233110 0 233166 800 6 ch_out[148]
port 307 nsew signal output
rlabel metal1 s 235286 0 235342 800 6 ch_out[149]
port 308 nsew signal output
rlabel metal1 s 207678 11200 207734 12000 6 ch_out[14]
port 309 nsew signal output
rlabel metal1 s 237462 0 237518 800 6 ch_out[150]
port 310 nsew signal output
rlabel metal1 s 239638 0 239694 800 6 ch_out[151]
port 311 nsew signal output
rlabel metal1 s 241814 0 241870 800 6 ch_out[152]
port 312 nsew signal output
rlabel metal1 s 243990 0 244046 800 6 ch_out[153]
port 313 nsew signal output
rlabel metal1 s 246166 0 246222 800 6 ch_out[154]
port 314 nsew signal output
rlabel metal1 s 248342 0 248398 800 6 ch_out[155]
port 315 nsew signal output
rlabel metal1 s 250518 0 250574 800 6 ch_out[156]
port 316 nsew signal output
rlabel metal1 s 252694 0 252750 800 6 ch_out[157]
port 317 nsew signal output
rlabel metal1 s 254870 0 254926 800 6 ch_out[158]
port 318 nsew signal output
rlabel metal1 s 257046 0 257102 800 6 ch_out[159]
port 319 nsew signal output
rlabel metal1 s 208222 11200 208278 12000 6 ch_out[15]
port 320 nsew signal output
rlabel metal1 s 259222 0 259278 800 6 ch_out[160]
port 321 nsew signal output
rlabel metal1 s 261398 0 261454 800 6 ch_out[161]
port 322 nsew signal output
rlabel metal1 s 263574 0 263630 800 6 ch_out[162]
port 323 nsew signal output
rlabel metal1 s 265750 0 265806 800 6 ch_out[163]
port 324 nsew signal output
rlabel metal1 s 267926 0 267982 800 6 ch_out[164]
port 325 nsew signal output
rlabel metal1 s 270102 0 270158 800 6 ch_out[165]
port 326 nsew signal output
rlabel metal1 s 272278 0 272334 800 6 ch_out[166]
port 327 nsew signal output
rlabel metal1 s 274454 0 274510 800 6 ch_out[167]
port 328 nsew signal output
rlabel metal1 s 276630 0 276686 800 6 ch_out[168]
port 329 nsew signal output
rlabel metal1 s 278806 0 278862 800 6 ch_out[169]
port 330 nsew signal output
rlabel metal1 s 17482 0 17538 800 6 ch_out[16]
port 331 nsew signal output
rlabel metal1 s 280982 0 281038 800 6 ch_out[170]
port 332 nsew signal output
rlabel metal1 s 283158 0 283214 800 6 ch_out[171]
port 333 nsew signal output
rlabel metal1 s 285334 0 285390 800 6 ch_out[172]
port 334 nsew signal output
rlabel metal1 s 287510 0 287566 800 6 ch_out[173]
port 335 nsew signal output
rlabel metal1 s 289686 0 289742 800 6 ch_out[174]
port 336 nsew signal output
rlabel metal1 s 291862 0 291918 800 6 ch_out[175]
port 337 nsew signal output
rlabel metal1 s 294038 0 294094 800 6 ch_out[176]
port 338 nsew signal output
rlabel metal1 s 296214 0 296270 800 6 ch_out[177]
port 339 nsew signal output
rlabel metal1 s 298390 0 298446 800 6 ch_out[178]
port 340 nsew signal output
rlabel metal1 s 300566 0 300622 800 6 ch_out[179]
port 341 nsew signal output
rlabel metal1 s 209310 11200 209366 12000 6 ch_out[17]
port 342 nsew signal output
rlabel metal1 s 302742 0 302798 800 6 ch_out[180]
port 343 nsew signal output
rlabel metal1 s 304918 0 304974 800 6 ch_out[181]
port 344 nsew signal output
rlabel metal1 s 307094 0 307150 800 6 ch_out[182]
port 345 nsew signal output
rlabel metal1 s 309270 0 309326 800 6 ch_out[183]
port 346 nsew signal output
rlabel metal1 s 311446 0 311502 800 6 ch_out[184]
port 347 nsew signal output
rlabel metal1 s 313622 0 313678 800 6 ch_out[185]
port 348 nsew signal output
rlabel metal1 s 315798 0 315854 800 6 ch_out[186]
port 349 nsew signal output
rlabel metal1 s 317974 0 318030 800 6 ch_out[187]
port 350 nsew signal output
rlabel metal1 s 360066 0 360122 800 6 ch_out[188]
port 351 nsew signal output
rlabel metal1 s 362242 0 362298 800 6 ch_out[189]
port 352 nsew signal output
rlabel metal1 s 209854 11200 209910 12000 6 ch_out[18]
port 353 nsew signal output
rlabel metal1 s 364418 0 364474 800 6 ch_out[190]
port 354 nsew signal output
rlabel metal1 s 366594 0 366650 800 6 ch_out[191]
port 355 nsew signal output
rlabel metal1 s 368770 0 368826 800 6 ch_out[192]
port 356 nsew signal output
rlabel metal1 s 370946 0 371002 800 6 ch_out[193]
port 357 nsew signal output
rlabel metal1 s 373122 0 373178 800 6 ch_out[194]
port 358 nsew signal output
rlabel metal1 s 375298 0 375354 800 6 ch_out[195]
port 359 nsew signal output
rlabel metal1 s 377474 0 377530 800 6 ch_out[196]
port 360 nsew signal output
rlabel metal1 s 379650 0 379706 800 6 ch_out[197]
port 361 nsew signal output
rlabel metal1 s 381826 0 381882 800 6 ch_out[198]
port 362 nsew signal output
rlabel metal1 s 384002 0 384058 800 6 ch_out[199]
port 363 nsew signal output
rlabel metal1 s 210398 11200 210454 12000 6 ch_out[19]
port 364 nsew signal output
rlabel metal1 s 200606 11200 200662 12000 6 ch_out[1]
port 365 nsew signal output
rlabel metal1 s 386178 0 386234 800 6 ch_out[200]
port 366 nsew signal output
rlabel metal1 s 388354 0 388410 800 6 ch_out[201]
port 367 nsew signal output
rlabel metal1 s 390530 0 390586 800 6 ch_out[202]
port 368 nsew signal output
rlabel metal1 s 392706 0 392762 800 6 ch_out[203]
port 369 nsew signal output
rlabel metal1 s 394882 0 394938 800 6 ch_out[204]
port 370 nsew signal output
rlabel metal1 s 397058 0 397114 800 6 ch_out[205]
port 371 nsew signal output
rlabel metal1 s 399234 0 399290 800 6 ch_out[206]
port 372 nsew signal output
rlabel metal1 s 401410 0 401466 800 6 ch_out[207]
port 373 nsew signal output
rlabel metal1 s 403586 0 403642 800 6 ch_out[208]
port 374 nsew signal output
rlabel metal1 s 405762 0 405818 800 6 ch_out[209]
port 375 nsew signal output
rlabel metal1 s 21834 0 21890 800 6 ch_out[20]
port 376 nsew signal output
rlabel metal1 s 407938 0 407994 800 6 ch_out[210]
port 377 nsew signal output
rlabel metal1 s 410114 0 410170 800 6 ch_out[211]
port 378 nsew signal output
rlabel metal1 s 412290 0 412346 800 6 ch_out[212]
port 379 nsew signal output
rlabel metal1 s 414466 0 414522 800 6 ch_out[213]
port 380 nsew signal output
rlabel metal1 s 416642 0 416698 800 6 ch_out[214]
port 381 nsew signal output
rlabel metal1 s 418818 0 418874 800 6 ch_out[215]
port 382 nsew signal output
rlabel metal1 s 420994 0 421050 800 6 ch_out[216]
port 383 nsew signal output
rlabel metal1 s 423170 0 423226 800 6 ch_out[217]
port 384 nsew signal output
rlabel metal1 s 425346 0 425402 800 6 ch_out[218]
port 385 nsew signal output
rlabel metal1 s 427522 0 427578 800 6 ch_out[219]
port 386 nsew signal output
rlabel metal1 s 211486 11200 211542 12000 6 ch_out[21]
port 387 nsew signal output
rlabel metal1 s 429698 0 429754 800 6 ch_out[220]
port 388 nsew signal output
rlabel metal1 s 431874 0 431930 800 6 ch_out[221]
port 389 nsew signal output
rlabel metal1 s 434050 0 434106 800 6 ch_out[222]
port 390 nsew signal output
rlabel metal1 s 436226 0 436282 800 6 ch_out[223]
port 391 nsew signal output
rlabel metal1 s 438402 0 438458 800 6 ch_out[224]
port 392 nsew signal output
rlabel metal1 s 440578 0 440634 800 6 ch_out[225]
port 393 nsew signal output
rlabel metal1 s 442754 0 442810 800 6 ch_out[226]
port 394 nsew signal output
rlabel metal1 s 444930 0 444986 800 6 ch_out[227]
port 395 nsew signal output
rlabel metal1 s 447106 0 447162 800 6 ch_out[228]
port 396 nsew signal output
rlabel metal1 s 449282 0 449338 800 6 ch_out[229]
port 397 nsew signal output
rlabel metal1 s 212030 11200 212086 12000 6 ch_out[22]
port 398 nsew signal output
rlabel metal1 s 451458 0 451514 800 6 ch_out[230]
port 399 nsew signal output
rlabel metal1 s 453634 0 453690 800 6 ch_out[231]
port 400 nsew signal output
rlabel metal1 s 455810 0 455866 800 6 ch_out[232]
port 401 nsew signal output
rlabel metal1 s 457986 0 458042 800 6 ch_out[233]
port 402 nsew signal output
rlabel metal1 s 460162 0 460218 800 6 ch_out[234]
port 403 nsew signal output
rlabel metal1 s 462338 0 462394 800 6 ch_out[235]
port 404 nsew signal output
rlabel metal1 s 464514 0 464570 800 6 ch_out[236]
port 405 nsew signal output
rlabel metal1 s 466690 0 466746 800 6 ch_out[237]
port 406 nsew signal output
rlabel metal1 s 468866 0 468922 800 6 ch_out[238]
port 407 nsew signal output
rlabel metal1 s 471042 0 471098 800 6 ch_out[239]
port 408 nsew signal output
rlabel metal1 s 212574 11200 212630 12000 6 ch_out[23]
port 409 nsew signal output
rlabel metal1 s 473218 0 473274 800 6 ch_out[240]
port 410 nsew signal output
rlabel metal1 s 475394 0 475450 800 6 ch_out[241]
port 411 nsew signal output
rlabel metal1 s 477570 0 477626 800 6 ch_out[242]
port 412 nsew signal output
rlabel metal1 s 479746 0 479802 800 6 ch_out[243]
port 413 nsew signal output
rlabel metal1 s 481922 0 481978 800 6 ch_out[244]
port 414 nsew signal output
rlabel metal1 s 484098 0 484154 800 6 ch_out[245]
port 415 nsew signal output
rlabel metal1 s 486274 0 486330 800 6 ch_out[246]
port 416 nsew signal output
rlabel metal1 s 488450 0 488506 800 6 ch_out[247]
port 417 nsew signal output
rlabel metal1 s 490626 0 490682 800 6 ch_out[248]
port 418 nsew signal output
rlabel metal1 s 492802 0 492858 800 6 ch_out[249]
port 419 nsew signal output
rlabel metal1 s 26186 0 26242 800 6 ch_out[24]
port 420 nsew signal output
rlabel metal1 s 494978 0 495034 800 6 ch_out[250]
port 421 nsew signal output
rlabel metal1 s 497154 0 497210 800 6 ch_out[251]
port 422 nsew signal output
rlabel metal1 s 488722 11200 488778 12000 6 ch_out[252]
port 423 nsew signal output
rlabel metal1 s 213662 11200 213718 12000 6 ch_out[25]
port 424 nsew signal output
rlabel metal1 s 214206 11200 214262 12000 6 ch_out[26]
port 425 nsew signal output
rlabel metal1 s 29450 0 29506 800 6 ch_out[27]
port 426 nsew signal output
rlabel metal1 s 215294 11200 215350 12000 6 ch_out[28]
port 427 nsew signal output
rlabel metal1 s 215838 11200 215894 12000 6 ch_out[29]
port 428 nsew signal output
rlabel metal1 s 2250 0 2306 800 6 ch_out[2]
port 429 nsew signal output
rlabel metal1 s 32714 0 32770 800 6 ch_out[30]
port 430 nsew signal output
rlabel metal1 s 216926 11200 216982 12000 6 ch_out[31]
port 431 nsew signal output
rlabel metal1 s 217470 11200 217526 12000 6 ch_out[32]
port 432 nsew signal output
rlabel metal1 s 35978 0 36034 800 6 ch_out[33]
port 433 nsew signal output
rlabel metal1 s 218558 11200 218614 12000 6 ch_out[34]
port 434 nsew signal output
rlabel metal1 s 219102 11200 219158 12000 6 ch_out[35]
port 435 nsew signal output
rlabel metal1 s 39242 0 39298 800 6 ch_out[36]
port 436 nsew signal output
rlabel metal1 s 220190 11200 220246 12000 6 ch_out[37]
port 437 nsew signal output
rlabel metal1 s 220734 11200 220790 12000 6 ch_out[38]
port 438 nsew signal output
rlabel metal1 s 42506 0 42562 800 6 ch_out[39]
port 439 nsew signal output
rlabel metal1 s 201694 11200 201750 12000 6 ch_out[3]
port 440 nsew signal output
rlabel metal1 s 221822 11200 221878 12000 6 ch_out[40]
port 441 nsew signal output
rlabel metal1 s 222366 11200 222422 12000 6 ch_out[41]
port 442 nsew signal output
rlabel metal1 s 45770 0 45826 800 6 ch_out[42]
port 443 nsew signal output
rlabel metal1 s 223454 11200 223510 12000 6 ch_out[43]
port 444 nsew signal output
rlabel metal1 s 223998 11200 224054 12000 6 ch_out[44]
port 445 nsew signal output
rlabel metal1 s 49034 0 49090 800 6 ch_out[45]
port 446 nsew signal output
rlabel metal1 s 225086 11200 225142 12000 6 ch_out[46]
port 447 nsew signal output
rlabel metal1 s 225630 11200 225686 12000 6 ch_out[47]
port 448 nsew signal output
rlabel metal1 s 52298 0 52354 800 6 ch_out[48]
port 449 nsew signal output
rlabel metal1 s 226718 11200 226774 12000 6 ch_out[49]
port 450 nsew signal output
rlabel metal1 s 202238 11200 202294 12000 6 ch_out[4]
port 451 nsew signal output
rlabel metal1 s 227262 11200 227318 12000 6 ch_out[50]
port 452 nsew signal output
rlabel metal1 s 55562 0 55618 800 6 ch_out[51]
port 453 nsew signal output
rlabel metal1 s 228350 11200 228406 12000 6 ch_out[52]
port 454 nsew signal output
rlabel metal1 s 228894 11200 228950 12000 6 ch_out[53]
port 455 nsew signal output
rlabel metal1 s 58826 0 58882 800 6 ch_out[54]
port 456 nsew signal output
rlabel metal1 s 229982 11200 230038 12000 6 ch_out[55]
port 457 nsew signal output
rlabel metal1 s 230526 11200 230582 12000 6 ch_out[56]
port 458 nsew signal output
rlabel metal1 s 62090 0 62146 800 6 ch_out[57]
port 459 nsew signal output
rlabel metal1 s 231614 11200 231670 12000 6 ch_out[58]
port 460 nsew signal output
rlabel metal1 s 232158 11200 232214 12000 6 ch_out[59]
port 461 nsew signal output
rlabel metal1 s 202782 11200 202838 12000 6 ch_out[5]
port 462 nsew signal output
rlabel metal1 s 65354 0 65410 800 6 ch_out[60]
port 463 nsew signal output
rlabel metal1 s 233246 11200 233302 12000 6 ch_out[61]
port 464 nsew signal output
rlabel metal1 s 233790 11200 233846 12000 6 ch_out[62]
port 465 nsew signal output
rlabel metal1 s 68618 0 68674 800 6 ch_out[63]
port 466 nsew signal output
rlabel metal1 s 234878 11200 234934 12000 6 ch_out[64]
port 467 nsew signal output
rlabel metal1 s 235422 11200 235478 12000 6 ch_out[65]
port 468 nsew signal output
rlabel metal1 s 71882 0 71938 800 6 ch_out[66]
port 469 nsew signal output
rlabel metal1 s 236510 11200 236566 12000 6 ch_out[67]
port 470 nsew signal output
rlabel metal1 s 237054 11200 237110 12000 6 ch_out[68]
port 471 nsew signal output
rlabel metal1 s 75146 0 75202 800 6 ch_out[69]
port 472 nsew signal output
rlabel metal1 s 203326 11200 203382 12000 6 ch_out[6]
port 473 nsew signal output
rlabel metal1 s 238142 11200 238198 12000 6 ch_out[70]
port 474 nsew signal output
rlabel metal1 s 238686 11200 238742 12000 6 ch_out[71]
port 475 nsew signal output
rlabel metal1 s 78410 0 78466 800 6 ch_out[72]
port 476 nsew signal output
rlabel metal1 s 239774 11200 239830 12000 6 ch_out[73]
port 477 nsew signal output
rlabel metal1 s 240318 11200 240374 12000 6 ch_out[74]
port 478 nsew signal output
rlabel metal1 s 81674 0 81730 800 6 ch_out[75]
port 479 nsew signal output
rlabel metal1 s 241406 11200 241462 12000 6 ch_out[76]
port 480 nsew signal output
rlabel metal1 s 241950 11200 242006 12000 6 ch_out[77]
port 481 nsew signal output
rlabel metal1 s 84938 0 84994 800 6 ch_out[78]
port 482 nsew signal output
rlabel metal1 s 243038 11200 243094 12000 6 ch_out[79]
port 483 nsew signal output
rlabel metal1 s 203870 11200 203926 12000 6 ch_out[7]
port 484 nsew signal output
rlabel metal1 s 243582 11200 243638 12000 6 ch_out[80]
port 485 nsew signal output
rlabel metal1 s 88202 0 88258 800 6 ch_out[81]
port 486 nsew signal output
rlabel metal1 s 244670 11200 244726 12000 6 ch_out[82]
port 487 nsew signal output
rlabel metal1 s 245214 11200 245270 12000 6 ch_out[83]
port 488 nsew signal output
rlabel metal1 s 91466 0 91522 800 6 ch_out[84]
port 489 nsew signal output
rlabel metal1 s 246302 11200 246358 12000 6 ch_out[85]
port 490 nsew signal output
rlabel metal1 s 246846 11200 246902 12000 6 ch_out[86]
port 491 nsew signal output
rlabel metal1 s 94730 0 94786 800 6 ch_out[87]
port 492 nsew signal output
rlabel metal1 s 247934 11200 247990 12000 6 ch_out[88]
port 493 nsew signal output
rlabel metal1 s 248478 11200 248534 12000 6 ch_out[89]
port 494 nsew signal output
rlabel metal1 s 8778 0 8834 800 6 ch_out[8]
port 495 nsew signal output
rlabel metal1 s 97994 0 98050 800 6 ch_out[90]
port 496 nsew signal output
rlabel metal1 s 249566 11200 249622 12000 6 ch_out[91]
port 497 nsew signal output
rlabel metal1 s 250110 11200 250166 12000 6 ch_out[92]
port 498 nsew signal output
rlabel metal1 s 101258 0 101314 800 6 ch_out[93]
port 499 nsew signal output
rlabel metal1 s 251198 11200 251254 12000 6 ch_out[94]
port 500 nsew signal output
rlabel metal1 s 251742 11200 251798 12000 6 ch_out[95]
port 501 nsew signal output
rlabel metal1 s 104522 0 104578 800 6 ch_out[96]
port 502 nsew signal output
rlabel metal1 s 252830 11200 252886 12000 6 ch_out[97]
port 503 nsew signal output
rlabel metal1 s 253374 11200 253430 12000 6 ch_out[98]
port 504 nsew signal output
rlabel metal1 s 107786 0 107842 800 6 ch_out[99]
port 505 nsew signal output
rlabel metal1 s 204958 11200 205014 12000 6 ch_out[9]
port 506 nsew signal output
rlabel metal2 s -416 656 -96 11312 4 vccd1
port 507 nsew power bidirectional
rlabel metal3 s -416 656 530336 976 6 vccd1
port 507 nsew power bidirectional
rlabel metal3 s -416 10992 530336 11312 6 vccd1
port 507 nsew power bidirectional
rlabel metal2 s 530016 656 530336 11312 6 vccd1
port 507 nsew power bidirectional
rlabel metal2 s 66908 -4 67228 11972 6 vccd1
port 507 nsew power bidirectional
rlabel metal2 s 198836 -4 199156 11972 6 vccd1
port 507 nsew power bidirectional
rlabel metal2 s 330764 -4 331084 11972 6 vccd1
port 507 nsew power bidirectional
rlabel metal2 s 462692 -4 463012 11972 6 vccd1
port 507 nsew power bidirectional
rlabel metal3 s -1076 2968 530996 3288 6 vccd1
port 507 nsew power bidirectional
rlabel metal3 s -1076 4872 530996 5192 6 vccd1
port 507 nsew power bidirectional
rlabel metal3 s -1076 6776 530996 7096 6 vccd1
port 507 nsew power bidirectional
rlabel metal3 s -1076 8680 530996 9000 6 vccd1
port 507 nsew power bidirectional
rlabel metal2 s -1076 -4 -756 11972 4 vssd1
port 508 nsew ground bidirectional
rlabel metal3 s -1076 -4 530996 316 6 vssd1
port 508 nsew ground bidirectional
rlabel metal3 s -1076 11652 530996 11972 6 vssd1
port 508 nsew ground bidirectional
rlabel metal2 s 530676 -4 530996 11972 6 vssd1
port 508 nsew ground bidirectional
rlabel metal2 s 67568 -4 67888 11972 6 vssd1
port 508 nsew ground bidirectional
rlabel metal2 s 199496 -4 199816 11972 6 vssd1
port 508 nsew ground bidirectional
rlabel metal2 s 331424 -4 331744 11972 6 vssd1
port 508 nsew ground bidirectional
rlabel metal2 s 463352 -4 463672 11972 6 vssd1
port 508 nsew ground bidirectional
rlabel metal3 s -1076 3628 530996 3948 6 vssd1
port 508 nsew ground bidirectional
rlabel metal3 s -1076 5532 530996 5852 6 vssd1
port 508 nsew ground bidirectional
rlabel metal3 s -1076 7436 530996 7756 6 vssd1
port 508 nsew ground bidirectional
rlabel metal3 s -1076 9340 530996 9660 6 vssd1
port 508 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 530000 12000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2703810
string GDS_FILE /home/lx/projects/caravel_env/caravel_usb_test/openlane/bus_rep_south/runs/bus_rep_south/results/signoff/bus_rep_south.magic.gds
string GDS_START 54436
<< end >>

