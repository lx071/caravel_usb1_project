magic
tech sky130A
magscale 1 2
timestamp 1698804403
<< viali >>
rect 107853 7429 107887 7463
rect 117605 7429 117639 7463
rect 120641 7429 120675 7463
rect 213377 7429 213411 7463
rect 216045 7429 216079 7463
rect 32689 7361 32723 7395
rect 33241 7361 33275 7395
rect 33517 7361 33551 7395
rect 35265 7361 35299 7395
rect 36829 7361 36863 7395
rect 37473 7361 37507 7395
rect 56609 7361 56643 7395
rect 57069 7361 57103 7395
rect 57345 7361 57379 7395
rect 59369 7361 59403 7395
rect 60933 7361 60967 7395
rect 61485 7361 61519 7395
rect 63509 7361 63543 7395
rect 64797 7361 64831 7395
rect 65901 7361 65935 7395
rect 66453 7361 66487 7395
rect 71973 7361 72007 7395
rect 72525 7361 72559 7395
rect 72801 7361 72835 7395
rect 74089 7361 74123 7395
rect 74641 7361 74675 7395
rect 74917 7361 74951 7395
rect 76113 7361 76147 7395
rect 76665 7361 76699 7395
rect 76941 7361 76975 7395
rect 78045 7361 78079 7395
rect 78781 7361 78815 7395
rect 80069 7361 80103 7395
rect 104633 7361 104667 7395
rect 105277 7361 105311 7395
rect 105829 7361 105863 7395
rect 107301 7361 107335 7395
rect 110153 7361 110187 7395
rect 110797 7361 110831 7395
rect 117881 7361 117915 7395
rect 119261 7361 119295 7395
rect 120089 7361 120123 7395
rect 121469 7361 121503 7395
rect 121837 7361 121871 7395
rect 122849 7361 122883 7395
rect 123217 7361 123251 7395
rect 123861 7361 123895 7395
rect 125333 7361 125367 7395
rect 125977 7361 126011 7395
rect 151185 7361 151219 7395
rect 153485 7361 153519 7395
rect 154773 7361 154807 7395
rect 166457 7361 166491 7395
rect 168205 7361 168239 7395
rect 168941 7361 168975 7395
rect 170137 7361 170171 7395
rect 197921 7361 197955 7395
rect 198565 7361 198599 7395
rect 200129 7361 200163 7395
rect 200773 7361 200807 7395
rect 214021 7361 214055 7395
rect 217241 7361 217275 7395
rect 219725 7361 219759 7395
rect 244381 7361 244415 7395
rect 244933 7361 244967 7395
rect 260389 7361 260423 7395
rect 35541 7293 35575 7327
rect 37749 7293 37783 7327
rect 59645 7293 59679 7327
rect 61761 7293 61795 7327
rect 63785 7293 63819 7327
rect 65073 7293 65107 7327
rect 66729 7293 66763 7327
rect 79333 7293 79367 7327
rect 80621 7293 80655 7327
rect 111349 7293 111383 7327
rect 118709 7293 118743 7327
rect 124413 7293 124447 7327
rect 126529 7293 126563 7327
rect 151737 7293 151771 7327
rect 154037 7293 154071 7327
rect 155325 7293 155359 7327
rect 167009 7293 167043 7327
rect 169493 7293 169527 7327
rect 170689 7293 170723 7327
rect 199117 7293 199151 7327
rect 201325 7293 201359 7327
rect 214573 7293 214607 7327
rect 218529 7293 218563 7327
rect 245485 7293 245519 7327
rect 260757 7293 260791 7327
rect 58817 7225 58851 7259
rect 259745 7225 259779 7259
rect 152749 7157 152783 7191
rect 217885 7157 217919 7191
rect 220461 7157 220495 7191
rect 166273 6953 166307 6987
rect 169953 6953 169987 6987
rect 35173 6885 35207 6919
rect 64613 6885 64647 6919
rect 107117 6885 107151 6919
rect 118985 6885 119019 6919
rect 122941 6885 122975 6919
rect 151001 6885 151035 6919
rect 154589 6885 154623 6919
rect 119629 6817 119663 6851
rect 123493 6817 123527 6851
rect 63325 6749 63359 6783
rect 79793 6749 79827 6783
rect 81541 6749 81575 6783
rect 108497 6749 108531 6783
rect 109141 6749 109175 6783
rect 116685 6749 116719 6783
rect 120181 6749 120215 6783
rect 121377 6749 121411 6783
rect 124045 6749 124079 6783
rect 125241 6749 125275 6783
rect 125885 6749 125919 6783
rect 156429 6749 156463 6783
rect 171655 6749 171689 6783
rect 215999 6749 216033 6783
rect 218713 6749 218747 6783
rect 246773 6749 246807 6783
rect 262045 6749 262079 6783
rect 82093 6681 82127 6715
rect 109693 6681 109727 6715
rect 116133 6681 116167 6715
rect 120825 6681 120859 6715
rect 124689 6681 124723 6715
rect 156981 6681 157015 6715
rect 172253 6681 172287 6715
rect 216597 6681 216631 6715
rect 217517 6681 217551 6715
rect 247325 6681 247359 6715
rect 262597 6681 262631 6715
rect 117421 6613 117455 6647
rect 117973 6613 118007 6647
rect 155785 6613 155819 6647
rect 171057 6613 171091 6647
rect 215493 6613 215527 6647
rect 219265 6613 219299 6647
rect 246129 6613 246163 6647
rect 307493 6409 307527 6443
rect 111165 6341 111199 6375
rect 123769 6341 123803 6375
rect 124321 6341 124355 6375
rect 353585 6341 353619 6375
rect 111809 6273 111843 6307
rect 122573 6273 122607 6307
rect 123033 6273 123067 6307
rect 126989 6273 127023 6307
rect 202429 6273 202463 6307
rect 213469 6273 213503 6307
rect 214665 6273 214699 6307
rect 215861 6273 215895 6307
rect 217885 6273 217919 6307
rect 292773 6273 292807 6307
rect 308137 6273 308171 6307
rect 310897 6273 310931 6307
rect 311725 6273 311759 6307
rect 313197 6273 313231 6307
rect 338865 6273 338899 6307
rect 354229 6273 354263 6307
rect 112361 6205 112395 6239
rect 127541 6205 127575 6239
rect 201693 6205 201727 6239
rect 202797 6205 202831 6239
rect 212917 6205 212951 6239
rect 214113 6205 214147 6239
rect 215309 6205 215343 6239
rect 217149 6205 217183 6239
rect 218437 6205 218471 6239
rect 261769 6205 261803 6239
rect 293325 6205 293359 6239
rect 308689 6205 308723 6239
rect 312369 6205 312403 6239
rect 339417 6205 339451 6239
rect 354597 6205 354631 6239
rect 126345 6137 126379 6171
rect 292129 6137 292163 6171
rect 81265 6069 81299 6103
rect 119353 6069 119387 6103
rect 120457 6069 120491 6103
rect 121469 6069 121503 6103
rect 122021 6069 122055 6103
rect 216505 6069 216539 6103
rect 313749 6069 313783 6103
rect 338221 6069 338255 6103
rect 172069 5729 172103 5763
rect 293693 5729 293727 5763
rect 310069 5729 310103 5763
rect 115029 5661 115063 5695
rect 115673 5661 115707 5695
rect 156705 5661 156739 5695
rect 157349 5661 157383 5695
rect 172713 5661 172747 5695
rect 211537 5661 211571 5695
rect 212089 5661 212123 5695
rect 247601 5661 247635 5695
rect 248153 5661 248187 5695
rect 262965 5661 262999 5695
rect 263517 5661 263551 5695
rect 294245 5661 294279 5695
rect 310897 5661 310931 5695
rect 114477 5593 114511 5627
rect 157901 5593 157935 5627
rect 173265 5593 173299 5627
rect 248981 5593 249015 5627
rect 264345 5593 264379 5627
rect 295073 5593 295107 5627
rect 122481 5525 122515 5559
rect 212733 5525 212767 5559
rect 213745 5525 213779 5559
rect 215309 5525 215343 5559
rect 311909 5525 311943 5559
rect 401149 5321 401183 5355
rect 203349 5185 203383 5219
rect 218621 5185 218655 5219
rect 309333 5185 309367 5219
rect 339877 5185 339911 5219
rect 354873 5185 354907 5219
rect 355333 5185 355367 5219
rect 386245 5185 386279 5219
rect 401701 5185 401735 5219
rect 406669 5185 406703 5219
rect 432153 5185 432187 5219
rect 432613 5185 432647 5219
rect 447977 5185 448011 5219
rect 202705 5117 202739 5151
rect 203901 5117 203935 5151
rect 219173 5117 219207 5151
rect 308781 5117 308815 5151
rect 309977 5117 310011 5151
rect 311081 5117 311115 5151
rect 340705 5117 340739 5151
rect 355977 5117 356011 5151
rect 387073 5117 387107 5151
rect 402529 5117 402563 5151
rect 406117 5117 406151 5151
rect 433257 5117 433291 5151
rect 448805 5117 448839 5151
rect 385693 5049 385727 5083
rect 218069 4981 218103 5015
rect 339325 4981 339359 5015
rect 407313 4981 407347 5015
rect 447425 4981 447459 5015
rect 248705 4777 248739 4811
rect 264069 4777 264103 4811
rect 112637 4573 112671 4607
rect 113189 4573 113223 4607
rect 210709 4573 210743 4607
rect 249349 4573 249383 4607
rect 264713 4573 264747 4607
rect 294797 4573 294831 4607
rect 295441 4573 295475 4607
rect 308597 4573 308631 4607
rect 309517 4573 309551 4607
rect 311081 4573 311115 4607
rect 405197 4573 405231 4607
rect 112361 4505 112395 4539
rect 210157 4505 210191 4539
rect 249717 4505 249751 4539
rect 265265 4505 265299 4539
rect 295993 4505 296027 4539
rect 308045 4505 308079 4539
rect 310345 4505 310379 4539
rect 311633 4505 311667 4539
rect 404645 4505 404679 4539
rect 211353 4437 211387 4471
rect 405933 4437 405967 4471
rect 309333 4233 309367 4267
rect 310805 4165 310839 4199
rect 499957 4165 499991 4199
rect 306481 4097 306515 4131
rect 341533 4097 341567 4131
rect 356897 4097 356931 4131
rect 387809 4097 387843 4131
rect 403265 4097 403299 4131
rect 434177 4097 434211 4131
rect 448989 4097 449023 4131
rect 449633 4097 449667 4131
rect 480545 4097 480579 4131
rect 496001 4097 496035 4131
rect 500509 4097 500543 4131
rect 526913 4097 526947 4131
rect 305929 4029 305963 4063
rect 342729 4029 342763 4063
rect 356253 4029 356287 4063
rect 358093 4029 358127 4063
rect 389005 4029 389039 4063
rect 404461 4029 404495 4063
rect 435373 4029 435407 4063
rect 450829 4029 450863 4063
rect 481741 4029 481775 4063
rect 497197 4029 497231 4063
rect 526269 4029 526303 4063
rect 528109 4029 528143 4063
rect 433533 3961 433567 3995
rect 307125 3893 307159 3927
rect 308873 3893 308907 3927
rect 387165 3893 387199 3927
rect 402621 3893 402655 3927
rect 479901 3893 479935 3927
rect 495449 3893 495483 3927
rect 501245 3893 501279 3927
rect 341349 3553 341383 3587
rect 208409 3485 208443 3519
rect 208961 3485 208995 3519
rect 402805 3485 402839 3519
rect 404185 3485 404219 3519
rect 404829 3485 404863 3519
rect 499221 3485 499255 3519
rect 541909 3485 541943 3519
rect 208133 3417 208167 3451
rect 402253 3417 402287 3451
rect 403633 3417 403667 3451
rect 498669 3417 498703 3451
rect 543105 3417 543139 3451
rect 499865 3349 499899 3383
rect 541357 3349 541391 3383
rect 32505 3145 32539 3179
rect 202521 3145 202555 3179
rect 295349 3145 295383 3179
rect 305469 3145 305503 3179
rect 449909 3145 449943 3179
rect 542553 3145 542587 3179
rect 573465 3145 573499 3179
rect 588921 3145 588955 3179
rect 619833 3145 619867 3179
rect 635289 3145 635323 3179
rect 109785 3077 109819 3111
rect 264345 3077 264379 3111
rect 357081 3077 357115 3111
rect 387993 3077 388027 3111
rect 434361 3077 434395 3111
rect 527189 3077 527223 3111
rect 594073 3077 594107 3111
rect 125241 3009 125275 3043
rect 218069 3009 218103 3043
rect 304641 3009 304675 3043
rect 401057 3009 401091 3043
rect 496185 3009 496219 3043
rect 497289 3009 497323 3043
rect 497565 3009 497599 3043
rect 594349 3009 594383 3043
rect 78873 2941 78907 2975
rect 171609 2941 171643 2975
rect 304365 2941 304399 2975
rect 310713 2941 310747 2975
rect 400781 2941 400815 2975
rect 403357 2941 403391 2975
rect 63509 2873 63543 2907
rect 156153 2873 156187 2907
rect 1593 2805 1627 2839
rect 47961 2805 47995 2839
rect 94329 2805 94363 2839
rect 140789 2805 140823 2839
rect 186881 2805 186915 2839
rect 233525 2805 233559 2839
rect 248889 2805 248923 2839
rect 279617 2805 279651 2839
rect 326261 2805 326295 2839
rect 341717 2805 341751 2839
rect 372629 2805 372663 2839
rect 401609 2805 401643 2839
rect 465273 2805 465307 2839
rect 480729 2805 480763 2839
rect 558009 2805 558043 2839
rect 18061 2601 18095 2635
rect 419365 2601 419399 2635
rect 512101 2601 512135 2635
rect 604837 2601 604871 2635
rect 94605 2533 94639 2567
rect 233617 2533 233651 2567
rect 326353 2533 326387 2567
rect 187157 2465 187191 2499
rect 279893 2465 279927 2499
rect 402621 2465 402655 2499
rect 2053 2397 2087 2431
rect 17509 2397 17543 2431
rect 32965 2397 32999 2431
rect 48421 2397 48455 2431
rect 63877 2397 63911 2431
rect 79333 2397 79367 2431
rect 94789 2397 94823 2431
rect 110245 2397 110279 2431
rect 125701 2397 125735 2431
rect 156613 2397 156647 2431
rect 172069 2397 172103 2431
rect 202981 2397 203015 2431
rect 218437 2397 218471 2431
rect 249349 2397 249383 2431
rect 264805 2397 264839 2431
rect 295717 2397 295751 2431
rect 311173 2397 311207 2431
rect 342085 2397 342119 2431
rect 357541 2397 357575 2431
rect 372997 2397 373031 2431
rect 388453 2397 388487 2431
rect 403909 2397 403943 2431
rect 419181 2397 419215 2431
rect 419825 2397 419859 2431
rect 434821 2397 434855 2431
rect 450277 2397 450311 2431
rect 465733 2397 465767 2431
rect 481189 2397 481223 2431
rect 496645 2397 496679 2431
rect 511917 2397 511951 2431
rect 512561 2397 512595 2431
rect 527557 2397 527591 2431
rect 543013 2397 543047 2431
rect 558469 2397 558503 2431
rect 573925 2397 573959 2431
rect 589381 2397 589415 2431
rect 604653 2397 604687 2431
rect 605297 2397 605331 2431
rect 620293 2397 620327 2431
rect 635749 2397 635783 2431
rect 140881 2329 140915 2363
rect 141065 2329 141099 2363
rect 187433 2329 187467 2363
rect 233801 2329 233835 2363
rect 280169 2329 280203 2363
rect 326537 2329 326571 2363
rect 1869 2261 1903 2295
rect 17325 2261 17359 2295
rect 32781 2261 32815 2295
rect 48237 2261 48271 2295
rect 63693 2261 63727 2295
rect 79149 2261 79183 2295
rect 110061 2261 110095 2295
rect 125517 2261 125551 2295
rect 156429 2261 156463 2295
rect 171885 2261 171919 2295
rect 202797 2261 202831 2295
rect 218253 2261 218287 2295
rect 249165 2261 249199 2295
rect 264621 2261 264655 2295
rect 295533 2261 295567 2295
rect 310989 2261 311023 2295
rect 341901 2261 341935 2295
rect 357357 2261 357391 2295
rect 372813 2261 372847 2295
rect 388269 2261 388303 2295
rect 403725 2261 403759 2295
rect 434637 2261 434671 2295
rect 450093 2261 450127 2295
rect 465549 2261 465583 2295
rect 481005 2261 481039 2295
rect 496461 2261 496495 2295
rect 527373 2261 527407 2295
rect 542829 2261 542863 2295
rect 558285 2261 558319 2295
rect 573741 2261 573775 2295
rect 589197 2261 589231 2295
rect 620109 2261 620143 2295
rect 635565 2261 635599 2295
<< metal1 >>
rect 19702 9188 19708 9240
rect 19760 9228 19766 9240
rect 20066 9228 20122 10000
rect 19760 9200 20122 9228
rect 19760 9188 19766 9200
rect 20162 9188 20168 9240
rect 20220 9228 20226 9240
rect 20338 9228 20394 10000
rect 20610 9228 20666 10000
rect 20220 9200 20394 9228
rect 20548 9200 20666 9228
rect 20882 9228 20938 10000
rect 20990 9228 20996 9240
rect 20882 9200 20996 9228
rect 20220 9188 20226 9200
rect 20548 9160 20576 9200
rect 20990 9188 20996 9200
rect 21048 9188 21054 9240
rect 21154 9228 21210 10000
rect 21266 9228 21272 9240
rect 21154 9200 21272 9228
rect 21266 9188 21272 9200
rect 21324 9188 21330 9240
rect 21426 9228 21482 10000
rect 21376 9200 21482 9228
rect 21698 9228 21754 10000
rect 21970 9228 22026 10000
rect 22242 9228 22298 10000
rect 22514 9228 22570 10000
rect 22786 9228 22842 10000
rect 22922 9228 22928 9240
rect 21698 9200 21772 9228
rect 21970 9200 22048 9228
rect 22242 9200 22324 9228
rect 22514 9200 22600 9228
rect 22786 9200 22928 9228
rect 21376 9160 21404 9200
rect 21744 9160 21772 9200
rect 22020 9160 22048 9200
rect 22296 9160 22324 9200
rect 22572 9160 22600 9200
rect 22922 9188 22928 9200
rect 22980 9188 22986 9240
rect 23058 9228 23114 10000
rect 23198 9228 23204 9240
rect 23058 9200 23204 9228
rect 23198 9188 23204 9200
rect 23256 9188 23262 9240
rect 23330 9228 23386 10000
rect 23602 9228 23658 10000
rect 23750 9228 23756 9240
rect 23330 9200 23428 9228
rect 23602 9200 23756 9228
rect 23400 9172 23428 9200
rect 23750 9188 23756 9200
rect 23808 9188 23814 9240
rect 23874 9228 23930 10000
rect 24146 9228 24202 10000
rect 24302 9228 24308 9240
rect 23874 9200 23980 9228
rect 24146 9200 24308 9228
rect 20548 9132 20652 9160
rect 21376 9132 21468 9160
rect 20624 8900 20652 9132
rect 20622 8848 20628 8900
rect 20680 8848 20686 8900
rect 21440 8888 21468 9132
rect 21698 9132 21772 9160
rect 21974 9132 22048 9160
rect 22250 9132 22324 9160
rect 22526 9132 22600 9160
rect 21698 8956 21726 9132
rect 21974 8968 22002 9132
rect 21818 8956 21824 8968
rect 21698 8928 21824 8956
rect 21818 8916 21824 8928
rect 21876 8916 21882 8968
rect 21974 8928 22008 8968
rect 22002 8916 22008 8928
rect 22060 8916 22066 8968
rect 21910 8888 21916 8900
rect 21440 8860 21916 8888
rect 21910 8848 21916 8860
rect 21968 8848 21974 8900
rect 22250 8412 22278 9132
rect 22526 8956 22554 9132
rect 23382 9120 23388 9172
rect 23440 9120 23446 9172
rect 23952 9160 23980 9200
rect 24302 9188 24308 9200
rect 24360 9188 24366 9240
rect 24418 9228 24474 10000
rect 24578 9228 24584 9240
rect 24418 9200 24584 9228
rect 24578 9188 24584 9200
rect 24636 9188 24642 9240
rect 24690 9228 24746 10000
rect 24962 9228 25018 10000
rect 25130 9228 25136 9240
rect 24690 9200 24808 9228
rect 24962 9200 25136 9228
rect 24780 9172 24808 9200
rect 25130 9188 25136 9200
rect 25188 9188 25194 9240
rect 25234 9228 25290 10000
rect 25506 9228 25562 10000
rect 25682 9228 25688 9240
rect 25234 9200 25360 9228
rect 25506 9200 25688 9228
rect 23888 9132 23980 9160
rect 23290 8956 23296 8968
rect 22526 8928 23296 8956
rect 23290 8916 23296 8928
rect 23348 8916 23354 8968
rect 23888 8616 23916 9132
rect 24762 9120 24768 9172
rect 24820 9120 24826 9172
rect 25332 9160 25360 9200
rect 25682 9188 25688 9200
rect 25740 9188 25746 9240
rect 25778 9228 25834 10000
rect 25958 9228 25964 9240
rect 25778 9200 25964 9228
rect 25958 9188 25964 9200
rect 26016 9188 26022 9240
rect 26050 9228 26106 10000
rect 26142 9228 26148 9240
rect 26050 9200 26148 9228
rect 26142 9188 26148 9200
rect 26200 9188 26206 9240
rect 26322 9228 26378 10000
rect 26252 9200 26378 9228
rect 26594 9228 26650 10000
rect 26694 9228 26700 9240
rect 26594 9200 26700 9228
rect 25240 9132 25360 9160
rect 26252 9160 26280 9200
rect 26694 9188 26700 9200
rect 26752 9188 26758 9240
rect 26866 9228 26922 10000
rect 26804 9200 26922 9228
rect 27138 9228 27194 10000
rect 27246 9228 27252 9240
rect 27138 9200 27252 9228
rect 26804 9160 26832 9200
rect 27246 9188 27252 9200
rect 27304 9188 27310 9240
rect 27410 9228 27466 10000
rect 27522 9228 27528 9240
rect 27410 9200 27528 9228
rect 27522 9188 27528 9200
rect 27580 9188 27586 9240
rect 27682 9228 27738 10000
rect 27798 9228 27804 9240
rect 27682 9200 27804 9228
rect 27798 9188 27804 9200
rect 27856 9188 27862 9240
rect 27954 9228 28010 10000
rect 28074 9228 28080 9240
rect 27954 9200 28080 9228
rect 28074 9188 28080 9200
rect 28132 9188 28138 9240
rect 28226 9228 28282 10000
rect 28350 9228 28356 9240
rect 28226 9200 28356 9228
rect 28350 9188 28356 9200
rect 28408 9188 28414 9240
rect 28498 9228 28554 10000
rect 28770 9228 28826 10000
rect 28902 9228 28908 9240
rect 28498 9200 28672 9228
rect 28770 9200 28908 9228
rect 28644 9160 28672 9200
rect 28902 9188 28908 9200
rect 28960 9188 28966 9240
rect 29042 9228 29098 10000
rect 29178 9228 29184 9240
rect 29042 9200 29184 9228
rect 29178 9188 29184 9200
rect 29236 9188 29242 9240
rect 29314 9228 29370 10000
rect 29454 9228 29460 9240
rect 29314 9200 29460 9228
rect 29454 9188 29460 9200
rect 29512 9188 29518 9240
rect 29586 9228 29642 10000
rect 29730 9228 29736 9240
rect 29586 9200 29736 9228
rect 29730 9188 29736 9200
rect 29788 9188 29794 9240
rect 29858 9228 29914 10000
rect 30006 9228 30012 9240
rect 29858 9200 30012 9228
rect 30006 9188 30012 9200
rect 30064 9188 30070 9240
rect 30130 9228 30186 10000
rect 30402 9228 30458 10000
rect 30674 9228 30730 10000
rect 30834 9228 30840 9240
rect 30130 9200 30328 9228
rect 30402 9200 30604 9228
rect 30674 9200 30840 9228
rect 30098 9160 30104 9172
rect 26252 9132 26372 9160
rect 26804 9132 26908 9160
rect 28644 9132 30104 9160
rect 25240 8956 25268 9132
rect 25240 8928 26280 8956
rect 26252 8684 26280 8928
rect 26344 8820 26372 9132
rect 26880 8956 26908 9132
rect 30098 9120 30104 9132
rect 30156 9120 30162 9172
rect 30300 9160 30328 9200
rect 30466 9160 30472 9172
rect 30300 9132 30472 9160
rect 30466 9120 30472 9132
rect 30524 9120 30530 9172
rect 30576 9160 30604 9200
rect 30834 9188 30840 9200
rect 30892 9188 30898 9240
rect 30946 9228 31002 10000
rect 31110 9228 31116 9240
rect 30946 9200 31116 9228
rect 31110 9188 31116 9200
rect 31168 9188 31174 9240
rect 31218 9228 31274 10000
rect 31478 9228 31484 9240
rect 31218 9200 31484 9228
rect 31478 9188 31484 9200
rect 31536 9188 31542 9240
rect 118970 9160 118976 9172
rect 30576 9132 118976 9160
rect 118970 9120 118976 9132
rect 119028 9120 119034 9172
rect 30282 9052 30288 9104
rect 30340 9092 30346 9104
rect 110138 9092 110144 9104
rect 30340 9064 110144 9092
rect 30340 9052 30346 9064
rect 110138 9052 110144 9064
rect 110196 9052 110202 9104
rect 108482 9024 108488 9036
rect 30300 8996 108488 9024
rect 30300 8956 30328 8996
rect 108482 8984 108488 8996
rect 108540 8984 108546 9036
rect 26880 8928 30328 8956
rect 30374 8916 30380 8968
rect 30432 8956 30438 8968
rect 107286 8956 107292 8968
rect 30432 8928 107292 8956
rect 30432 8916 30438 8928
rect 107286 8916 107292 8928
rect 107344 8916 107350 8968
rect 30466 8848 30472 8900
rect 30524 8888 30530 8900
rect 104618 8888 104624 8900
rect 30524 8860 104624 8888
rect 30524 8848 30530 8860
rect 104618 8848 104624 8860
rect 104676 8848 104682 8900
rect 78030 8820 78036 8832
rect 26344 8792 78036 8820
rect 78030 8780 78036 8792
rect 78088 8780 78094 8832
rect 29730 8712 29736 8764
rect 29788 8752 29794 8764
rect 74074 8752 74080 8764
rect 29788 8724 74080 8752
rect 29788 8712 29794 8724
rect 74074 8712 74080 8724
rect 74132 8712 74138 8764
rect 30282 8684 30288 8696
rect 26252 8656 30288 8684
rect 30282 8644 30288 8656
rect 30340 8644 30346 8696
rect 30374 8644 30380 8696
rect 30432 8684 30438 8696
rect 62574 8684 62580 8696
rect 30432 8656 62580 8684
rect 30432 8644 30438 8656
rect 62574 8644 62580 8656
rect 62632 8644 62638 8696
rect 35250 8616 35256 8628
rect 23888 8588 30328 8616
rect 26142 8508 26148 8560
rect 26200 8548 26206 8560
rect 30190 8548 30196 8560
rect 26200 8520 30196 8548
rect 26200 8508 26206 8520
rect 30190 8508 30196 8520
rect 30248 8508 30254 8560
rect 30300 8548 30328 8588
rect 30576 8588 35256 8616
rect 30576 8548 30604 8588
rect 35250 8576 35256 8588
rect 35308 8576 35314 8628
rect 36814 8616 36820 8628
rect 35866 8588 36820 8616
rect 30300 8520 30604 8548
rect 30650 8508 30656 8560
rect 30708 8548 30714 8560
rect 35866 8548 35894 8588
rect 36814 8576 36820 8588
rect 36872 8576 36878 8628
rect 30708 8520 35894 8548
rect 30708 8508 30714 8520
rect 25682 8440 25688 8492
rect 25740 8480 25746 8492
rect 32674 8480 32680 8492
rect 25740 8452 32680 8480
rect 25740 8440 25746 8452
rect 32674 8440 32680 8452
rect 32732 8440 32738 8492
rect 22250 8384 27200 8412
rect 27172 8276 27200 8384
rect 27246 8372 27252 8424
rect 27304 8412 27310 8424
rect 123846 8412 123852 8424
rect 27304 8384 123852 8412
rect 27304 8372 27310 8384
rect 123846 8372 123852 8384
rect 123904 8372 123910 8424
rect 30650 8276 30656 8288
rect 27172 8248 30656 8276
rect 30650 8236 30656 8248
rect 30708 8236 30714 8288
rect 57330 8236 57336 8288
rect 57388 8276 57394 8288
rect 151170 8276 151176 8288
rect 57388 8248 151176 8276
rect 57388 8236 57394 8248
rect 151170 8236 151176 8248
rect 151228 8236 151234 8288
rect 74902 8168 74908 8220
rect 74960 8208 74966 8220
rect 168190 8208 168196 8220
rect 74960 8180 168196 8208
rect 74960 8168 74966 8180
rect 168190 8168 168196 8180
rect 168248 8168 168254 8220
rect 22922 8100 22928 8152
rect 22980 8140 22986 8152
rect 65886 8140 65892 8152
rect 22980 8112 65892 8140
rect 22980 8100 22986 8112
rect 65886 8100 65892 8112
rect 65944 8100 65950 8152
rect 72786 8100 72792 8152
rect 72844 8140 72850 8152
rect 166442 8140 166448 8152
rect 72844 8112 166448 8140
rect 72844 8100 72850 8112
rect 166442 8100 166448 8112
rect 166500 8100 166506 8152
rect 28074 8032 28080 8084
rect 28132 8072 28138 8084
rect 76098 8072 76104 8084
rect 28132 8044 76104 8072
rect 28132 8032 28138 8044
rect 76098 8032 76104 8044
rect 76156 8032 76162 8084
rect 24762 7964 24768 8016
rect 24820 8004 24826 8016
rect 79962 8004 79968 8016
rect 24820 7976 79968 8004
rect 24820 7964 24826 7976
rect 79962 7964 79968 7976
rect 80020 7964 80026 8016
rect 31110 7896 31116 7948
rect 31168 7936 31174 7948
rect 56594 7936 56600 7948
rect 31168 7908 56600 7936
rect 31168 7896 31174 7908
rect 56594 7896 56600 7908
rect 56652 7896 56658 7948
rect 76926 7896 76932 7948
rect 76984 7936 76990 7948
rect 170122 7936 170128 7948
rect 76984 7908 170128 7936
rect 76984 7896 76990 7908
rect 170122 7896 170128 7908
rect 170180 7896 170186 7948
rect 33502 7828 33508 7880
rect 33560 7868 33566 7880
rect 125318 7868 125324 7880
rect 33560 7840 125324 7868
rect 33560 7828 33566 7840
rect 125318 7828 125324 7840
rect 125376 7828 125382 7880
rect 27798 7760 27804 7812
rect 27856 7800 27862 7812
rect 60918 7800 60924 7812
rect 27856 7772 60924 7800
rect 27856 7760 27862 7772
rect 60918 7760 60924 7772
rect 60976 7760 60982 7812
rect 107838 7760 107844 7812
rect 107896 7800 107902 7812
rect 200114 7800 200120 7812
rect 107896 7772 200120 7800
rect 107896 7760 107902 7772
rect 200114 7760 200120 7772
rect 200172 7760 200178 7812
rect 31478 7692 31484 7744
rect 31536 7732 31542 7744
rect 71958 7732 71964 7744
rect 31536 7704 71964 7732
rect 31536 7692 31542 7704
rect 71958 7692 71964 7704
rect 72016 7692 72022 7744
rect 105814 7692 105820 7744
rect 105872 7732 105878 7744
rect 197906 7732 197912 7744
rect 105872 7704 197912 7732
rect 105872 7692 105878 7704
rect 197906 7692 197912 7704
rect 197964 7692 197970 7744
rect 1104 7642 648876 7664
rect 1104 7590 82581 7642
rect 82633 7590 82645 7642
rect 82697 7590 82709 7642
rect 82761 7590 82773 7642
rect 82825 7590 82837 7642
rect 82889 7590 244524 7642
rect 244576 7590 244588 7642
rect 244640 7590 244652 7642
rect 244704 7590 244716 7642
rect 244768 7590 244780 7642
rect 244832 7590 406467 7642
rect 406519 7590 406531 7642
rect 406583 7590 406595 7642
rect 406647 7590 406659 7642
rect 406711 7590 406723 7642
rect 406775 7590 568410 7642
rect 568462 7590 568474 7642
rect 568526 7590 568538 7642
rect 568590 7590 568602 7642
rect 568654 7590 568666 7642
rect 568718 7590 648876 7642
rect 1104 7568 648876 7590
rect 25130 7488 25136 7540
rect 25188 7528 25194 7540
rect 25188 7500 117636 7528
rect 25188 7488 25194 7500
rect 25958 7420 25964 7472
rect 26016 7460 26022 7472
rect 26016 7432 107792 7460
rect 26016 7420 26022 7432
rect 32674 7352 32680 7404
rect 32732 7392 32738 7404
rect 33229 7395 33287 7401
rect 33229 7392 33241 7395
rect 32732 7364 33241 7392
rect 32732 7352 32738 7364
rect 33229 7361 33241 7364
rect 33275 7361 33287 7395
rect 33229 7355 33287 7361
rect 33502 7352 33508 7404
rect 33560 7352 33566 7404
rect 35250 7352 35256 7404
rect 35308 7352 35314 7404
rect 36814 7352 36820 7404
rect 36872 7392 36878 7404
rect 37461 7395 37519 7401
rect 37461 7392 37473 7395
rect 36872 7364 37473 7392
rect 36872 7352 36878 7364
rect 37461 7361 37473 7364
rect 37507 7361 37519 7395
rect 37461 7355 37519 7361
rect 56594 7352 56600 7404
rect 56652 7392 56658 7404
rect 57057 7395 57115 7401
rect 57057 7392 57069 7395
rect 56652 7364 57069 7392
rect 56652 7352 56658 7364
rect 57057 7361 57069 7364
rect 57103 7361 57115 7395
rect 57057 7355 57115 7361
rect 57330 7352 57336 7404
rect 57388 7352 57394 7404
rect 59357 7395 59415 7401
rect 59357 7392 59369 7395
rect 58820 7364 59369 7392
rect 35526 7284 35532 7336
rect 35584 7284 35590 7336
rect 37734 7284 37740 7336
rect 37792 7284 37798 7336
rect 29454 7216 29460 7268
rect 29512 7256 29518 7268
rect 58820 7265 58848 7364
rect 59357 7361 59369 7364
rect 59403 7361 59415 7395
rect 59357 7355 59415 7361
rect 60918 7352 60924 7404
rect 60976 7392 60982 7404
rect 61473 7395 61531 7401
rect 61473 7392 61485 7395
rect 60976 7364 61485 7392
rect 60976 7352 60982 7364
rect 61473 7361 61485 7364
rect 61519 7361 61531 7395
rect 61473 7355 61531 7361
rect 62574 7352 62580 7404
rect 62632 7392 62638 7404
rect 63034 7392 63040 7404
rect 62632 7364 63040 7392
rect 62632 7352 62638 7364
rect 63034 7352 63040 7364
rect 63092 7392 63098 7404
rect 63497 7395 63555 7401
rect 63497 7392 63509 7395
rect 63092 7364 63509 7392
rect 63092 7352 63098 7364
rect 63497 7361 63509 7364
rect 63543 7361 63555 7395
rect 63497 7355 63555 7361
rect 64782 7352 64788 7404
rect 64840 7352 64846 7404
rect 65886 7352 65892 7404
rect 65944 7392 65950 7404
rect 66441 7395 66499 7401
rect 66441 7392 66453 7395
rect 65944 7364 66453 7392
rect 65944 7352 65950 7364
rect 66441 7361 66453 7364
rect 66487 7361 66499 7395
rect 66441 7355 66499 7361
rect 71958 7352 71964 7404
rect 72016 7392 72022 7404
rect 72513 7395 72571 7401
rect 72513 7392 72525 7395
rect 72016 7364 72525 7392
rect 72016 7352 72022 7364
rect 72513 7361 72525 7364
rect 72559 7361 72571 7395
rect 72513 7355 72571 7361
rect 72786 7352 72792 7404
rect 72844 7352 72850 7404
rect 74074 7352 74080 7404
rect 74132 7392 74138 7404
rect 74629 7395 74687 7401
rect 74629 7392 74641 7395
rect 74132 7364 74641 7392
rect 74132 7352 74138 7364
rect 74629 7361 74641 7364
rect 74675 7361 74687 7395
rect 74629 7355 74687 7361
rect 74902 7352 74908 7404
rect 74960 7352 74966 7404
rect 76098 7352 76104 7404
rect 76156 7392 76162 7404
rect 76653 7395 76711 7401
rect 76653 7392 76665 7395
rect 76156 7364 76665 7392
rect 76156 7352 76162 7364
rect 76653 7361 76665 7364
rect 76699 7361 76711 7395
rect 76653 7355 76711 7361
rect 76926 7352 76932 7404
rect 76984 7352 76990 7404
rect 78030 7352 78036 7404
rect 78088 7392 78094 7404
rect 78769 7395 78827 7401
rect 78769 7392 78781 7395
rect 78088 7364 78781 7392
rect 78088 7352 78094 7364
rect 78769 7361 78781 7364
rect 78815 7361 78827 7395
rect 78769 7355 78827 7361
rect 79594 7352 79600 7404
rect 79652 7392 79658 7404
rect 79962 7392 79968 7404
rect 79652 7364 79968 7392
rect 79652 7352 79658 7364
rect 79962 7352 79968 7364
rect 80020 7392 80026 7404
rect 80057 7395 80115 7401
rect 80057 7392 80069 7395
rect 80020 7364 80069 7392
rect 80020 7352 80026 7364
rect 80057 7361 80069 7364
rect 80103 7361 80115 7395
rect 80057 7355 80115 7361
rect 104618 7352 104624 7404
rect 104676 7392 104682 7404
rect 105265 7395 105323 7401
rect 105265 7392 105277 7395
rect 104676 7364 105277 7392
rect 104676 7352 104682 7364
rect 105265 7361 105277 7364
rect 105311 7361 105323 7395
rect 105265 7355 105323 7361
rect 105814 7352 105820 7404
rect 105872 7352 105878 7404
rect 107286 7352 107292 7404
rect 107344 7352 107350 7404
rect 107764 7392 107792 7432
rect 107838 7420 107844 7472
rect 107896 7420 107902 7472
rect 117608 7469 117636 7500
rect 123202 7488 123208 7540
rect 123260 7528 123266 7540
rect 123260 7500 215294 7528
rect 123260 7488 123266 7500
rect 117593 7463 117651 7469
rect 108040 7432 113174 7460
rect 108040 7392 108068 7432
rect 107764 7364 108068 7392
rect 110138 7352 110144 7404
rect 110196 7392 110202 7404
rect 110785 7395 110843 7401
rect 110785 7392 110797 7395
rect 110196 7364 110797 7392
rect 110196 7352 110202 7364
rect 110785 7361 110797 7364
rect 110831 7361 110843 7395
rect 110785 7355 110843 7361
rect 59630 7284 59636 7336
rect 59688 7284 59694 7336
rect 61749 7327 61807 7333
rect 61749 7293 61761 7327
rect 61795 7293 61807 7327
rect 61749 7287 61807 7293
rect 58805 7259 58863 7265
rect 58805 7256 58817 7259
rect 29512 7228 58817 7256
rect 29512 7216 29518 7228
rect 58805 7225 58817 7228
rect 58851 7225 58863 7259
rect 61764 7256 61792 7287
rect 63770 7284 63776 7336
rect 63828 7284 63834 7336
rect 65058 7284 65064 7336
rect 65116 7284 65122 7336
rect 66714 7284 66720 7336
rect 66772 7284 66778 7336
rect 79318 7284 79324 7336
rect 79376 7284 79382 7336
rect 80606 7284 80612 7336
rect 80664 7284 80670 7336
rect 111334 7284 111340 7336
rect 111392 7284 111398 7336
rect 113146 7324 113174 7432
rect 117593 7429 117605 7463
rect 117639 7429 117651 7463
rect 117593 7423 117651 7429
rect 120629 7463 120687 7469
rect 120629 7429 120641 7463
rect 120675 7460 120687 7463
rect 213365 7463 213423 7469
rect 213365 7460 213377 7463
rect 120675 7432 213377 7460
rect 120675 7429 120687 7432
rect 120629 7423 120687 7429
rect 213365 7429 213377 7432
rect 213411 7429 213423 7463
rect 215266 7460 215294 7500
rect 216033 7463 216091 7469
rect 216033 7460 216045 7463
rect 215266 7432 216045 7460
rect 213365 7423 213423 7429
rect 216033 7429 216045 7432
rect 216079 7429 216091 7463
rect 216033 7423 216091 7429
rect 117869 7395 117927 7401
rect 117869 7361 117881 7395
rect 117915 7392 117927 7395
rect 117958 7392 117964 7404
rect 117915 7364 117964 7392
rect 117915 7361 117927 7364
rect 117869 7355 117927 7361
rect 117958 7352 117964 7364
rect 118016 7352 118022 7404
rect 119249 7395 119307 7401
rect 119249 7361 119261 7395
rect 119295 7392 119307 7395
rect 119338 7392 119344 7404
rect 119295 7364 119344 7392
rect 119295 7361 119307 7364
rect 119249 7355 119307 7361
rect 119338 7352 119344 7364
rect 119396 7352 119402 7404
rect 120077 7395 120135 7401
rect 120077 7361 120089 7395
rect 120123 7361 120135 7395
rect 120077 7355 120135 7361
rect 118697 7327 118755 7333
rect 118697 7324 118709 7327
rect 113146 7296 118709 7324
rect 118697 7293 118709 7296
rect 118743 7293 118755 7327
rect 118697 7287 118755 7293
rect 118970 7284 118976 7336
rect 119028 7324 119034 7336
rect 120092 7324 120120 7355
rect 121454 7352 121460 7404
rect 121512 7352 121518 7404
rect 121822 7352 121828 7404
rect 121880 7352 121886 7404
rect 122834 7352 122840 7404
rect 122892 7352 122898 7404
rect 123202 7352 123208 7404
rect 123260 7352 123266 7404
rect 123846 7352 123852 7404
rect 123904 7352 123910 7404
rect 125318 7352 125324 7404
rect 125376 7392 125382 7404
rect 125965 7395 126023 7401
rect 125965 7392 125977 7395
rect 125376 7364 125977 7392
rect 125376 7352 125382 7364
rect 125965 7361 125977 7364
rect 126011 7361 126023 7395
rect 125965 7355 126023 7361
rect 151170 7352 151176 7404
rect 151228 7352 151234 7404
rect 152734 7352 152740 7404
rect 152792 7392 152798 7404
rect 153473 7395 153531 7401
rect 153473 7392 153485 7395
rect 152792 7364 153485 7392
rect 152792 7352 152798 7364
rect 153473 7361 153485 7364
rect 153519 7361 153531 7395
rect 154761 7395 154819 7401
rect 154761 7392 154773 7395
rect 153473 7355 153531 7361
rect 154592 7364 154773 7392
rect 119028 7296 120120 7324
rect 124401 7327 124459 7333
rect 119028 7284 119034 7296
rect 124401 7293 124413 7327
rect 124447 7324 124459 7327
rect 125502 7324 125508 7336
rect 124447 7296 125508 7324
rect 124447 7293 124459 7296
rect 124401 7287 124459 7293
rect 125502 7284 125508 7296
rect 125560 7284 125566 7336
rect 126514 7284 126520 7336
rect 126572 7284 126578 7336
rect 151722 7284 151728 7336
rect 151780 7284 151786 7336
rect 154025 7327 154083 7333
rect 154025 7293 154037 7327
rect 154071 7324 154083 7327
rect 154482 7324 154488 7336
rect 154071 7296 154488 7324
rect 154071 7293 154083 7296
rect 154025 7287 154083 7293
rect 154482 7284 154488 7296
rect 154540 7284 154546 7336
rect 154592 7268 154620 7364
rect 154761 7361 154773 7364
rect 154807 7361 154819 7395
rect 154761 7355 154819 7361
rect 166442 7352 166448 7404
rect 166500 7352 166506 7404
rect 168190 7352 168196 7404
rect 168248 7392 168254 7404
rect 168929 7395 168987 7401
rect 168929 7392 168941 7395
rect 168248 7364 168941 7392
rect 168248 7352 168254 7364
rect 168929 7361 168941 7364
rect 168975 7361 168987 7395
rect 168929 7355 168987 7361
rect 170122 7352 170128 7404
rect 170180 7352 170186 7404
rect 197906 7352 197912 7404
rect 197964 7392 197970 7404
rect 198553 7395 198611 7401
rect 198553 7392 198565 7395
rect 197964 7364 198565 7392
rect 197964 7352 197970 7364
rect 198553 7361 198565 7364
rect 198599 7361 198611 7395
rect 198553 7355 198611 7361
rect 200114 7352 200120 7404
rect 200172 7392 200178 7404
rect 200761 7395 200819 7401
rect 200761 7392 200773 7395
rect 200172 7364 200773 7392
rect 200172 7352 200178 7364
rect 200761 7361 200773 7364
rect 200807 7361 200819 7395
rect 213380 7392 213408 7423
rect 214009 7395 214067 7401
rect 214009 7392 214021 7395
rect 213380 7364 214021 7392
rect 200761 7355 200819 7361
rect 214009 7361 214021 7364
rect 214055 7361 214067 7395
rect 214009 7355 214067 7361
rect 217229 7395 217287 7401
rect 217229 7361 217241 7395
rect 217275 7392 217287 7395
rect 217870 7392 217876 7404
rect 217275 7364 217876 7392
rect 217275 7361 217287 7364
rect 217229 7355 217287 7361
rect 217870 7352 217876 7364
rect 217928 7352 217934 7404
rect 219713 7395 219771 7401
rect 219713 7361 219725 7395
rect 219759 7392 219771 7395
rect 220446 7392 220452 7404
rect 219759 7364 220452 7392
rect 219759 7361 219771 7364
rect 219713 7355 219771 7361
rect 220446 7352 220452 7364
rect 220504 7352 220510 7404
rect 244366 7352 244372 7404
rect 244424 7392 244430 7404
rect 244921 7395 244979 7401
rect 244921 7392 244933 7395
rect 244424 7364 244933 7392
rect 244424 7352 244430 7364
rect 244921 7361 244933 7364
rect 244967 7361 244979 7395
rect 260377 7395 260435 7401
rect 260377 7392 260389 7395
rect 244921 7355 244979 7361
rect 259748 7364 260389 7392
rect 155313 7327 155371 7333
rect 155313 7293 155325 7327
rect 155359 7324 155371 7327
rect 157334 7324 157340 7336
rect 155359 7296 157340 7324
rect 155359 7293 155371 7296
rect 155313 7287 155371 7293
rect 157334 7284 157340 7296
rect 157392 7284 157398 7336
rect 166997 7327 167055 7333
rect 166997 7293 167009 7327
rect 167043 7293 167055 7327
rect 166997 7287 167055 7293
rect 154574 7256 154580 7268
rect 61764 7228 154580 7256
rect 58805 7219 58863 7225
rect 154574 7216 154580 7228
rect 154632 7216 154638 7268
rect 167012 7256 167040 7287
rect 169478 7284 169484 7336
rect 169536 7284 169542 7336
rect 170674 7284 170680 7336
rect 170732 7284 170738 7336
rect 199102 7284 199108 7336
rect 199160 7284 199166 7336
rect 201310 7284 201316 7336
rect 201368 7284 201374 7336
rect 214558 7284 214564 7336
rect 214616 7284 214622 7336
rect 214742 7284 214748 7336
rect 214800 7324 214806 7336
rect 218517 7327 218575 7333
rect 218517 7324 218529 7327
rect 214800 7296 218529 7324
rect 214800 7284 214806 7296
rect 218517 7293 218529 7296
rect 218563 7293 218575 7327
rect 218517 7287 218575 7293
rect 245470 7284 245476 7336
rect 245528 7284 245534 7336
rect 259748 7265 259776 7364
rect 260377 7361 260389 7364
rect 260423 7361 260435 7395
rect 260377 7355 260435 7361
rect 260742 7284 260748 7336
rect 260800 7284 260806 7336
rect 259733 7259 259791 7265
rect 259733 7256 259745 7259
rect 167012 7228 259745 7256
rect 259733 7225 259745 7228
rect 259779 7225 259791 7259
rect 259733 7219 259791 7225
rect 152734 7148 152740 7200
rect 152792 7148 152798 7200
rect 217870 7148 217876 7200
rect 217928 7148 217934 7200
rect 220446 7148 220452 7200
rect 220504 7148 220510 7200
rect 1104 7098 648876 7120
rect 1104 7046 81921 7098
rect 81973 7046 81985 7098
rect 82037 7046 82049 7098
rect 82101 7046 82113 7098
rect 82165 7046 82177 7098
rect 82229 7046 243864 7098
rect 243916 7046 243928 7098
rect 243980 7046 243992 7098
rect 244044 7046 244056 7098
rect 244108 7046 244120 7098
rect 244172 7046 405807 7098
rect 405859 7046 405871 7098
rect 405923 7046 405935 7098
rect 405987 7046 405999 7098
rect 406051 7046 406063 7098
rect 406115 7046 567750 7098
rect 567802 7046 567814 7098
rect 567866 7046 567878 7098
rect 567930 7046 567942 7098
rect 567994 7046 568006 7098
rect 568058 7046 648876 7098
rect 1104 7024 648876 7046
rect 24578 6944 24584 6996
rect 24636 6984 24642 6996
rect 24636 6956 35894 6984
rect 24636 6944 24642 6956
rect 35161 6919 35219 6925
rect 35161 6885 35173 6919
rect 35207 6916 35219 6919
rect 35250 6916 35256 6928
rect 35207 6888 35256 6916
rect 35207 6885 35219 6888
rect 35161 6879 35219 6885
rect 35250 6876 35256 6888
rect 35308 6876 35314 6928
rect 35866 6916 35894 6956
rect 59630 6944 59636 6996
rect 59688 6984 59694 6996
rect 152734 6984 152740 6996
rect 59688 6956 152740 6984
rect 59688 6944 59694 6956
rect 152734 6944 152740 6956
rect 152792 6944 152798 6996
rect 166261 6987 166319 6993
rect 154408 6956 157334 6984
rect 64601 6919 64659 6925
rect 64601 6916 64613 6919
rect 35866 6888 64613 6916
rect 64601 6885 64613 6888
rect 64647 6916 64659 6919
rect 64782 6916 64788 6928
rect 64647 6888 64788 6916
rect 64647 6885 64659 6888
rect 64601 6879 64659 6885
rect 64782 6876 64788 6888
rect 64840 6876 64846 6928
rect 107105 6919 107163 6925
rect 107105 6885 107117 6919
rect 107151 6916 107163 6919
rect 107286 6916 107292 6928
rect 107151 6888 107292 6916
rect 107151 6885 107163 6888
rect 107105 6879 107163 6885
rect 107286 6876 107292 6888
rect 107344 6876 107350 6928
rect 118970 6876 118976 6928
rect 119028 6876 119034 6928
rect 122929 6919 122987 6925
rect 122929 6885 122941 6919
rect 122975 6916 122987 6919
rect 123202 6916 123208 6928
rect 122975 6888 123208 6916
rect 122975 6885 122987 6888
rect 122929 6879 122987 6885
rect 123202 6876 123208 6888
rect 123260 6876 123266 6928
rect 150989 6919 151047 6925
rect 150989 6885 151001 6919
rect 151035 6916 151047 6919
rect 151170 6916 151176 6928
rect 151035 6888 151176 6916
rect 151035 6885 151047 6888
rect 150989 6879 151047 6885
rect 151170 6876 151176 6888
rect 151228 6876 151234 6928
rect 151722 6876 151728 6928
rect 151780 6916 151786 6928
rect 154408 6916 154436 6956
rect 151780 6888 154436 6916
rect 151780 6876 151786 6888
rect 154574 6876 154580 6928
rect 154632 6876 154638 6928
rect 157306 6916 157334 6956
rect 166261 6953 166273 6987
rect 166307 6984 166319 6987
rect 166442 6984 166448 6996
rect 166307 6956 166448 6984
rect 166307 6953 166319 6956
rect 166261 6947 166319 6953
rect 166442 6944 166448 6956
rect 166500 6944 166506 6996
rect 169941 6987 169999 6993
rect 169941 6953 169953 6987
rect 169987 6984 169999 6987
rect 170122 6984 170128 6996
rect 169987 6956 170128 6984
rect 169987 6953 169999 6956
rect 169941 6947 169999 6953
rect 170122 6944 170128 6956
rect 170180 6944 170186 6996
rect 170214 6944 170220 6996
rect 170272 6984 170278 6996
rect 172330 6984 172336 6996
rect 170272 6956 172336 6984
rect 170272 6944 170278 6956
rect 172330 6944 172336 6956
rect 172388 6944 172394 6996
rect 215294 6944 215300 6996
rect 215352 6984 215358 6996
rect 218790 6984 218796 6996
rect 215352 6956 218796 6984
rect 215352 6944 215358 6956
rect 218790 6944 218796 6956
rect 218848 6944 218854 6996
rect 215846 6916 215852 6928
rect 157306 6888 215852 6916
rect 215846 6876 215852 6888
rect 215904 6876 215910 6928
rect 216030 6876 216036 6928
rect 216088 6916 216094 6928
rect 244366 6916 244372 6928
rect 216088 6888 244372 6916
rect 216088 6876 216094 6888
rect 244366 6876 244372 6888
rect 244424 6876 244430 6928
rect 17862 6808 17868 6860
rect 17920 6848 17926 6860
rect 19702 6848 19708 6860
rect 17920 6820 19708 6848
rect 17920 6808 17926 6820
rect 19702 6808 19708 6820
rect 19760 6808 19766 6860
rect 26694 6808 26700 6860
rect 26752 6848 26758 6860
rect 119617 6851 119675 6857
rect 119617 6848 119629 6851
rect 26752 6820 119629 6848
rect 26752 6808 26758 6820
rect 119617 6817 119629 6820
rect 119663 6817 119675 6851
rect 123481 6851 123539 6857
rect 123481 6848 123493 6851
rect 119617 6811 119675 6817
rect 120092 6820 123493 6848
rect 18046 6740 18052 6792
rect 18104 6780 18110 6792
rect 20162 6780 20168 6792
rect 18104 6752 20168 6780
rect 18104 6740 18110 6752
rect 20162 6740 20168 6752
rect 20220 6740 20226 6792
rect 63034 6740 63040 6792
rect 63092 6780 63098 6792
rect 63313 6783 63371 6789
rect 63313 6780 63325 6783
rect 63092 6752 63325 6780
rect 63092 6740 63098 6752
rect 63313 6749 63325 6752
rect 63359 6749 63371 6783
rect 63313 6743 63371 6749
rect 79594 6740 79600 6792
rect 79652 6780 79658 6792
rect 79781 6783 79839 6789
rect 79781 6780 79793 6783
rect 79652 6752 79793 6780
rect 79652 6740 79658 6752
rect 79781 6749 79793 6752
rect 79827 6749 79839 6783
rect 79781 6743 79839 6749
rect 81526 6740 81532 6792
rect 81584 6740 81590 6792
rect 81636 6752 84194 6780
rect 30006 6672 30012 6724
rect 30064 6712 30070 6724
rect 81636 6712 81664 6752
rect 30064 6684 81664 6712
rect 82081 6715 82139 6721
rect 30064 6672 30070 6684
rect 82081 6681 82093 6715
rect 82127 6712 82139 6715
rect 82446 6712 82452 6724
rect 82127 6684 82452 6712
rect 82127 6681 82139 6684
rect 82081 6675 82139 6681
rect 82446 6672 82452 6684
rect 82504 6672 82510 6724
rect 84166 6712 84194 6752
rect 108482 6740 108488 6792
rect 108540 6780 108546 6792
rect 109129 6783 109187 6789
rect 109129 6780 109141 6783
rect 108540 6752 109141 6780
rect 108540 6740 108546 6752
rect 109129 6749 109141 6752
rect 109175 6749 109187 6783
rect 116673 6783 116731 6789
rect 109129 6743 109187 6749
rect 109236 6752 116256 6780
rect 109236 6712 109264 6752
rect 84166 6684 109264 6712
rect 109681 6715 109739 6721
rect 109681 6681 109693 6715
rect 109727 6712 109739 6715
rect 109727 6684 113174 6712
rect 109727 6681 109739 6684
rect 109681 6675 109739 6681
rect 113146 6644 113174 6684
rect 116118 6672 116124 6724
rect 116176 6672 116182 6724
rect 116228 6712 116256 6752
rect 116673 6749 116685 6783
rect 116719 6780 116731 6783
rect 117038 6780 117044 6792
rect 116719 6752 117044 6780
rect 116719 6749 116731 6752
rect 116673 6743 116731 6749
rect 117038 6740 117044 6752
rect 117096 6740 117102 6792
rect 120092 6780 120120 6820
rect 123481 6817 123493 6820
rect 123527 6817 123539 6851
rect 170214 6848 170220 6860
rect 123481 6811 123539 6817
rect 142126 6820 162256 6848
rect 117148 6752 120120 6780
rect 120169 6783 120227 6789
rect 117148 6712 117176 6752
rect 120169 6749 120181 6783
rect 120215 6780 120227 6783
rect 120442 6780 120448 6792
rect 120215 6752 120448 6780
rect 120215 6749 120227 6752
rect 120169 6743 120227 6749
rect 120442 6740 120448 6752
rect 120500 6740 120506 6792
rect 121365 6783 121423 6789
rect 121365 6749 121377 6783
rect 121411 6780 121423 6783
rect 121454 6780 121460 6792
rect 121411 6752 121460 6780
rect 121411 6749 121423 6752
rect 121365 6743 121423 6749
rect 121454 6740 121460 6752
rect 121512 6740 121518 6792
rect 124030 6740 124036 6792
rect 124088 6740 124094 6792
rect 125229 6783 125287 6789
rect 125229 6749 125241 6783
rect 125275 6780 125287 6783
rect 125873 6783 125931 6789
rect 125873 6780 125885 6783
rect 125275 6752 125885 6780
rect 125275 6749 125287 6752
rect 125229 6743 125287 6749
rect 125873 6749 125885 6752
rect 125919 6780 125931 6783
rect 125919 6752 132494 6780
rect 125919 6749 125931 6752
rect 125873 6743 125931 6749
rect 116228 6684 117176 6712
rect 117240 6684 118096 6712
rect 117240 6644 117268 6684
rect 113146 6616 117268 6644
rect 117406 6604 117412 6656
rect 117464 6604 117470 6656
rect 117958 6604 117964 6656
rect 118016 6604 118022 6656
rect 118068 6644 118096 6684
rect 118666 6684 119108 6712
rect 118666 6644 118694 6684
rect 118068 6616 118694 6644
rect 119080 6644 119108 6684
rect 120810 6672 120816 6724
rect 120868 6672 120874 6724
rect 122668 6684 122972 6712
rect 122668 6644 122696 6684
rect 119080 6616 122696 6644
rect 122944 6644 122972 6684
rect 124674 6672 124680 6724
rect 124732 6672 124738 6724
rect 132466 6712 132494 6752
rect 142126 6712 142154 6820
rect 155770 6740 155776 6792
rect 155828 6780 155834 6792
rect 156417 6783 156475 6789
rect 156417 6780 156429 6783
rect 155828 6752 156429 6780
rect 155828 6740 155834 6752
rect 156417 6749 156429 6752
rect 156463 6749 156475 6783
rect 156417 6743 156475 6749
rect 132466 6684 142154 6712
rect 154592 6684 155908 6712
rect 154592 6644 154620 6684
rect 122944 6616 154620 6644
rect 155770 6604 155776 6656
rect 155828 6604 155834 6656
rect 155880 6644 155908 6684
rect 156966 6672 156972 6724
rect 157024 6672 157030 6724
rect 162228 6712 162256 6820
rect 164206 6820 170220 6848
rect 164206 6712 164234 6820
rect 170214 6808 170220 6820
rect 170272 6808 170278 6860
rect 170674 6808 170680 6860
rect 170732 6848 170738 6860
rect 215754 6848 215760 6860
rect 170732 6820 215760 6848
rect 170732 6808 170738 6820
rect 215754 6808 215760 6820
rect 215812 6808 215818 6860
rect 216214 6808 216220 6860
rect 216272 6848 216278 6860
rect 262950 6848 262956 6860
rect 216272 6820 262956 6848
rect 216272 6808 216278 6820
rect 262950 6808 262956 6820
rect 263008 6808 263014 6860
rect 171042 6740 171048 6792
rect 171100 6780 171106 6792
rect 171643 6783 171701 6789
rect 171643 6780 171655 6783
rect 171100 6752 171655 6780
rect 171100 6740 171106 6752
rect 171643 6749 171655 6752
rect 171689 6749 171701 6783
rect 171643 6743 171701 6749
rect 173066 6740 173072 6792
rect 173124 6780 173130 6792
rect 215294 6780 215300 6792
rect 173124 6752 215300 6780
rect 173124 6740 173130 6752
rect 215294 6740 215300 6752
rect 215352 6740 215358 6792
rect 215987 6783 216045 6789
rect 215987 6780 215999 6783
rect 215496 6752 215999 6780
rect 162228 6684 164234 6712
rect 169036 6684 171640 6712
rect 169036 6644 169064 6684
rect 155880 6616 169064 6644
rect 171042 6604 171048 6656
rect 171100 6604 171106 6656
rect 171612 6644 171640 6684
rect 172238 6672 172244 6724
rect 172296 6672 172302 6724
rect 172330 6672 172336 6724
rect 172388 6712 172394 6724
rect 214742 6712 214748 6724
rect 172388 6684 214748 6712
rect 172388 6672 172394 6684
rect 214742 6672 214748 6684
rect 214800 6672 214806 6724
rect 190546 6644 190552 6656
rect 171612 6616 190552 6644
rect 190546 6604 190552 6616
rect 190604 6604 190610 6656
rect 190638 6604 190644 6656
rect 190696 6644 190702 6656
rect 213270 6644 213276 6656
rect 190696 6616 213276 6644
rect 190696 6604 190702 6616
rect 213270 6604 213276 6616
rect 213328 6604 213334 6656
rect 213362 6604 213368 6656
rect 213420 6644 213426 6656
rect 215496 6653 215524 6752
rect 215987 6749 215999 6752
rect 216033 6749 216045 6783
rect 215987 6743 216045 6749
rect 218701 6783 218759 6789
rect 218701 6749 218713 6783
rect 218747 6749 218759 6783
rect 218701 6743 218759 6749
rect 216582 6672 216588 6724
rect 216640 6672 216646 6724
rect 217502 6672 217508 6724
rect 217560 6672 217566 6724
rect 215481 6647 215539 6653
rect 215481 6644 215493 6647
rect 213420 6616 215493 6644
rect 213420 6604 213426 6616
rect 215481 6613 215493 6616
rect 215527 6613 215539 6647
rect 218716 6644 218744 6743
rect 218790 6740 218796 6792
rect 218848 6780 218854 6792
rect 218848 6752 246712 6780
rect 218848 6740 218854 6752
rect 246684 6712 246712 6752
rect 246758 6740 246764 6792
rect 246816 6740 246822 6792
rect 261754 6780 261760 6792
rect 246868 6752 261760 6780
rect 246868 6712 246896 6752
rect 261754 6740 261760 6752
rect 261812 6780 261818 6792
rect 262033 6783 262091 6789
rect 262033 6780 262045 6783
rect 261812 6752 262045 6780
rect 261812 6740 261818 6752
rect 262033 6749 262045 6752
rect 262079 6749 262091 6783
rect 262033 6743 262091 6749
rect 234586 6684 246620 6712
rect 246684 6684 246896 6712
rect 219253 6647 219311 6653
rect 219253 6644 219265 6647
rect 218716 6616 219265 6644
rect 215481 6607 215539 6613
rect 219253 6613 219265 6616
rect 219299 6644 219311 6647
rect 234586 6644 234614 6684
rect 219299 6616 234614 6644
rect 219299 6613 219311 6616
rect 219253 6607 219311 6613
rect 246114 6604 246120 6656
rect 246172 6604 246178 6656
rect 246592 6644 246620 6684
rect 247310 6672 247316 6724
rect 247368 6672 247374 6724
rect 262582 6672 262588 6724
rect 262640 6672 262646 6724
rect 310882 6644 310888 6656
rect 246592 6616 310888 6644
rect 310882 6604 310888 6616
rect 310940 6604 310946 6656
rect 1104 6554 648876 6576
rect 1104 6502 82581 6554
rect 82633 6502 82645 6554
rect 82697 6502 82709 6554
rect 82761 6502 82773 6554
rect 82825 6502 82837 6554
rect 82889 6502 244524 6554
rect 244576 6502 244588 6554
rect 244640 6502 244652 6554
rect 244704 6502 244716 6554
rect 244768 6502 244780 6554
rect 244832 6502 406467 6554
rect 406519 6502 406531 6554
rect 406583 6502 406595 6554
rect 406647 6502 406659 6554
rect 406711 6502 406723 6554
rect 406775 6502 568410 6554
rect 568462 6502 568474 6554
rect 568526 6502 568538 6554
rect 568590 6502 568602 6554
rect 568654 6502 568666 6554
rect 568718 6502 648876 6554
rect 1104 6480 648876 6502
rect 63770 6400 63776 6452
rect 63828 6440 63834 6452
rect 155770 6440 155776 6452
rect 63828 6412 155776 6440
rect 63828 6400 63834 6412
rect 155770 6400 155776 6412
rect 155828 6400 155834 6452
rect 157334 6400 157340 6452
rect 157392 6440 157398 6452
rect 167178 6440 167184 6452
rect 157392 6412 167184 6440
rect 157392 6400 157398 6412
rect 167178 6400 167184 6412
rect 167236 6400 167242 6452
rect 169478 6400 169484 6452
rect 169536 6440 169542 6452
rect 173066 6440 173072 6452
rect 169536 6412 173072 6440
rect 169536 6400 169542 6412
rect 173066 6400 173072 6412
rect 173124 6400 173130 6452
rect 173158 6400 173164 6452
rect 173216 6440 173222 6452
rect 190638 6440 190644 6452
rect 173216 6412 190644 6440
rect 173216 6400 173222 6412
rect 190638 6400 190644 6412
rect 190696 6400 190702 6452
rect 190730 6400 190736 6452
rect 190788 6440 190794 6452
rect 200574 6440 200580 6452
rect 190788 6412 200580 6440
rect 190788 6400 190794 6412
rect 200574 6400 200580 6412
rect 200632 6400 200638 6452
rect 200684 6412 209774 6440
rect 23750 6332 23756 6384
rect 23808 6372 23814 6384
rect 111153 6375 111211 6381
rect 111153 6372 111165 6375
rect 23808 6344 111165 6372
rect 23808 6332 23814 6344
rect 111153 6341 111165 6344
rect 111199 6341 111211 6375
rect 111153 6335 111211 6341
rect 123757 6375 123815 6381
rect 123757 6341 123769 6375
rect 123803 6372 123815 6375
rect 123846 6372 123852 6384
rect 123803 6344 123852 6372
rect 123803 6341 123815 6344
rect 123757 6335 123815 6341
rect 27522 6264 27528 6316
rect 27580 6304 27586 6316
rect 111168 6304 111196 6335
rect 123846 6332 123852 6344
rect 123904 6332 123910 6384
rect 124030 6332 124036 6384
rect 124088 6372 124094 6384
rect 124309 6375 124367 6381
rect 124309 6372 124321 6375
rect 124088 6344 124321 6372
rect 124088 6332 124094 6344
rect 124309 6341 124321 6344
rect 124355 6372 124367 6375
rect 200684 6372 200712 6412
rect 209746 6372 209774 6412
rect 214558 6400 214564 6452
rect 214616 6440 214622 6452
rect 307481 6443 307539 6449
rect 307481 6440 307493 6443
rect 214616 6412 307493 6440
rect 214616 6400 214622 6412
rect 307481 6409 307493 6412
rect 307527 6409 307539 6443
rect 307481 6403 307539 6409
rect 217502 6372 217508 6384
rect 124355 6344 200712 6372
rect 200776 6344 205634 6372
rect 209746 6344 217508 6372
rect 124355 6341 124367 6344
rect 124309 6335 124367 6341
rect 111797 6307 111855 6313
rect 111797 6304 111809 6307
rect 27580 6276 103514 6304
rect 111168 6276 111809 6304
rect 27580 6264 27586 6276
rect 103486 6236 103514 6276
rect 111797 6273 111809 6276
rect 111843 6273 111855 6307
rect 120810 6304 120816 6316
rect 111797 6267 111855 6273
rect 111904 6276 120816 6304
rect 111904 6236 111932 6276
rect 120810 6264 120816 6276
rect 120868 6264 120874 6316
rect 122558 6264 122564 6316
rect 122616 6264 122622 6316
rect 123021 6307 123079 6313
rect 123021 6273 123033 6307
rect 123067 6304 123079 6307
rect 123067 6276 126744 6304
rect 123067 6273 123079 6276
rect 123021 6267 123079 6273
rect 103486 6208 111932 6236
rect 112346 6196 112352 6248
rect 112404 6196 112410 6248
rect 126716 6236 126744 6276
rect 126882 6264 126888 6316
rect 126940 6304 126946 6316
rect 126977 6307 127035 6313
rect 126977 6304 126989 6307
rect 126940 6276 126989 6304
rect 126940 6264 126946 6276
rect 126977 6273 126989 6276
rect 127023 6273 127035 6307
rect 200776 6304 200804 6344
rect 202417 6307 202475 6313
rect 202417 6304 202429 6307
rect 126977 6267 127035 6273
rect 127176 6276 200804 6304
rect 201696 6276 202429 6304
rect 127176 6236 127204 6276
rect 126716 6208 127204 6236
rect 127526 6196 127532 6248
rect 127584 6196 127590 6248
rect 127618 6196 127624 6248
rect 127676 6236 127682 6248
rect 127676 6208 198780 6236
rect 127676 6196 127682 6208
rect 20622 6128 20628 6180
rect 20680 6168 20686 6180
rect 32490 6168 32496 6180
rect 20680 6140 32496 6168
rect 20680 6128 20686 6140
rect 32490 6128 32496 6140
rect 32548 6128 32554 6180
rect 35526 6128 35532 6180
rect 35584 6168 35590 6180
rect 126333 6171 126391 6177
rect 126333 6168 126345 6171
rect 35584 6140 126345 6168
rect 35584 6128 35590 6140
rect 126333 6137 126345 6140
rect 126379 6168 126391 6171
rect 126882 6168 126888 6180
rect 126379 6140 126888 6168
rect 126379 6137 126391 6140
rect 126333 6131 126391 6137
rect 126882 6128 126888 6140
rect 126940 6128 126946 6180
rect 126974 6128 126980 6180
rect 127032 6168 127038 6180
rect 171042 6168 171048 6180
rect 127032 6140 171048 6168
rect 127032 6128 127038 6140
rect 171042 6128 171048 6140
rect 171100 6128 171106 6180
rect 198752 6168 198780 6208
rect 200574 6196 200580 6248
rect 200632 6236 200638 6248
rect 201696 6245 201724 6276
rect 202417 6273 202429 6276
rect 202463 6273 202475 6307
rect 205606 6304 205634 6344
rect 217502 6332 217508 6344
rect 217560 6332 217566 6384
rect 260742 6332 260748 6384
rect 260800 6372 260806 6384
rect 260800 6344 302234 6372
rect 260800 6332 260806 6344
rect 213362 6304 213368 6316
rect 205606 6276 213368 6304
rect 202417 6267 202475 6273
rect 213362 6264 213368 6276
rect 213420 6264 213426 6316
rect 213457 6307 213515 6313
rect 213457 6273 213469 6307
rect 213503 6304 213515 6307
rect 213638 6304 213644 6316
rect 213503 6276 213644 6304
rect 213503 6273 213515 6276
rect 213457 6267 213515 6273
rect 213638 6264 213644 6276
rect 213696 6264 213702 6316
rect 214653 6307 214711 6313
rect 213748 6276 214420 6304
rect 201681 6239 201739 6245
rect 201681 6236 201693 6239
rect 200632 6208 201693 6236
rect 200632 6196 200638 6208
rect 201681 6205 201693 6208
rect 201727 6205 201739 6239
rect 201681 6199 201739 6205
rect 202782 6196 202788 6248
rect 202840 6196 202846 6248
rect 211522 6236 211528 6248
rect 203076 6208 211528 6236
rect 203076 6168 203104 6208
rect 211522 6196 211528 6208
rect 211580 6196 211586 6248
rect 212902 6196 212908 6248
rect 212960 6196 212966 6248
rect 213270 6196 213276 6248
rect 213328 6236 213334 6248
rect 213748 6236 213776 6276
rect 213328 6208 213776 6236
rect 213328 6196 213334 6208
rect 214098 6196 214104 6248
rect 214156 6196 214162 6248
rect 214392 6236 214420 6276
rect 214653 6273 214665 6307
rect 214699 6304 214711 6307
rect 214926 6304 214932 6316
rect 214699 6276 214932 6304
rect 214699 6273 214711 6276
rect 214653 6267 214711 6273
rect 214926 6264 214932 6276
rect 214984 6264 214990 6316
rect 215849 6307 215907 6313
rect 215036 6276 215616 6304
rect 215036 6236 215064 6276
rect 214392 6208 215064 6236
rect 215110 6196 215116 6248
rect 215168 6236 215174 6248
rect 215297 6239 215355 6245
rect 215297 6236 215309 6239
rect 215168 6208 215309 6236
rect 215168 6196 215174 6208
rect 215297 6205 215309 6208
rect 215343 6205 215355 6239
rect 215588 6236 215616 6276
rect 215849 6273 215861 6307
rect 215895 6304 215907 6307
rect 216490 6304 216496 6316
rect 215895 6276 216496 6304
rect 215895 6273 215907 6276
rect 215849 6267 215907 6273
rect 216490 6264 216496 6276
rect 216548 6264 216554 6316
rect 217873 6307 217931 6313
rect 217873 6273 217885 6307
rect 217919 6273 217931 6307
rect 217873 6267 217931 6273
rect 217137 6239 217195 6245
rect 217137 6236 217149 6239
rect 215588 6208 217149 6236
rect 215297 6199 215355 6205
rect 217137 6205 217149 6208
rect 217183 6236 217195 6239
rect 217888 6236 217916 6267
rect 220446 6264 220452 6316
rect 220504 6304 220510 6316
rect 292574 6304 292580 6316
rect 220504 6276 292580 6304
rect 220504 6264 220510 6276
rect 292574 6264 292580 6276
rect 292632 6264 292638 6316
rect 292758 6264 292764 6316
rect 292816 6264 292822 6316
rect 217183 6208 217916 6236
rect 217183 6205 217195 6208
rect 217137 6199 217195 6205
rect 218422 6196 218428 6248
rect 218480 6196 218486 6248
rect 261754 6196 261760 6248
rect 261812 6196 261818 6248
rect 293310 6196 293316 6248
rect 293368 6196 293374 6248
rect 302206 6236 302234 6344
rect 307496 6304 307524 6403
rect 353573 6375 353631 6381
rect 353573 6372 353585 6375
rect 308232 6344 353585 6372
rect 308125 6307 308183 6313
rect 308125 6304 308137 6307
rect 307496 6276 308137 6304
rect 308125 6273 308137 6276
rect 308171 6273 308183 6307
rect 308125 6267 308183 6273
rect 308232 6236 308260 6344
rect 353573 6341 353585 6344
rect 353619 6341 353631 6375
rect 353573 6335 353631 6341
rect 310882 6264 310888 6316
rect 310940 6264 310946 6316
rect 311713 6307 311771 6313
rect 311713 6273 311725 6307
rect 311759 6304 311771 6307
rect 311894 6304 311900 6316
rect 311759 6276 311900 6304
rect 311759 6273 311771 6276
rect 311713 6267 311771 6273
rect 311894 6264 311900 6276
rect 311952 6264 311958 6316
rect 313185 6307 313243 6313
rect 313185 6273 313197 6307
rect 313231 6304 313243 6307
rect 313734 6304 313740 6316
rect 313231 6276 313740 6304
rect 313231 6273 313243 6276
rect 313185 6267 313243 6273
rect 313734 6264 313740 6276
rect 313792 6264 313798 6316
rect 338853 6307 338911 6313
rect 338853 6304 338865 6307
rect 338224 6276 338865 6304
rect 302206 6208 308260 6236
rect 308674 6196 308680 6248
rect 308732 6196 308738 6248
rect 312357 6239 312415 6245
rect 312357 6236 312369 6239
rect 311866 6208 312369 6236
rect 180766 6140 195974 6168
rect 198752 6140 203104 6168
rect 23198 6060 23204 6112
rect 23256 6100 23262 6112
rect 81253 6103 81311 6109
rect 81253 6100 81265 6103
rect 23256 6072 81265 6100
rect 23256 6060 23262 6072
rect 81253 6069 81265 6072
rect 81299 6100 81311 6103
rect 81526 6100 81532 6112
rect 81299 6072 81532 6100
rect 81299 6069 81311 6072
rect 81253 6063 81311 6069
rect 81526 6060 81532 6072
rect 81584 6060 81590 6112
rect 119338 6060 119344 6112
rect 119396 6060 119402 6112
rect 120442 6060 120448 6112
rect 120500 6060 120506 6112
rect 121454 6060 121460 6112
rect 121512 6060 121518 6112
rect 121822 6060 121828 6112
rect 121880 6100 121886 6112
rect 122009 6103 122067 6109
rect 122009 6100 122021 6103
rect 121880 6072 122021 6100
rect 121880 6060 121886 6072
rect 122009 6069 122021 6072
rect 122055 6100 122067 6103
rect 180766 6100 180794 6140
rect 122055 6072 180794 6100
rect 195946 6100 195974 6140
rect 203150 6128 203156 6180
rect 203208 6168 203214 6180
rect 292117 6171 292175 6177
rect 292117 6168 292129 6171
rect 203208 6140 215064 6168
rect 203208 6128 203214 6140
rect 214926 6100 214932 6112
rect 195946 6072 214932 6100
rect 122055 6069 122067 6072
rect 122009 6063 122067 6069
rect 214926 6060 214932 6072
rect 214984 6060 214990 6112
rect 215036 6100 215064 6140
rect 215266 6140 292129 6168
rect 215266 6100 215294 6140
rect 292117 6137 292129 6140
rect 292163 6168 292175 6171
rect 292163 6140 292574 6168
rect 292163 6137 292175 6140
rect 292117 6131 292175 6137
rect 215036 6072 215294 6100
rect 216490 6060 216496 6112
rect 216548 6060 216554 6112
rect 292546 6100 292574 6140
rect 292666 6128 292672 6180
rect 292724 6168 292730 6180
rect 311866 6168 311894 6208
rect 312357 6205 312369 6208
rect 312403 6205 312415 6239
rect 312357 6199 312415 6205
rect 292724 6140 311894 6168
rect 292724 6128 292730 6140
rect 338224 6112 338252 6276
rect 338853 6273 338865 6276
rect 338899 6273 338911 6307
rect 353588 6304 353616 6335
rect 354217 6307 354275 6313
rect 354217 6304 354229 6307
rect 353588 6276 354229 6304
rect 338853 6267 338911 6273
rect 354217 6273 354229 6276
rect 354263 6273 354275 6307
rect 354217 6267 354275 6273
rect 339402 6196 339408 6248
rect 339460 6196 339466 6248
rect 354582 6196 354588 6248
rect 354640 6196 354646 6248
rect 292758 6100 292764 6112
rect 292546 6072 292764 6100
rect 292758 6060 292764 6072
rect 292816 6060 292822 6112
rect 313734 6060 313740 6112
rect 313792 6060 313798 6112
rect 338206 6060 338212 6112
rect 338264 6060 338270 6112
rect 1104 6010 648876 6032
rect 1104 5958 81921 6010
rect 81973 5958 81985 6010
rect 82037 5958 82049 6010
rect 82101 5958 82113 6010
rect 82165 5958 82177 6010
rect 82229 5958 243864 6010
rect 243916 5958 243928 6010
rect 243980 5958 243992 6010
rect 244044 5958 244056 6010
rect 244108 5958 244120 6010
rect 244172 5958 405807 6010
rect 405859 5958 405871 6010
rect 405923 5958 405935 6010
rect 405987 5958 405999 6010
rect 406051 5958 406063 6010
rect 406115 5958 567750 6010
rect 567802 5958 567814 6010
rect 567866 5958 567878 6010
rect 567930 5958 567942 6010
rect 567994 5958 568006 6010
rect 568058 5958 648876 6010
rect 1104 5936 648876 5958
rect 24302 5856 24308 5908
rect 24360 5896 24366 5908
rect 116118 5896 116124 5908
rect 24360 5868 116124 5896
rect 24360 5856 24366 5868
rect 116118 5856 116124 5868
rect 116176 5856 116182 5908
rect 120442 5856 120448 5908
rect 120500 5896 120506 5908
rect 212902 5896 212908 5908
rect 120500 5868 212908 5896
rect 120500 5856 120506 5868
rect 212902 5856 212908 5868
rect 212960 5856 212966 5908
rect 245470 5856 245476 5908
rect 245528 5896 245534 5908
rect 338206 5896 338212 5908
rect 245528 5868 338212 5896
rect 245528 5856 245534 5868
rect 338206 5856 338212 5868
rect 338264 5856 338270 5908
rect 121454 5788 121460 5840
rect 121512 5828 121518 5840
rect 214098 5828 214104 5840
rect 121512 5800 214104 5828
rect 121512 5788 121518 5800
rect 214098 5788 214104 5800
rect 214156 5788 214162 5840
rect 217870 5788 217876 5840
rect 217928 5828 217934 5840
rect 217928 5800 302234 5828
rect 217928 5788 217934 5800
rect 80606 5720 80612 5772
rect 80664 5760 80670 5772
rect 172057 5763 172115 5769
rect 172057 5760 172069 5763
rect 80664 5732 172069 5760
rect 80664 5720 80670 5732
rect 172057 5729 172069 5732
rect 172103 5760 172115 5763
rect 172103 5732 172744 5760
rect 172103 5729 172115 5732
rect 172057 5723 172115 5729
rect 65058 5652 65064 5704
rect 65116 5692 65122 5704
rect 115017 5695 115075 5701
rect 65116 5664 114968 5692
rect 65116 5652 65122 5664
rect 23382 5584 23388 5636
rect 23440 5624 23446 5636
rect 114465 5627 114523 5633
rect 114465 5624 114477 5627
rect 23440 5596 114477 5624
rect 23440 5584 23446 5596
rect 114465 5593 114477 5596
rect 114511 5593 114523 5627
rect 114940 5624 114968 5664
rect 115017 5661 115029 5695
rect 115063 5692 115075 5695
rect 115658 5692 115664 5704
rect 115063 5664 115664 5692
rect 115063 5661 115075 5664
rect 115017 5655 115075 5661
rect 115658 5652 115664 5664
rect 115716 5652 115722 5704
rect 172716 5701 172744 5732
rect 199102 5720 199108 5772
rect 199160 5760 199166 5772
rect 203150 5760 203156 5772
rect 199160 5732 203156 5760
rect 199160 5720 199166 5732
rect 203150 5720 203156 5732
rect 203208 5720 203214 5772
rect 293681 5763 293739 5769
rect 293681 5760 293693 5763
rect 205606 5732 293693 5760
rect 156693 5695 156751 5701
rect 156693 5692 156705 5695
rect 118666 5664 156705 5692
rect 118666 5624 118694 5664
rect 156693 5661 156705 5664
rect 156739 5692 156751 5695
rect 157337 5695 157395 5701
rect 157337 5692 157349 5695
rect 156739 5664 157349 5692
rect 156739 5661 156751 5664
rect 156693 5655 156751 5661
rect 157337 5661 157349 5664
rect 157383 5661 157395 5695
rect 157337 5655 157395 5661
rect 172701 5695 172759 5701
rect 172701 5661 172713 5695
rect 172747 5661 172759 5695
rect 172701 5655 172759 5661
rect 201310 5652 201316 5704
rect 201368 5692 201374 5704
rect 205606 5692 205634 5732
rect 293681 5729 293693 5732
rect 293727 5760 293739 5763
rect 302206 5760 302234 5800
rect 310057 5763 310115 5769
rect 310057 5760 310069 5763
rect 293727 5732 294276 5760
rect 302206 5732 310069 5760
rect 293727 5729 293739 5732
rect 293681 5723 293739 5729
rect 201368 5664 205634 5692
rect 201368 5652 201374 5664
rect 211522 5652 211528 5704
rect 211580 5652 211586 5704
rect 212077 5695 212135 5701
rect 212077 5661 212089 5695
rect 212123 5692 212135 5695
rect 212123 5664 212764 5692
rect 212123 5661 212135 5664
rect 212077 5655 212135 5661
rect 114940 5596 118694 5624
rect 114465 5587 114523 5593
rect 119338 5584 119344 5636
rect 119396 5624 119402 5636
rect 127618 5624 127624 5636
rect 119396 5596 127624 5624
rect 119396 5584 119402 5596
rect 127618 5584 127624 5596
rect 127676 5584 127682 5636
rect 157886 5584 157892 5636
rect 157944 5584 157950 5636
rect 166994 5584 167000 5636
rect 167052 5624 167058 5636
rect 173158 5624 173164 5636
rect 167052 5596 173164 5624
rect 167052 5584 167058 5596
rect 173158 5584 173164 5596
rect 173216 5584 173222 5636
rect 173250 5584 173256 5636
rect 173308 5584 173314 5636
rect 212736 5568 212764 5664
rect 247586 5652 247592 5704
rect 247644 5692 247650 5704
rect 248141 5695 248199 5701
rect 248141 5692 248153 5695
rect 247644 5664 248153 5692
rect 247644 5652 247650 5664
rect 248141 5661 248153 5664
rect 248187 5661 248199 5695
rect 248141 5655 248199 5661
rect 262950 5652 262956 5704
rect 263008 5692 263014 5704
rect 294248 5701 294276 5732
rect 310057 5729 310069 5732
rect 310103 5729 310115 5763
rect 310057 5723 310115 5729
rect 263505 5695 263563 5701
rect 263505 5692 263517 5695
rect 263008 5664 263517 5692
rect 263008 5652 263014 5664
rect 263505 5661 263517 5664
rect 263551 5661 263563 5695
rect 263505 5655 263563 5661
rect 294233 5695 294291 5701
rect 294233 5661 294245 5695
rect 294279 5661 294291 5695
rect 294233 5655 294291 5661
rect 310885 5695 310943 5701
rect 310885 5661 310897 5695
rect 310931 5692 310943 5695
rect 311066 5692 311072 5704
rect 310931 5664 311072 5692
rect 310931 5661 310943 5664
rect 310885 5655 310943 5661
rect 311066 5652 311072 5664
rect 311124 5652 311130 5704
rect 248966 5584 248972 5636
rect 249024 5584 249030 5636
rect 264330 5584 264336 5636
rect 264388 5584 264394 5636
rect 295058 5584 295064 5636
rect 295116 5584 295122 5636
rect 28902 5516 28908 5568
rect 28960 5556 28966 5568
rect 122469 5559 122527 5565
rect 122469 5556 122481 5559
rect 28960 5528 122481 5556
rect 28960 5516 28966 5528
rect 122469 5525 122481 5528
rect 122515 5556 122527 5559
rect 122558 5556 122564 5568
rect 122515 5528 122564 5556
rect 122515 5525 122527 5528
rect 122469 5519 122527 5525
rect 122558 5516 122564 5528
rect 122616 5516 122622 5568
rect 212718 5516 212724 5568
rect 212776 5516 212782 5568
rect 213730 5516 213736 5568
rect 213788 5516 213794 5568
rect 215294 5516 215300 5568
rect 215352 5516 215358 5568
rect 311894 5516 311900 5568
rect 311952 5516 311958 5568
rect 1104 5466 648876 5488
rect 1104 5414 82581 5466
rect 82633 5414 82645 5466
rect 82697 5414 82709 5466
rect 82761 5414 82773 5466
rect 82825 5414 82837 5466
rect 82889 5414 244524 5466
rect 244576 5414 244588 5466
rect 244640 5414 244652 5466
rect 244704 5414 244716 5466
rect 244768 5414 244780 5466
rect 244832 5414 406467 5466
rect 406519 5414 406531 5466
rect 406583 5414 406595 5466
rect 406647 5414 406659 5466
rect 406711 5414 406723 5466
rect 406775 5414 568410 5466
rect 568462 5414 568474 5466
rect 568526 5414 568538 5466
rect 568590 5414 568602 5466
rect 568654 5414 568666 5466
rect 568718 5414 648876 5466
rect 1104 5392 648876 5414
rect 308674 5312 308680 5364
rect 308732 5352 308738 5364
rect 401137 5355 401195 5361
rect 401137 5352 401149 5355
rect 308732 5324 401149 5352
rect 308732 5312 308738 5324
rect 401137 5321 401149 5324
rect 401183 5321 401195 5355
rect 401137 5315 401195 5321
rect 216490 5244 216496 5296
rect 216548 5284 216554 5296
rect 216548 5256 224954 5284
rect 216548 5244 216554 5256
rect 203337 5219 203395 5225
rect 203337 5216 203349 5219
rect 202708 5188 203349 5216
rect 202708 5157 202736 5188
rect 203337 5185 203349 5188
rect 203383 5185 203395 5219
rect 218609 5219 218667 5225
rect 218609 5216 218621 5219
rect 203337 5179 203395 5185
rect 218072 5188 218621 5216
rect 202693 5151 202751 5157
rect 202693 5148 202705 5151
rect 180766 5120 202705 5148
rect 111334 5040 111340 5092
rect 111392 5080 111398 5092
rect 180766 5080 180794 5120
rect 202693 5117 202705 5120
rect 202739 5117 202751 5151
rect 202693 5111 202751 5117
rect 203886 5108 203892 5160
rect 203944 5108 203950 5160
rect 111392 5052 180794 5080
rect 195946 5052 209774 5080
rect 111392 5040 111398 5052
rect 126514 4972 126520 5024
rect 126572 5012 126578 5024
rect 195946 5012 195974 5052
rect 126572 4984 195974 5012
rect 209746 5012 209774 5052
rect 218072 5021 218100 5188
rect 218609 5185 218621 5188
rect 218655 5185 218667 5219
rect 218609 5179 218667 5185
rect 219158 5108 219164 5160
rect 219216 5108 219222 5160
rect 224926 5148 224954 5256
rect 262582 5244 262588 5296
rect 262640 5284 262646 5296
rect 262640 5256 354674 5284
rect 262640 5244 262646 5256
rect 309321 5219 309379 5225
rect 309321 5185 309333 5219
rect 309367 5216 309379 5219
rect 309367 5188 310008 5216
rect 309367 5185 309379 5188
rect 309321 5179 309379 5185
rect 309980 5160 310008 5188
rect 339862 5176 339868 5228
rect 339920 5176 339926 5228
rect 354646 5216 354674 5256
rect 354861 5219 354919 5225
rect 354861 5216 354873 5219
rect 354646 5188 354873 5216
rect 354861 5185 354873 5188
rect 354907 5216 354919 5219
rect 355321 5219 355379 5225
rect 355321 5216 355333 5219
rect 354907 5188 355333 5216
rect 354907 5185 354919 5188
rect 354861 5179 354919 5185
rect 355321 5185 355333 5188
rect 355367 5185 355379 5219
rect 386233 5219 386291 5225
rect 386233 5216 386245 5219
rect 355321 5179 355379 5185
rect 385696 5188 386245 5216
rect 308769 5151 308827 5157
rect 308769 5148 308781 5151
rect 224926 5120 308781 5148
rect 308769 5117 308781 5120
rect 308815 5117 308827 5151
rect 308769 5111 308827 5117
rect 309962 5108 309968 5160
rect 310020 5108 310026 5160
rect 311066 5108 311072 5160
rect 311124 5108 311130 5160
rect 338086 5120 339632 5148
rect 293310 5040 293316 5092
rect 293368 5080 293374 5092
rect 338086 5080 338114 5120
rect 293368 5052 338114 5080
rect 339604 5080 339632 5120
rect 340690 5108 340696 5160
rect 340748 5108 340754 5160
rect 355962 5108 355968 5160
rect 356020 5108 356026 5160
rect 385696 5089 385724 5188
rect 386233 5185 386245 5188
rect 386279 5185 386291 5219
rect 401152 5216 401180 5315
rect 401689 5219 401747 5225
rect 401689 5216 401701 5219
rect 401152 5188 401701 5216
rect 386233 5179 386291 5185
rect 401689 5185 401701 5188
rect 401735 5185 401747 5219
rect 401689 5179 401747 5185
rect 406657 5219 406715 5225
rect 406657 5185 406669 5219
rect 406703 5216 406715 5219
rect 406703 5188 407344 5216
rect 406703 5185 406715 5188
rect 406657 5179 406715 5185
rect 387058 5108 387064 5160
rect 387116 5108 387122 5160
rect 402514 5108 402520 5160
rect 402572 5108 402578 5160
rect 404538 5108 404544 5160
rect 404596 5148 404602 5160
rect 406105 5151 406163 5157
rect 406105 5148 406117 5151
rect 404596 5120 406117 5148
rect 404596 5108 404602 5120
rect 406105 5117 406117 5120
rect 406151 5117 406163 5151
rect 406105 5111 406163 5117
rect 385681 5083 385739 5089
rect 385681 5080 385693 5083
rect 339604 5052 385693 5080
rect 293368 5040 293374 5052
rect 385681 5049 385693 5052
rect 385727 5049 385739 5083
rect 385681 5043 385739 5049
rect 407316 5024 407344 5188
rect 432138 5176 432144 5228
rect 432196 5216 432202 5228
rect 432601 5219 432659 5225
rect 432601 5216 432613 5219
rect 432196 5188 432613 5216
rect 432196 5176 432202 5188
rect 432601 5185 432613 5188
rect 432647 5185 432659 5219
rect 447965 5219 448023 5225
rect 447965 5216 447977 5219
rect 432601 5179 432659 5185
rect 447428 5188 447977 5216
rect 433242 5108 433248 5160
rect 433300 5108 433306 5160
rect 447428 5024 447456 5188
rect 447965 5185 447977 5188
rect 448011 5185 448023 5219
rect 447965 5179 448023 5185
rect 448790 5108 448796 5160
rect 448848 5108 448854 5160
rect 218057 5015 218115 5021
rect 218057 5012 218069 5015
rect 209746 4984 218069 5012
rect 126572 4972 126578 4984
rect 218057 4981 218069 4984
rect 218103 4981 218115 5015
rect 218057 4975 218115 4981
rect 247310 4972 247316 5024
rect 247368 5012 247374 5024
rect 339313 5015 339371 5021
rect 339313 5012 339325 5015
rect 247368 4984 339325 5012
rect 247368 4972 247374 4984
rect 339313 4981 339325 4984
rect 339359 5012 339371 5015
rect 339862 5012 339868 5024
rect 339359 4984 339868 5012
rect 339359 4981 339371 4984
rect 339313 4975 339371 4981
rect 339862 4972 339868 4984
rect 339920 4972 339926 5024
rect 407298 4972 407304 5024
rect 407356 4972 407362 5024
rect 447410 4972 447416 5024
rect 447468 4972 447474 5024
rect 1104 4922 648876 4944
rect 1104 4870 81921 4922
rect 81973 4870 81985 4922
rect 82037 4870 82049 4922
rect 82101 4870 82113 4922
rect 82165 4870 82177 4922
rect 82229 4870 243864 4922
rect 243916 4870 243928 4922
rect 243980 4870 243992 4922
rect 244044 4870 244056 4922
rect 244108 4870 244120 4922
rect 244172 4870 405807 4922
rect 405859 4870 405871 4922
rect 405923 4870 405935 4922
rect 405987 4870 405999 4922
rect 406051 4870 406063 4922
rect 406115 4870 567750 4922
rect 567802 4870 567814 4922
rect 567866 4870 567878 4922
rect 567930 4870 567942 4922
rect 567994 4870 568006 4922
rect 568058 4870 648876 4922
rect 1104 4848 648876 4870
rect 233878 4768 233884 4820
rect 233936 4808 233942 4820
rect 248693 4811 248751 4817
rect 248693 4808 248705 4811
rect 233936 4780 248705 4808
rect 233936 4768 233942 4780
rect 248693 4777 248705 4780
rect 248739 4808 248751 4811
rect 249334 4808 249340 4820
rect 248739 4780 249340 4808
rect 248739 4777 248751 4780
rect 248693 4771 248751 4777
rect 249334 4768 249340 4780
rect 249392 4768 249398 4820
rect 264057 4811 264115 4817
rect 264057 4808 264069 4811
rect 258046 4780 264069 4808
rect 172238 4700 172244 4752
rect 172296 4740 172302 4752
rect 239306 4740 239312 4752
rect 172296 4712 239312 4740
rect 172296 4700 172302 4712
rect 239306 4700 239312 4712
rect 239364 4700 239370 4752
rect 239490 4700 239496 4752
rect 239548 4740 239554 4752
rect 258046 4740 258074 4780
rect 264057 4777 264069 4780
rect 264103 4808 264115 4811
rect 264698 4808 264704 4820
rect 264103 4780 264704 4808
rect 264103 4777 264115 4780
rect 264057 4771 264115 4777
rect 264698 4768 264704 4780
rect 264756 4768 264762 4820
rect 277366 4780 302234 4808
rect 239548 4712 258074 4740
rect 262784 4712 267734 4740
rect 239548 4700 239554 4712
rect 156966 4632 156972 4684
rect 157024 4672 157030 4684
rect 233878 4672 233884 4684
rect 157024 4644 233884 4672
rect 157024 4632 157030 4644
rect 233878 4632 233884 4644
rect 233936 4632 233942 4684
rect 262784 4672 262812 4712
rect 244246 4644 262812 4672
rect 263060 4644 265572 4672
rect 112625 4607 112683 4613
rect 112625 4573 112637 4607
rect 112671 4604 112683 4607
rect 113177 4607 113235 4613
rect 113177 4604 113189 4607
rect 112671 4576 113189 4604
rect 112671 4573 112683 4576
rect 112625 4567 112683 4573
rect 113177 4573 113189 4576
rect 113223 4604 113235 4607
rect 114462 4604 114468 4616
rect 113223 4576 114468 4604
rect 113223 4573 113235 4576
rect 113177 4567 113235 4573
rect 114462 4564 114468 4576
rect 114520 4564 114526 4616
rect 210697 4607 210755 4613
rect 210697 4573 210709 4607
rect 210743 4604 210755 4607
rect 211338 4604 211344 4616
rect 210743 4576 211344 4604
rect 210743 4573 210755 4576
rect 210697 4567 210755 4573
rect 211338 4564 211344 4576
rect 211396 4564 211402 4616
rect 216582 4564 216588 4616
rect 216640 4604 216646 4616
rect 244246 4604 244274 4644
rect 216640 4576 244274 4604
rect 248708 4576 249104 4604
rect 216640 4564 216646 4576
rect 23290 4496 23296 4548
rect 23348 4536 23354 4548
rect 112349 4539 112407 4545
rect 112349 4536 112361 4539
rect 23348 4508 112361 4536
rect 23348 4496 23354 4508
rect 112349 4505 112361 4508
rect 112395 4505 112407 4539
rect 112349 4499 112407 4505
rect 117958 4496 117964 4548
rect 118016 4536 118022 4548
rect 210145 4539 210203 4545
rect 210145 4536 210157 4539
rect 118016 4508 210157 4536
rect 118016 4496 118022 4508
rect 210145 4505 210157 4508
rect 210191 4505 210203 4539
rect 210145 4499 210203 4505
rect 211172 4508 212212 4536
rect 202782 4428 202788 4480
rect 202840 4468 202846 4480
rect 211172 4468 211200 4508
rect 202840 4440 211200 4468
rect 202840 4428 202846 4440
rect 211338 4428 211344 4480
rect 211396 4428 211402 4480
rect 212184 4468 212212 4508
rect 215294 4496 215300 4548
rect 215352 4536 215358 4548
rect 239398 4536 239404 4548
rect 215352 4508 239404 4536
rect 215352 4496 215358 4508
rect 239398 4496 239404 4508
rect 239456 4496 239462 4548
rect 248708 4536 248736 4576
rect 239508 4508 248736 4536
rect 239508 4468 239536 4508
rect 212184 4440 239536 4468
rect 239582 4428 239588 4480
rect 239640 4468 239646 4480
rect 248782 4468 248788 4480
rect 239640 4440 248788 4468
rect 239640 4428 239646 4440
rect 248782 4428 248788 4440
rect 248840 4428 248846 4480
rect 249076 4468 249104 4576
rect 249334 4564 249340 4616
rect 249392 4564 249398 4616
rect 249702 4496 249708 4548
rect 249760 4496 249766 4548
rect 249794 4496 249800 4548
rect 249852 4536 249858 4548
rect 263060 4536 263088 4644
rect 264698 4564 264704 4616
rect 264756 4564 264762 4616
rect 249852 4508 263088 4536
rect 249852 4496 249858 4508
rect 265250 4496 265256 4548
rect 265308 4496 265314 4548
rect 265544 4536 265572 4644
rect 267706 4604 267734 4712
rect 277366 4604 277394 4780
rect 267706 4576 277394 4604
rect 291856 4712 297404 4740
rect 291856 4536 291884 4712
rect 294785 4607 294843 4613
rect 294785 4604 294797 4607
rect 265544 4508 291884 4536
rect 292500 4576 294797 4604
rect 292500 4468 292528 4576
rect 294785 4573 294797 4576
rect 294831 4604 294843 4607
rect 295429 4607 295487 4613
rect 295429 4604 295441 4607
rect 294831 4576 295441 4604
rect 294831 4573 294843 4576
rect 294785 4567 294843 4573
rect 295429 4573 295441 4576
rect 295475 4573 295487 4607
rect 297376 4604 297404 4712
rect 302206 4672 302234 4780
rect 407298 4768 407304 4820
rect 407356 4808 407362 4820
rect 499942 4808 499948 4820
rect 407356 4780 499948 4808
rect 407356 4768 407362 4780
rect 499942 4768 499948 4780
rect 500000 4768 500006 4820
rect 339402 4700 339408 4752
rect 339460 4740 339466 4752
rect 432138 4740 432144 4752
rect 339460 4712 432144 4740
rect 339460 4700 339466 4712
rect 432138 4700 432144 4712
rect 432196 4700 432202 4752
rect 309318 4672 309324 4684
rect 302206 4644 309324 4672
rect 309318 4632 309324 4644
rect 309376 4672 309382 4684
rect 309376 4644 309548 4672
rect 309376 4632 309382 4644
rect 308585 4607 308643 4613
rect 297376 4576 302234 4604
rect 295429 4567 295487 4573
rect 295978 4496 295984 4548
rect 296036 4496 296042 4548
rect 302206 4536 302234 4576
rect 308585 4573 308597 4607
rect 308631 4604 308643 4607
rect 308858 4604 308864 4616
rect 308631 4576 308864 4604
rect 308631 4573 308643 4576
rect 308585 4567 308643 4573
rect 308858 4564 308864 4576
rect 308916 4564 308922 4616
rect 309520 4613 309548 4644
rect 354582 4632 354588 4684
rect 354640 4672 354646 4684
rect 447410 4672 447416 4684
rect 354640 4644 447416 4672
rect 354640 4632 354646 4644
rect 447410 4632 447416 4644
rect 447468 4632 447474 4684
rect 309505 4607 309563 4613
rect 309505 4573 309517 4607
rect 309551 4573 309563 4607
rect 309505 4567 309563 4573
rect 310790 4564 310796 4616
rect 310848 4604 310854 4616
rect 311069 4607 311127 4613
rect 311069 4604 311081 4607
rect 310848 4576 311081 4604
rect 310848 4564 310854 4576
rect 311069 4573 311081 4576
rect 311115 4573 311127 4607
rect 311069 4567 311127 4573
rect 405185 4607 405243 4613
rect 405185 4573 405197 4607
rect 405231 4604 405243 4607
rect 405231 4576 405964 4604
rect 405231 4573 405243 4576
rect 405185 4567 405243 4573
rect 308033 4539 308091 4545
rect 308033 4536 308045 4539
rect 302206 4508 308045 4536
rect 308033 4505 308045 4508
rect 308079 4505 308091 4539
rect 308033 4499 308091 4505
rect 310330 4496 310336 4548
rect 310388 4496 310394 4548
rect 311618 4496 311624 4548
rect 311676 4496 311682 4548
rect 311894 4496 311900 4548
rect 311952 4536 311958 4548
rect 404633 4539 404691 4545
rect 404633 4536 404645 4539
rect 311952 4508 404645 4536
rect 311952 4496 311958 4508
rect 404633 4505 404645 4508
rect 404679 4505 404691 4539
rect 404633 4499 404691 4505
rect 249076 4440 292528 4468
rect 313734 4428 313740 4480
rect 313792 4468 313798 4480
rect 404538 4468 404544 4480
rect 313792 4440 404544 4468
rect 313792 4428 313798 4440
rect 404538 4428 404544 4440
rect 404596 4428 404602 4480
rect 405936 4477 405964 4576
rect 405921 4471 405979 4477
rect 405921 4437 405933 4471
rect 405967 4468 405979 4471
rect 406194 4468 406200 4480
rect 405967 4440 406200 4468
rect 405967 4437 405979 4440
rect 405921 4431 405979 4437
rect 406194 4428 406200 4440
rect 406252 4428 406258 4480
rect 1104 4378 648876 4400
rect 1104 4326 82581 4378
rect 82633 4326 82645 4378
rect 82697 4326 82709 4378
rect 82761 4326 82773 4378
rect 82825 4326 82837 4378
rect 82889 4326 244524 4378
rect 244576 4326 244588 4378
rect 244640 4326 244652 4378
rect 244704 4326 244716 4378
rect 244768 4326 244780 4378
rect 244832 4326 406467 4378
rect 406519 4326 406531 4378
rect 406583 4326 406595 4378
rect 406647 4326 406659 4378
rect 406711 4326 406723 4378
rect 406775 4326 568410 4378
rect 568462 4326 568474 4378
rect 568526 4326 568538 4378
rect 568590 4326 568602 4378
rect 568654 4326 568666 4378
rect 568718 4326 648876 4378
rect 1104 4304 648876 4326
rect 248782 4224 248788 4276
rect 248840 4264 248846 4276
rect 249794 4264 249800 4276
rect 248840 4236 249800 4264
rect 248840 4224 248846 4236
rect 249794 4224 249800 4236
rect 249852 4224 249858 4276
rect 309318 4224 309324 4276
rect 309376 4224 309382 4276
rect 218422 4156 218428 4208
rect 218480 4196 218486 4208
rect 310790 4196 310796 4208
rect 218480 4168 310796 4196
rect 218480 4156 218486 4168
rect 310790 4156 310796 4168
rect 310848 4156 310854 4208
rect 356808 4168 357020 4196
rect 248966 4088 248972 4140
rect 249024 4128 249030 4140
rect 249024 4100 306420 4128
rect 249024 4088 249030 4100
rect 264330 4020 264336 4072
rect 264388 4060 264394 4072
rect 264388 4032 294644 4060
rect 264388 4020 264394 4032
rect 213730 3952 213736 4004
rect 213788 3992 213794 4004
rect 294616 3992 294644 4032
rect 296714 4020 296720 4072
rect 296772 4060 296778 4072
rect 305917 4063 305975 4069
rect 305917 4060 305929 4063
rect 296772 4032 305929 4060
rect 296772 4020 296778 4032
rect 305917 4029 305929 4032
rect 305963 4029 305975 4063
rect 306392 4060 306420 4100
rect 306466 4088 306472 4140
rect 306524 4088 306530 4140
rect 341334 4128 341340 4140
rect 306576 4100 341340 4128
rect 306576 4060 306604 4100
rect 341334 4088 341340 4100
rect 341392 4128 341398 4140
rect 341521 4131 341579 4137
rect 341521 4128 341533 4131
rect 341392 4100 341533 4128
rect 341392 4088 341398 4100
rect 341521 4097 341533 4100
rect 341567 4097 341579 4131
rect 341521 4091 341579 4097
rect 342180 4100 350534 4128
rect 306392 4032 306604 4060
rect 306668 4032 331214 4060
rect 305917 4023 305975 4029
rect 306668 3992 306696 4032
rect 213788 3964 289814 3992
rect 294616 3964 306696 3992
rect 213788 3952 213794 3964
rect 289786 3924 289814 3964
rect 307018 3952 307024 4004
rect 307076 3992 307082 4004
rect 331186 3992 331214 4032
rect 340690 4020 340696 4072
rect 340748 4060 340754 4072
rect 342070 4060 342076 4072
rect 340748 4032 342076 4060
rect 340748 4020 340754 4032
rect 342070 4020 342076 4032
rect 342128 4020 342134 4072
rect 342180 3992 342208 4100
rect 342714 4020 342720 4072
rect 342772 4020 342778 4072
rect 350506 4060 350534 4100
rect 355962 4088 355968 4140
rect 356020 4128 356026 4140
rect 356808 4128 356836 4168
rect 356020 4100 356836 4128
rect 356885 4131 356943 4137
rect 356020 4088 356026 4100
rect 356885 4097 356897 4131
rect 356931 4097 356943 4131
rect 356992 4128 357020 4168
rect 434088 4168 434300 4196
rect 356992 4100 373994 4128
rect 356885 4091 356943 4097
rect 356241 4063 356299 4069
rect 356241 4060 356253 4063
rect 350506 4032 356253 4060
rect 356241 4029 356253 4032
rect 356287 4060 356299 4063
rect 356900 4060 356928 4091
rect 356287 4032 356928 4060
rect 356287 4029 356299 4032
rect 356241 4023 356299 4029
rect 358078 4020 358084 4072
rect 358136 4020 358142 4072
rect 373966 4060 373994 4100
rect 387794 4088 387800 4140
rect 387852 4088 387858 4140
rect 387904 4100 393314 4128
rect 387904 4060 387932 4100
rect 373966 4032 387932 4060
rect 388990 4020 388996 4072
rect 389048 4020 389054 4072
rect 393286 4060 393314 4100
rect 402606 4088 402612 4140
rect 402664 4128 402670 4140
rect 403253 4131 403311 4137
rect 403253 4128 403265 4131
rect 402664 4100 403265 4128
rect 402664 4088 402670 4100
rect 403253 4097 403265 4100
rect 403299 4097 403311 4131
rect 434088 4128 434116 4168
rect 403253 4091 403311 4097
rect 404372 4100 434116 4128
rect 434165 4131 434223 4137
rect 404372 4060 404400 4100
rect 434165 4097 434177 4131
rect 434211 4097 434223 4131
rect 434272 4128 434300 4168
rect 499942 4156 499948 4208
rect 500000 4156 500006 4208
rect 448977 4131 449035 4137
rect 448977 4128 448989 4131
rect 434272 4100 448989 4128
rect 434165 4091 434223 4097
rect 448977 4097 448989 4100
rect 449023 4128 449035 4131
rect 449621 4131 449679 4137
rect 449621 4128 449633 4131
rect 449023 4100 449633 4128
rect 449023 4097 449035 4100
rect 448977 4091 449035 4097
rect 449621 4097 449633 4100
rect 449667 4097 449679 4131
rect 449621 4091 449679 4097
rect 393286 4032 404400 4060
rect 404446 4020 404452 4072
rect 404504 4020 404510 4072
rect 307076 3964 311894 3992
rect 331186 3964 342208 3992
rect 307076 3952 307082 3964
rect 296714 3924 296720 3936
rect 289786 3896 296720 3924
rect 296714 3884 296720 3896
rect 296772 3884 296778 3936
rect 306466 3884 306472 3936
rect 306524 3924 306530 3936
rect 307110 3924 307116 3936
rect 306524 3896 307116 3924
rect 306524 3884 306530 3896
rect 307110 3884 307116 3896
rect 307168 3884 307174 3936
rect 308858 3884 308864 3936
rect 308916 3884 308922 3936
rect 311866 3924 311894 3964
rect 342254 3952 342260 4004
rect 342312 3992 342318 4004
rect 433521 3995 433579 4001
rect 433521 3992 433533 3995
rect 342312 3964 433533 3992
rect 342312 3952 342318 3964
rect 433521 3961 433533 3964
rect 433567 3992 433579 3995
rect 434180 3992 434208 4091
rect 479886 4088 479892 4140
rect 479944 4128 479950 4140
rect 480533 4131 480591 4137
rect 480533 4128 480545 4131
rect 479944 4100 480545 4128
rect 479944 4088 479950 4100
rect 480533 4097 480545 4100
rect 480579 4097 480591 4131
rect 480533 4091 480591 4097
rect 480916 4100 489914 4128
rect 435358 4020 435364 4072
rect 435416 4020 435422 4072
rect 450814 4020 450820 4072
rect 450872 4020 450878 4072
rect 480916 4060 480944 4100
rect 451246 4032 480944 4060
rect 481729 4063 481787 4069
rect 451246 3992 451274 4032
rect 481729 4029 481741 4063
rect 481775 4060 481787 4063
rect 489886 4060 489914 4100
rect 495434 4088 495440 4140
rect 495492 4128 495498 4140
rect 495989 4131 496047 4137
rect 495989 4128 496001 4131
rect 495492 4100 496001 4128
rect 495492 4088 495498 4100
rect 495989 4097 496001 4100
rect 496035 4097 496047 4131
rect 495989 4091 496047 4097
rect 496096 4100 499574 4128
rect 496096 4060 496124 4100
rect 481775 4032 485774 4060
rect 489886 4032 496124 4060
rect 481775 4029 481787 4032
rect 481729 4023 481787 4029
rect 433567 3964 434208 3992
rect 441586 3964 451274 3992
rect 485746 3992 485774 4032
rect 497182 4020 497188 4072
rect 497240 4020 497246 4072
rect 499546 4060 499574 4100
rect 500494 4088 500500 4140
rect 500552 4088 500558 4140
rect 526901 4131 526959 4137
rect 526901 4097 526913 4131
rect 526947 4097 526959 4131
rect 526901 4091 526959 4097
rect 526257 4063 526315 4069
rect 526257 4060 526269 4063
rect 499546 4032 526269 4060
rect 526257 4029 526269 4032
rect 526303 4060 526315 4063
rect 526916 4060 526944 4091
rect 526303 4032 526944 4060
rect 528097 4063 528155 4069
rect 526303 4029 526315 4032
rect 526257 4023 526315 4029
rect 528097 4029 528109 4063
rect 528143 4060 528155 4063
rect 619818 4060 619824 4072
rect 528143 4032 619824 4060
rect 528143 4029 528155 4032
rect 528097 4023 528155 4029
rect 619818 4020 619824 4032
rect 619876 4020 619882 4072
rect 573450 3992 573456 4004
rect 485746 3964 573456 3992
rect 433567 3961 433579 3964
rect 433521 3955 433579 3961
rect 387153 3927 387211 3933
rect 387153 3924 387165 3927
rect 311866 3896 387165 3924
rect 387153 3893 387165 3896
rect 387199 3924 387211 3927
rect 387794 3924 387800 3936
rect 387199 3896 387800 3924
rect 387199 3893 387211 3896
rect 387153 3887 387211 3893
rect 387794 3884 387800 3896
rect 387852 3884 387858 3936
rect 402606 3884 402612 3936
rect 402664 3884 402670 3936
rect 433242 3884 433248 3936
rect 433300 3924 433306 3936
rect 441586 3924 441614 3964
rect 573450 3952 573456 3964
rect 573508 3952 573514 4004
rect 433300 3896 441614 3924
rect 433300 3884 433306 3896
rect 479886 3884 479892 3936
rect 479944 3884 479950 3936
rect 495434 3884 495440 3936
rect 495492 3884 495498 3936
rect 500494 3884 500500 3936
rect 500552 3924 500558 3936
rect 501233 3927 501291 3933
rect 501233 3924 501245 3927
rect 500552 3896 501245 3924
rect 500552 3884 500558 3896
rect 501233 3893 501245 3896
rect 501279 3924 501291 3927
rect 594058 3924 594064 3936
rect 501279 3896 594064 3924
rect 501279 3893 501291 3896
rect 501233 3887 501291 3893
rect 594058 3884 594064 3896
rect 594116 3884 594122 3936
rect 1104 3834 648876 3856
rect 1104 3782 81921 3834
rect 81973 3782 81985 3834
rect 82037 3782 82049 3834
rect 82101 3782 82113 3834
rect 82165 3782 82177 3834
rect 82229 3782 243864 3834
rect 243916 3782 243928 3834
rect 243980 3782 243992 3834
rect 244044 3782 244056 3834
rect 244108 3782 244120 3834
rect 244172 3782 405807 3834
rect 405859 3782 405871 3834
rect 405923 3782 405935 3834
rect 405987 3782 405999 3834
rect 406051 3782 406063 3834
rect 406115 3782 567750 3834
rect 567802 3782 567814 3834
rect 567866 3782 567878 3834
rect 567930 3782 567942 3834
rect 567994 3782 568006 3834
rect 568058 3782 648876 3834
rect 1104 3760 648876 3782
rect 295058 3680 295064 3732
rect 295116 3720 295122 3732
rect 307018 3720 307024 3732
rect 295116 3692 307024 3720
rect 295116 3680 295122 3692
rect 307018 3680 307024 3692
rect 307076 3680 307082 3732
rect 310330 3680 310336 3732
rect 310388 3720 310394 3732
rect 402606 3720 402612 3732
rect 310388 3692 402612 3720
rect 310388 3680 310394 3692
rect 402606 3680 402612 3692
rect 402664 3680 402670 3732
rect 404446 3680 404452 3732
rect 404504 3720 404510 3732
rect 496170 3720 496176 3732
rect 404504 3692 496176 3720
rect 404504 3680 404510 3692
rect 496170 3680 496176 3692
rect 496228 3680 496234 3732
rect 497182 3680 497188 3732
rect 497240 3720 497246 3732
rect 588906 3720 588912 3732
rect 497240 3692 588912 3720
rect 497240 3680 497246 3692
rect 588906 3680 588912 3692
rect 588964 3680 588970 3732
rect 295978 3612 295984 3664
rect 296036 3652 296042 3664
rect 387978 3652 387984 3664
rect 296036 3624 309134 3652
rect 296036 3612 296042 3624
rect 309106 3584 309134 3624
rect 318766 3624 387984 3652
rect 318766 3584 318794 3624
rect 387978 3612 387984 3624
rect 388036 3612 388042 3664
rect 309106 3556 318794 3584
rect 341334 3544 341340 3596
rect 341392 3544 341398 3596
rect 387058 3544 387064 3596
rect 387116 3584 387122 3596
rect 479886 3584 479892 3596
rect 387116 3556 479892 3584
rect 387116 3544 387122 3556
rect 479886 3544 479892 3556
rect 479944 3544 479950 3596
rect 208397 3519 208455 3525
rect 208397 3485 208409 3519
rect 208443 3516 208455 3519
rect 208949 3519 209007 3525
rect 208949 3516 208961 3519
rect 208443 3488 208961 3516
rect 208443 3485 208455 3488
rect 208397 3479 208455 3485
rect 208949 3485 208961 3488
rect 208995 3516 209007 3519
rect 233602 3516 233608 3528
rect 208995 3488 233608 3516
rect 208995 3485 209007 3488
rect 208949 3479 209007 3485
rect 233602 3476 233608 3488
rect 233660 3476 233666 3528
rect 311066 3476 311072 3528
rect 311124 3516 311130 3528
rect 402793 3519 402851 3525
rect 311124 3488 402376 3516
rect 311124 3476 311130 3488
rect 117406 3408 117412 3460
rect 117464 3448 117470 3460
rect 208121 3451 208179 3457
rect 208121 3448 208133 3451
rect 117464 3420 208133 3448
rect 117464 3408 117470 3420
rect 208121 3417 208133 3420
rect 208167 3417 208179 3451
rect 208121 3411 208179 3417
rect 309962 3408 309968 3460
rect 310020 3448 310026 3460
rect 402241 3451 402299 3457
rect 402241 3448 402253 3451
rect 310020 3420 402253 3448
rect 310020 3408 310026 3420
rect 402241 3417 402253 3420
rect 402287 3417 402299 3451
rect 402348 3448 402376 3488
rect 402793 3485 402805 3519
rect 402839 3516 402851 3519
rect 403342 3516 403348 3528
rect 402839 3488 403348 3516
rect 402839 3485 402851 3488
rect 402793 3479 402851 3485
rect 403342 3476 403348 3488
rect 403400 3476 403406 3528
rect 404173 3519 404231 3525
rect 404173 3485 404185 3519
rect 404219 3516 404231 3519
rect 404817 3519 404875 3525
rect 404817 3516 404829 3519
rect 404219 3488 404829 3516
rect 404219 3485 404231 3488
rect 404173 3479 404231 3485
rect 404817 3485 404829 3488
rect 404863 3516 404875 3519
rect 497274 3516 497280 3528
rect 404863 3488 497280 3516
rect 404863 3485 404875 3488
rect 404817 3479 404875 3485
rect 497274 3476 497280 3488
rect 497332 3476 497338 3528
rect 499209 3519 499267 3525
rect 499209 3485 499221 3519
rect 499255 3516 499267 3519
rect 499850 3516 499856 3528
rect 499255 3488 499856 3516
rect 499255 3485 499267 3488
rect 499209 3479 499267 3485
rect 499850 3476 499856 3488
rect 499908 3476 499914 3528
rect 541897 3519 541955 3525
rect 541897 3516 541909 3519
rect 541360 3488 541909 3516
rect 403621 3451 403679 3457
rect 403621 3448 403633 3451
rect 402348 3420 403633 3448
rect 402241 3411 402299 3417
rect 403621 3417 403633 3420
rect 403667 3417 403679 3451
rect 403621 3411 403679 3417
rect 404648 3420 404860 3448
rect 342714 3340 342720 3392
rect 342772 3380 342778 3392
rect 404648 3380 404676 3420
rect 342772 3352 404676 3380
rect 404832 3380 404860 3420
rect 406194 3408 406200 3460
rect 406252 3448 406258 3460
rect 498657 3451 498715 3457
rect 498657 3448 498669 3451
rect 406252 3420 498669 3448
rect 406252 3408 406258 3420
rect 498657 3417 498669 3420
rect 498703 3417 498715 3451
rect 498657 3411 498715 3417
rect 499546 3420 509234 3448
rect 434346 3380 434352 3392
rect 404832 3352 434352 3380
rect 342772 3340 342778 3352
rect 434346 3340 434352 3352
rect 434404 3340 434410 3392
rect 448790 3340 448796 3392
rect 448848 3380 448854 3392
rect 499546 3380 499574 3420
rect 448848 3352 499574 3380
rect 448848 3340 448854 3352
rect 499850 3340 499856 3392
rect 499908 3340 499914 3392
rect 509206 3380 509234 3420
rect 541360 3389 541388 3488
rect 541897 3485 541909 3488
rect 541943 3485 541955 3519
rect 541897 3479 541955 3485
rect 543093 3451 543151 3457
rect 543093 3417 543105 3451
rect 543139 3448 543151 3451
rect 635274 3448 635280 3460
rect 543139 3420 635280 3448
rect 543139 3417 543151 3420
rect 543093 3411 543151 3417
rect 635274 3408 635280 3420
rect 635332 3408 635338 3460
rect 541345 3383 541403 3389
rect 541345 3380 541357 3383
rect 509206 3352 541357 3380
rect 541345 3349 541357 3352
rect 541391 3349 541403 3383
rect 541345 3343 541403 3349
rect 1104 3290 648876 3312
rect 1104 3238 82581 3290
rect 82633 3238 82645 3290
rect 82697 3238 82709 3290
rect 82761 3238 82773 3290
rect 82825 3238 82837 3290
rect 82889 3238 244524 3290
rect 244576 3238 244588 3290
rect 244640 3238 244652 3290
rect 244704 3238 244716 3290
rect 244768 3238 244780 3290
rect 244832 3238 406467 3290
rect 406519 3238 406531 3290
rect 406583 3238 406595 3290
rect 406647 3238 406659 3290
rect 406711 3238 406723 3290
rect 406775 3238 568410 3290
rect 568462 3238 568474 3290
rect 568526 3238 568538 3290
rect 568590 3238 568602 3290
rect 568654 3238 568666 3290
rect 568718 3238 648876 3290
rect 1104 3216 648876 3238
rect 32490 3136 32496 3188
rect 32548 3136 32554 3188
rect 112346 3136 112352 3188
rect 112404 3176 112410 3188
rect 202506 3176 202512 3188
rect 112404 3148 202512 3176
rect 112404 3136 112410 3148
rect 202506 3136 202512 3148
rect 202564 3136 202570 3188
rect 203886 3136 203892 3188
rect 203944 3176 203950 3188
rect 295337 3179 295395 3185
rect 295337 3176 295349 3179
rect 203944 3148 295349 3176
rect 203944 3136 203950 3148
rect 295337 3145 295349 3148
rect 295383 3176 295395 3179
rect 295702 3176 295708 3188
rect 295383 3148 295708 3176
rect 295383 3145 295395 3148
rect 295337 3139 295395 3145
rect 295702 3136 295708 3148
rect 295760 3136 295766 3188
rect 304810 3176 304816 3188
rect 299446 3148 304816 3176
rect 22002 3068 22008 3120
rect 22060 3108 22066 3120
rect 109773 3111 109831 3117
rect 109773 3108 109785 3111
rect 22060 3080 109785 3108
rect 22060 3068 22066 3080
rect 109773 3077 109785 3080
rect 109819 3108 109831 3111
rect 110230 3108 110236 3120
rect 109819 3080 110236 3108
rect 109819 3077 109831 3080
rect 109773 3071 109831 3077
rect 110230 3068 110236 3080
rect 110288 3068 110294 3120
rect 173250 3068 173256 3120
rect 173308 3108 173314 3120
rect 264333 3111 264391 3117
rect 264333 3108 264345 3111
rect 173308 3080 264345 3108
rect 173308 3068 173314 3080
rect 264333 3077 264345 3080
rect 264379 3108 264391 3111
rect 264790 3108 264796 3120
rect 264379 3080 264796 3108
rect 264379 3077 264391 3080
rect 264333 3071 264391 3077
rect 264790 3068 264796 3080
rect 264848 3068 264854 3120
rect 265250 3068 265256 3120
rect 265308 3108 265314 3120
rect 299446 3108 299474 3148
rect 304810 3136 304816 3148
rect 304868 3136 304874 3188
rect 305457 3179 305515 3185
rect 305457 3145 305469 3179
rect 305503 3176 305515 3179
rect 326338 3176 326344 3188
rect 305503 3148 326344 3176
rect 305503 3145 305515 3148
rect 305457 3139 305515 3145
rect 305472 3108 305500 3139
rect 326338 3136 326344 3148
rect 326396 3136 326402 3188
rect 358078 3136 358084 3188
rect 358136 3176 358142 3188
rect 449897 3179 449955 3185
rect 449897 3176 449909 3179
rect 358136 3148 449909 3176
rect 358136 3136 358142 3148
rect 449897 3145 449909 3148
rect 449943 3176 449955 3179
rect 450262 3176 450268 3188
rect 449943 3148 450268 3176
rect 449943 3145 449955 3148
rect 449897 3139 449955 3145
rect 450262 3136 450268 3148
rect 450320 3136 450326 3188
rect 450814 3136 450820 3188
rect 450872 3176 450878 3188
rect 542541 3179 542599 3185
rect 542541 3176 542553 3179
rect 450872 3148 542553 3176
rect 450872 3136 450878 3148
rect 542541 3145 542553 3148
rect 542587 3176 542599 3179
rect 542998 3176 543004 3188
rect 542587 3148 543004 3176
rect 542587 3145 542599 3148
rect 542541 3139 542599 3145
rect 542998 3136 543004 3148
rect 543056 3136 543062 3188
rect 573450 3136 573456 3188
rect 573508 3136 573514 3188
rect 588906 3136 588912 3188
rect 588964 3136 588970 3188
rect 619818 3136 619824 3188
rect 619876 3136 619882 3188
rect 635274 3136 635280 3188
rect 635332 3136 635338 3188
rect 357066 3108 357072 3120
rect 265308 3080 299474 3108
rect 304644 3080 305500 3108
rect 305564 3080 357072 3108
rect 265308 3068 265314 3080
rect 37734 3000 37740 3052
rect 37792 3040 37798 3052
rect 125226 3040 125232 3052
rect 37792 3012 125232 3040
rect 37792 3000 37798 3012
rect 125226 3000 125232 3012
rect 125284 3000 125290 3052
rect 127526 3000 127532 3052
rect 127584 3040 127590 3052
rect 218057 3043 218115 3049
rect 218057 3040 218069 3043
rect 127584 3012 218069 3040
rect 127584 3000 127590 3012
rect 218057 3009 218069 3012
rect 218103 3040 218115 3043
rect 218422 3040 218428 3052
rect 218103 3012 218428 3040
rect 218103 3009 218115 3012
rect 218057 3003 218115 3009
rect 218422 3000 218428 3012
rect 218480 3000 218486 3052
rect 219158 3000 219164 3052
rect 219216 3040 219222 3052
rect 304644 3049 304672 3080
rect 304629 3043 304687 3049
rect 219216 3012 304580 3040
rect 219216 3000 219222 3012
rect 21910 2932 21916 2984
rect 21968 2972 21974 2984
rect 78861 2975 78919 2981
rect 78861 2972 78873 2975
rect 21968 2944 78873 2972
rect 21968 2932 21974 2944
rect 78861 2941 78873 2944
rect 78907 2972 78919 2975
rect 79318 2972 79324 2984
rect 78907 2944 79324 2972
rect 78907 2941 78919 2944
rect 78861 2935 78919 2941
rect 79318 2932 79324 2944
rect 79376 2932 79382 2984
rect 82446 2932 82452 2984
rect 82504 2972 82510 2984
rect 171597 2975 171655 2981
rect 171597 2972 171609 2975
rect 82504 2944 171609 2972
rect 82504 2932 82510 2944
rect 171597 2941 171609 2944
rect 171643 2972 171655 2975
rect 172054 2972 172060 2984
rect 171643 2944 172060 2972
rect 171643 2941 171655 2944
rect 171597 2935 171655 2941
rect 172054 2932 172060 2944
rect 172112 2932 172118 2984
rect 212718 2932 212724 2984
rect 212776 2972 212782 2984
rect 304353 2975 304411 2981
rect 304353 2972 304365 2975
rect 212776 2944 304365 2972
rect 212776 2932 212782 2944
rect 304353 2941 304365 2944
rect 304399 2941 304411 2975
rect 304552 2972 304580 3012
rect 304629 3009 304641 3043
rect 304675 3009 304687 3043
rect 304629 3003 304687 3009
rect 304810 3000 304816 3052
rect 304868 3040 304874 3052
rect 305564 3040 305592 3080
rect 357066 3068 357072 3080
rect 357124 3068 357130 3120
rect 387978 3068 387984 3120
rect 388036 3068 388042 3120
rect 400876 3080 401732 3108
rect 304868 3012 305592 3040
rect 304868 3000 304874 3012
rect 308858 3000 308864 3052
rect 308916 3040 308922 3052
rect 308916 3012 311894 3040
rect 308916 3000 308922 3012
rect 310701 2975 310759 2981
rect 310701 2972 310713 2975
rect 304552 2944 310713 2972
rect 304353 2935 304411 2941
rect 310701 2941 310713 2944
rect 310747 2972 310759 2975
rect 311158 2972 311164 2984
rect 310747 2944 311164 2972
rect 310747 2941 310759 2944
rect 310701 2935 310759 2941
rect 311158 2932 311164 2944
rect 311216 2932 311222 2984
rect 311866 2972 311894 3012
rect 400769 2975 400827 2981
rect 400769 2972 400781 2975
rect 311866 2944 400781 2972
rect 400769 2941 400781 2944
rect 400815 2941 400827 2975
rect 400769 2935 400827 2941
rect 21266 2864 21272 2916
rect 21324 2904 21330 2916
rect 63497 2907 63555 2913
rect 63497 2904 63509 2907
rect 21324 2876 63509 2904
rect 21324 2864 21330 2876
rect 63497 2873 63509 2876
rect 63543 2904 63555 2907
rect 63862 2904 63868 2916
rect 63543 2876 63868 2904
rect 63543 2873 63555 2876
rect 63497 2867 63555 2873
rect 63862 2864 63868 2876
rect 63920 2864 63926 2916
rect 66714 2864 66720 2916
rect 66772 2904 66778 2916
rect 156141 2907 156199 2913
rect 156141 2904 156153 2907
rect 66772 2876 156153 2904
rect 66772 2864 66778 2876
rect 156141 2873 156153 2876
rect 156187 2904 156199 2907
rect 156598 2904 156604 2916
rect 156187 2876 156604 2904
rect 156187 2873 156199 2876
rect 156141 2867 156199 2873
rect 156598 2864 156604 2876
rect 156656 2864 156662 2916
rect 157886 2864 157892 2916
rect 157944 2904 157950 2916
rect 157944 2876 234614 2904
rect 157944 2864 157950 2876
rect 1578 2796 1584 2848
rect 1636 2796 1642 2848
rect 47946 2796 47952 2848
rect 48004 2796 48010 2848
rect 94314 2796 94320 2848
rect 94372 2796 94378 2848
rect 140777 2839 140835 2845
rect 140777 2805 140789 2839
rect 140823 2836 140835 2839
rect 141050 2836 141056 2848
rect 140823 2808 141056 2836
rect 140823 2805 140835 2808
rect 140777 2799 140835 2805
rect 141050 2796 141056 2808
rect 141108 2796 141114 2848
rect 186866 2796 186872 2848
rect 186924 2796 186930 2848
rect 233513 2839 233571 2845
rect 233513 2805 233525 2839
rect 233559 2836 233571 2839
rect 233786 2836 233792 2848
rect 233559 2808 233792 2836
rect 233559 2805 233571 2808
rect 233513 2799 233571 2805
rect 233786 2796 233792 2808
rect 233844 2796 233850 2848
rect 234586 2836 234614 2876
rect 249702 2864 249708 2916
rect 249760 2904 249766 2916
rect 249760 2876 331214 2904
rect 249760 2864 249766 2876
rect 248877 2839 248935 2845
rect 248877 2836 248889 2839
rect 234586 2808 248889 2836
rect 248877 2805 248889 2808
rect 248923 2836 248935 2839
rect 248966 2836 248972 2848
rect 248923 2808 248972 2836
rect 248923 2805 248935 2808
rect 248877 2799 248935 2805
rect 248966 2796 248972 2808
rect 249024 2796 249030 2848
rect 279602 2796 279608 2848
rect 279660 2796 279666 2848
rect 326249 2839 326307 2845
rect 326249 2805 326261 2839
rect 326295 2836 326307 2839
rect 326522 2836 326528 2848
rect 326295 2808 326528 2836
rect 326295 2805 326307 2808
rect 326249 2799 326307 2805
rect 326522 2796 326528 2808
rect 326580 2796 326586 2848
rect 331186 2836 331214 2876
rect 388990 2864 388996 2916
rect 389048 2904 389054 2916
rect 400876 2904 400904 3080
rect 401045 3043 401103 3049
rect 401045 3009 401057 3043
rect 401091 3040 401103 3043
rect 401091 3012 401640 3040
rect 401091 3009 401103 3012
rect 401045 3003 401103 3009
rect 389048 2876 400904 2904
rect 389048 2864 389054 2876
rect 341705 2839 341763 2845
rect 341705 2836 341717 2839
rect 331186 2808 341717 2836
rect 341705 2805 341717 2808
rect 341751 2836 341763 2839
rect 342070 2836 342076 2848
rect 341751 2808 342076 2836
rect 341751 2805 341763 2808
rect 341705 2799 341763 2805
rect 342070 2796 342076 2808
rect 342128 2796 342134 2848
rect 372614 2796 372620 2848
rect 372672 2796 372678 2848
rect 401612 2845 401640 3012
rect 401704 2904 401732 3080
rect 434346 3068 434352 3120
rect 434404 3068 434410 3120
rect 435358 3068 435364 3120
rect 435416 3108 435422 3120
rect 527177 3111 527235 3117
rect 527177 3108 527189 3111
rect 435416 3080 527189 3108
rect 435416 3068 435422 3080
rect 527177 3077 527189 3080
rect 527223 3108 527235 3111
rect 527542 3108 527548 3120
rect 527223 3080 527548 3108
rect 527223 3077 527235 3080
rect 527177 3071 527235 3077
rect 527542 3068 527548 3080
rect 527600 3068 527606 3120
rect 594058 3068 594064 3120
rect 594116 3068 594122 3120
rect 402514 3000 402520 3052
rect 402572 3040 402578 3052
rect 495434 3040 495440 3052
rect 402572 3012 495440 3040
rect 402572 3000 402578 3012
rect 495434 3000 495440 3012
rect 495492 3000 495498 3052
rect 496170 3000 496176 3052
rect 496228 3000 496234 3052
rect 497274 3000 497280 3052
rect 497332 3000 497338 3052
rect 497553 3043 497611 3049
rect 497553 3009 497565 3043
rect 497599 3040 497611 3043
rect 510522 3040 510528 3052
rect 497599 3012 510528 3040
rect 497599 3009 497611 3012
rect 497553 3003 497611 3009
rect 510522 3000 510528 3012
rect 510580 3000 510586 3052
rect 594337 3043 594395 3049
rect 594337 3009 594349 3043
rect 594383 3040 594395 3043
rect 602890 3040 602896 3052
rect 594383 3012 602896 3040
rect 594383 3009 594395 3012
rect 594337 3003 594395 3009
rect 602890 3000 602896 3012
rect 602948 3000 602954 3052
rect 403342 2932 403348 2984
rect 403400 2932 403406 2984
rect 401704 2876 470594 2904
rect 401597 2839 401655 2845
rect 401597 2805 401609 2839
rect 401643 2836 401655 2839
rect 415302 2836 415308 2848
rect 401643 2808 415308 2836
rect 401643 2805 401655 2808
rect 401597 2799 401655 2805
rect 415302 2796 415308 2808
rect 415360 2796 415366 2848
rect 465258 2796 465264 2848
rect 465316 2796 465322 2848
rect 470566 2836 470594 2876
rect 480717 2839 480775 2845
rect 480717 2836 480729 2839
rect 470566 2808 480729 2836
rect 480717 2805 480729 2808
rect 480763 2836 480775 2839
rect 480806 2836 480812 2848
rect 480763 2808 480812 2836
rect 480763 2805 480775 2808
rect 480717 2799 480775 2805
rect 480806 2796 480812 2808
rect 480864 2796 480870 2848
rect 557994 2796 558000 2848
rect 558052 2796 558058 2848
rect 1104 2746 648876 2768
rect 1104 2694 81921 2746
rect 81973 2694 81985 2746
rect 82037 2694 82049 2746
rect 82101 2694 82113 2746
rect 82165 2694 82177 2746
rect 82229 2694 243864 2746
rect 243916 2694 243928 2746
rect 243980 2694 243992 2746
rect 244044 2694 244056 2746
rect 244108 2694 244120 2746
rect 244172 2694 405807 2746
rect 405859 2694 405871 2746
rect 405923 2694 405935 2746
rect 405987 2694 405999 2746
rect 406051 2694 406063 2746
rect 406115 2694 567750 2746
rect 567802 2694 567814 2746
rect 567866 2694 567878 2746
rect 567930 2694 567942 2746
rect 567994 2694 568006 2746
rect 568058 2694 648876 2746
rect 1104 2672 648876 2694
rect 18046 2592 18052 2644
rect 18104 2592 18110 2644
rect 415302 2592 415308 2644
rect 415360 2632 415366 2644
rect 419353 2635 419411 2641
rect 419353 2632 419365 2635
rect 415360 2604 419365 2632
rect 415360 2592 415366 2604
rect 419353 2601 419365 2604
rect 419399 2601 419411 2635
rect 419353 2595 419411 2601
rect 510522 2592 510528 2644
rect 510580 2632 510586 2644
rect 512089 2635 512147 2641
rect 512089 2632 512101 2635
rect 510580 2604 512101 2632
rect 510580 2592 510586 2604
rect 512089 2601 512101 2604
rect 512135 2601 512147 2635
rect 512089 2595 512147 2601
rect 602890 2592 602896 2644
rect 602948 2632 602954 2644
rect 604825 2635 604883 2641
rect 604825 2632 604837 2635
rect 602948 2604 604837 2632
rect 602948 2592 602954 2604
rect 604825 2601 604837 2604
rect 604871 2601 604883 2635
rect 604825 2595 604883 2601
rect 94593 2567 94651 2573
rect 94593 2564 94605 2567
rect 84166 2536 94605 2564
rect 21818 2456 21824 2508
rect 21876 2496 21882 2508
rect 84166 2496 84194 2536
rect 94593 2533 94605 2536
rect 94639 2533 94651 2567
rect 94593 2527 94651 2533
rect 233602 2524 233608 2576
rect 233660 2524 233666 2576
rect 326338 2524 326344 2576
rect 326396 2524 326402 2576
rect 21876 2468 84194 2496
rect 21876 2456 21882 2468
rect 115658 2456 115664 2508
rect 115716 2496 115722 2508
rect 187145 2499 187203 2505
rect 187145 2496 187157 2499
rect 115716 2468 187157 2496
rect 115716 2456 115722 2468
rect 187145 2465 187157 2468
rect 187191 2465 187203 2499
rect 187145 2459 187203 2465
rect 211338 2456 211344 2508
rect 211396 2496 211402 2508
rect 279881 2499 279939 2505
rect 279881 2496 279893 2499
rect 211396 2468 279893 2496
rect 211396 2456 211402 2468
rect 279881 2465 279893 2468
rect 279927 2465 279939 2499
rect 279881 2459 279939 2465
rect 311618 2456 311624 2508
rect 311676 2496 311682 2508
rect 402609 2499 402667 2505
rect 402609 2496 402621 2499
rect 311676 2468 402621 2496
rect 311676 2456 311682 2468
rect 402609 2465 402621 2468
rect 402655 2496 402667 2499
rect 402655 2468 402974 2496
rect 402655 2465 402667 2468
rect 402609 2459 402667 2465
rect 1578 2388 1584 2440
rect 1636 2428 1642 2440
rect 2041 2431 2099 2437
rect 2041 2428 2053 2431
rect 1636 2400 2053 2428
rect 1636 2388 1642 2400
rect 2041 2397 2053 2400
rect 2087 2397 2099 2431
rect 2041 2391 2099 2397
rect 17497 2431 17555 2437
rect 17497 2397 17509 2431
rect 17543 2428 17555 2431
rect 18046 2428 18052 2440
rect 17543 2400 18052 2428
rect 17543 2397 17555 2400
rect 17497 2391 17555 2397
rect 18046 2388 18052 2400
rect 18104 2388 18110 2440
rect 32490 2388 32496 2440
rect 32548 2428 32554 2440
rect 32953 2431 33011 2437
rect 32953 2428 32965 2431
rect 32548 2400 32965 2428
rect 32548 2388 32554 2400
rect 32953 2397 32965 2400
rect 32999 2397 33011 2431
rect 32953 2391 33011 2397
rect 47946 2388 47952 2440
rect 48004 2428 48010 2440
rect 48409 2431 48467 2437
rect 48409 2428 48421 2431
rect 48004 2400 48421 2428
rect 48004 2388 48010 2400
rect 48409 2397 48421 2400
rect 48455 2397 48467 2431
rect 48409 2391 48467 2397
rect 63862 2388 63868 2440
rect 63920 2388 63926 2440
rect 79318 2388 79324 2440
rect 79376 2388 79382 2440
rect 94314 2388 94320 2440
rect 94372 2428 94378 2440
rect 94777 2431 94835 2437
rect 94777 2428 94789 2431
rect 94372 2400 94789 2428
rect 94372 2388 94378 2400
rect 94777 2397 94789 2400
rect 94823 2397 94835 2431
rect 94777 2391 94835 2397
rect 110230 2388 110236 2440
rect 110288 2388 110294 2440
rect 125226 2388 125232 2440
rect 125284 2428 125290 2440
rect 125689 2431 125747 2437
rect 125689 2428 125701 2431
rect 125284 2400 125701 2428
rect 125284 2388 125290 2400
rect 125689 2397 125701 2400
rect 125735 2397 125747 2431
rect 125689 2391 125747 2397
rect 156598 2388 156604 2440
rect 156656 2388 156662 2440
rect 172054 2388 172060 2440
rect 172112 2388 172118 2440
rect 202506 2388 202512 2440
rect 202564 2428 202570 2440
rect 202969 2431 203027 2437
rect 202969 2428 202981 2431
rect 202564 2400 202981 2428
rect 202564 2388 202570 2400
rect 202969 2397 202981 2400
rect 203015 2397 203027 2431
rect 202969 2391 203027 2397
rect 218422 2388 218428 2440
rect 218480 2388 218486 2440
rect 248966 2388 248972 2440
rect 249024 2428 249030 2440
rect 249337 2431 249395 2437
rect 249337 2428 249349 2431
rect 249024 2400 249349 2428
rect 249024 2388 249030 2400
rect 249337 2397 249349 2400
rect 249383 2397 249395 2431
rect 249337 2391 249395 2397
rect 264790 2388 264796 2440
rect 264848 2388 264854 2440
rect 295702 2388 295708 2440
rect 295760 2388 295766 2440
rect 311158 2388 311164 2440
rect 311216 2388 311222 2440
rect 316006 2400 335354 2428
rect 17862 2360 17868 2372
rect 6886 2332 17868 2360
rect 1857 2295 1915 2301
rect 1857 2261 1869 2295
rect 1903 2292 1915 2295
rect 6886 2292 6914 2332
rect 17862 2320 17868 2332
rect 17920 2320 17926 2372
rect 20990 2320 20996 2372
rect 21048 2360 21054 2372
rect 21048 2332 35894 2360
rect 21048 2320 21054 2332
rect 1903 2264 6914 2292
rect 1903 2261 1915 2264
rect 1857 2255 1915 2261
rect 15930 2252 15936 2304
rect 15988 2292 15994 2304
rect 17313 2295 17371 2301
rect 17313 2292 17325 2295
rect 15988 2264 17325 2292
rect 15988 2252 15994 2264
rect 17313 2261 17325 2264
rect 17359 2261 17371 2295
rect 17313 2255 17371 2261
rect 31662 2252 31668 2304
rect 31720 2292 31726 2304
rect 32769 2295 32827 2301
rect 32769 2292 32781 2295
rect 31720 2264 32781 2292
rect 31720 2252 31726 2264
rect 32769 2261 32781 2264
rect 32815 2261 32827 2295
rect 35866 2292 35894 2332
rect 114462 2320 114468 2372
rect 114520 2360 114526 2372
rect 140869 2363 140927 2369
rect 140869 2360 140881 2363
rect 114520 2332 140881 2360
rect 114520 2320 114526 2332
rect 140869 2329 140881 2332
rect 140915 2329 140927 2363
rect 140869 2323 140927 2329
rect 141050 2320 141056 2372
rect 141108 2320 141114 2372
rect 186866 2320 186872 2372
rect 186924 2360 186930 2372
rect 187421 2363 187479 2369
rect 187421 2360 187433 2363
rect 186924 2332 187433 2360
rect 186924 2320 186930 2332
rect 187421 2329 187433 2332
rect 187467 2329 187479 2363
rect 187421 2323 187479 2329
rect 233786 2320 233792 2372
rect 233844 2320 233850 2372
rect 279602 2320 279608 2372
rect 279660 2360 279666 2372
rect 280157 2363 280215 2369
rect 280157 2360 280169 2363
rect 279660 2332 280169 2360
rect 279660 2320 279666 2332
rect 280157 2329 280169 2332
rect 280203 2329 280215 2363
rect 280157 2323 280215 2329
rect 307110 2320 307116 2372
rect 307168 2360 307174 2372
rect 316006 2360 316034 2400
rect 307168 2332 316034 2360
rect 307168 2320 307174 2332
rect 326522 2320 326528 2372
rect 326580 2320 326586 2372
rect 335326 2360 335354 2400
rect 342070 2388 342076 2440
rect 342128 2388 342134 2440
rect 357066 2388 357072 2440
rect 357124 2428 357130 2440
rect 357529 2431 357587 2437
rect 357529 2428 357541 2431
rect 357124 2400 357541 2428
rect 357124 2388 357130 2400
rect 357529 2397 357541 2400
rect 357575 2397 357587 2431
rect 357529 2391 357587 2397
rect 372614 2388 372620 2440
rect 372672 2428 372678 2440
rect 372985 2431 373043 2437
rect 372985 2428 372997 2431
rect 372672 2400 372997 2428
rect 372672 2388 372678 2400
rect 372985 2397 372997 2400
rect 373031 2397 373043 2431
rect 372985 2391 373043 2397
rect 387978 2388 387984 2440
rect 388036 2428 388042 2440
rect 388441 2431 388499 2437
rect 388441 2428 388453 2431
rect 388036 2400 388453 2428
rect 388036 2388 388042 2400
rect 388441 2397 388453 2400
rect 388487 2397 388499 2431
rect 402946 2428 402974 2468
rect 403897 2431 403955 2437
rect 403897 2428 403909 2431
rect 402946 2400 403909 2428
rect 388441 2391 388499 2397
rect 403897 2397 403909 2400
rect 403943 2397 403955 2431
rect 403897 2391 403955 2397
rect 418062 2388 418068 2440
rect 418120 2428 418126 2440
rect 419169 2431 419227 2437
rect 419169 2428 419181 2431
rect 418120 2400 419181 2428
rect 418120 2388 418126 2400
rect 419169 2397 419181 2400
rect 419215 2428 419227 2431
rect 419813 2431 419871 2437
rect 419813 2428 419825 2431
rect 419215 2400 419825 2428
rect 419215 2397 419227 2400
rect 419169 2391 419227 2397
rect 419813 2397 419825 2400
rect 419859 2397 419871 2431
rect 419813 2391 419871 2397
rect 434346 2388 434352 2440
rect 434404 2428 434410 2440
rect 434809 2431 434867 2437
rect 434809 2428 434821 2431
rect 434404 2400 434821 2428
rect 434404 2388 434410 2400
rect 434809 2397 434821 2400
rect 434855 2397 434867 2431
rect 434809 2391 434867 2397
rect 450262 2388 450268 2440
rect 450320 2388 450326 2440
rect 465258 2388 465264 2440
rect 465316 2428 465322 2440
rect 465721 2431 465779 2437
rect 465721 2428 465733 2431
rect 465316 2400 465733 2428
rect 465316 2388 465322 2400
rect 465721 2397 465733 2400
rect 465767 2397 465779 2431
rect 465721 2391 465779 2397
rect 480806 2388 480812 2440
rect 480864 2428 480870 2440
rect 481177 2431 481235 2437
rect 481177 2428 481189 2431
rect 480864 2400 481189 2428
rect 480864 2388 480870 2400
rect 481177 2397 481189 2400
rect 481223 2397 481235 2431
rect 481177 2391 481235 2397
rect 496170 2388 496176 2440
rect 496228 2428 496234 2440
rect 496633 2431 496691 2437
rect 496633 2428 496645 2431
rect 496228 2400 496645 2428
rect 496228 2388 496234 2400
rect 496633 2397 496645 2400
rect 496679 2397 496691 2431
rect 496633 2391 496691 2397
rect 511902 2388 511908 2440
rect 511960 2428 511966 2440
rect 512549 2431 512607 2437
rect 512549 2428 512561 2431
rect 511960 2400 512561 2428
rect 511960 2388 511966 2400
rect 512549 2397 512561 2400
rect 512595 2397 512607 2431
rect 512549 2391 512607 2397
rect 527542 2388 527548 2440
rect 527600 2388 527606 2440
rect 542998 2388 543004 2440
rect 543056 2388 543062 2440
rect 557994 2388 558000 2440
rect 558052 2428 558058 2440
rect 558457 2431 558515 2437
rect 558457 2428 558469 2431
rect 558052 2400 558469 2428
rect 558052 2388 558058 2400
rect 558457 2397 558469 2400
rect 558503 2397 558515 2431
rect 558457 2391 558515 2397
rect 573450 2388 573456 2440
rect 573508 2428 573514 2440
rect 573913 2431 573971 2437
rect 573913 2428 573925 2431
rect 573508 2400 573925 2428
rect 573508 2388 573514 2400
rect 573913 2397 573925 2400
rect 573959 2397 573971 2431
rect 573913 2391 573971 2397
rect 588906 2388 588912 2440
rect 588964 2428 588970 2440
rect 589369 2431 589427 2437
rect 589369 2428 589381 2431
rect 588964 2400 589381 2428
rect 588964 2388 588970 2400
rect 589369 2397 589381 2400
rect 589415 2397 589427 2431
rect 589369 2391 589427 2397
rect 604362 2388 604368 2440
rect 604420 2428 604426 2440
rect 604641 2431 604699 2437
rect 604641 2428 604653 2431
rect 604420 2400 604653 2428
rect 604420 2388 604426 2400
rect 604641 2397 604653 2400
rect 604687 2428 604699 2431
rect 605285 2431 605343 2437
rect 605285 2428 605297 2431
rect 604687 2400 605297 2428
rect 604687 2397 604699 2400
rect 604641 2391 604699 2397
rect 605285 2397 605297 2400
rect 605331 2397 605343 2431
rect 605285 2391 605343 2397
rect 619818 2388 619824 2440
rect 619876 2428 619882 2440
rect 620281 2431 620339 2437
rect 620281 2428 620293 2431
rect 619876 2400 620293 2428
rect 619876 2388 619882 2400
rect 620281 2397 620293 2400
rect 620327 2397 620339 2431
rect 620281 2391 620339 2397
rect 635274 2388 635280 2440
rect 635332 2428 635338 2440
rect 635737 2431 635795 2437
rect 635737 2428 635749 2431
rect 635332 2400 635749 2428
rect 635332 2388 635338 2400
rect 635737 2397 635749 2400
rect 635783 2397 635795 2431
rect 635737 2391 635795 2397
rect 335326 2332 364334 2360
rect 48225 2295 48283 2301
rect 48225 2292 48237 2295
rect 35866 2264 48237 2292
rect 32769 2255 32827 2261
rect 48225 2261 48237 2264
rect 48271 2261 48283 2295
rect 48225 2255 48283 2261
rect 62022 2252 62028 2304
rect 62080 2292 62086 2304
rect 63681 2295 63739 2301
rect 63681 2292 63693 2295
rect 62080 2264 63693 2292
rect 62080 2252 62086 2264
rect 63681 2261 63693 2264
rect 63727 2261 63739 2295
rect 63681 2255 63739 2261
rect 77202 2252 77208 2304
rect 77260 2292 77266 2304
rect 79137 2295 79195 2301
rect 79137 2292 79149 2295
rect 77260 2264 79149 2292
rect 77260 2252 77266 2264
rect 79137 2261 79149 2264
rect 79183 2261 79195 2295
rect 79137 2255 79195 2261
rect 107562 2252 107568 2304
rect 107620 2292 107626 2304
rect 110049 2295 110107 2301
rect 110049 2292 110061 2295
rect 107620 2264 110061 2292
rect 107620 2252 107626 2264
rect 110049 2261 110061 2264
rect 110095 2261 110107 2295
rect 110049 2255 110107 2261
rect 122650 2252 122656 2304
rect 122708 2292 122714 2304
rect 125505 2295 125563 2301
rect 125505 2292 125517 2295
rect 122708 2264 125517 2292
rect 122708 2252 122714 2264
rect 125505 2261 125517 2264
rect 125551 2261 125563 2295
rect 125505 2255 125563 2261
rect 156414 2252 156420 2304
rect 156472 2252 156478 2304
rect 169662 2252 169668 2304
rect 169720 2292 169726 2304
rect 171873 2295 171931 2301
rect 171873 2292 171885 2295
rect 169720 2264 171885 2292
rect 169720 2252 169726 2264
rect 171873 2261 171885 2264
rect 171919 2261 171931 2295
rect 171873 2255 171931 2261
rect 199470 2252 199476 2304
rect 199528 2292 199534 2304
rect 202785 2295 202843 2301
rect 202785 2292 202797 2295
rect 199528 2264 202797 2292
rect 199528 2252 199534 2264
rect 202785 2261 202797 2264
rect 202831 2261 202843 2295
rect 202785 2255 202843 2261
rect 218238 2252 218244 2304
rect 218296 2252 218302 2304
rect 249150 2252 249156 2304
rect 249208 2252 249214 2304
rect 264606 2252 264612 2304
rect 264664 2252 264670 2304
rect 293954 2252 293960 2304
rect 294012 2292 294018 2304
rect 295521 2295 295579 2301
rect 295521 2292 295533 2295
rect 294012 2264 295533 2292
rect 294012 2252 294018 2264
rect 295521 2261 295533 2264
rect 295567 2261 295579 2295
rect 295521 2255 295579 2261
rect 309134 2252 309140 2304
rect 309192 2292 309198 2304
rect 310977 2295 311035 2301
rect 310977 2292 310989 2295
rect 309192 2264 310989 2292
rect 309192 2252 309198 2264
rect 310977 2261 310989 2264
rect 311023 2261 311035 2295
rect 310977 2255 311035 2261
rect 339494 2252 339500 2304
rect 339552 2292 339558 2304
rect 341889 2295 341947 2301
rect 341889 2292 341901 2295
rect 339552 2264 341901 2292
rect 339552 2252 339558 2264
rect 341889 2261 341901 2264
rect 341935 2261 341947 2295
rect 341889 2255 341947 2261
rect 357342 2252 357348 2304
rect 357400 2252 357406 2304
rect 364306 2292 364334 2332
rect 403342 2320 403348 2372
rect 403400 2360 403406 2372
rect 403400 2332 451274 2360
rect 403400 2320 403406 2332
rect 372801 2295 372859 2301
rect 372801 2292 372813 2295
rect 364306 2264 372813 2292
rect 372801 2261 372813 2264
rect 372847 2261 372859 2295
rect 372801 2255 372859 2261
rect 386414 2252 386420 2304
rect 386472 2292 386478 2304
rect 388257 2295 388315 2301
rect 388257 2292 388269 2295
rect 386472 2264 388269 2292
rect 386472 2252 386478 2264
rect 388257 2261 388269 2264
rect 388303 2261 388315 2295
rect 388257 2255 388315 2261
rect 402698 2252 402704 2304
rect 402756 2292 402762 2304
rect 403713 2295 403771 2301
rect 403713 2292 403725 2295
rect 402756 2264 403725 2292
rect 402756 2252 402762 2264
rect 403713 2261 403725 2264
rect 403759 2261 403771 2295
rect 403713 2255 403771 2261
rect 432782 2252 432788 2304
rect 432840 2292 432846 2304
rect 434625 2295 434683 2301
rect 434625 2292 434637 2295
rect 432840 2264 434637 2292
rect 432840 2252 432846 2264
rect 434625 2261 434637 2264
rect 434671 2261 434683 2295
rect 434625 2255 434683 2261
rect 450078 2252 450084 2304
rect 450136 2252 450142 2304
rect 451246 2292 451274 2332
rect 499850 2320 499856 2372
rect 499908 2360 499914 2372
rect 499908 2332 547874 2360
rect 499908 2320 499914 2332
rect 465537 2295 465595 2301
rect 465537 2292 465549 2295
rect 451246 2264 465549 2292
rect 465537 2261 465549 2264
rect 465583 2261 465595 2295
rect 465537 2255 465595 2261
rect 480990 2252 480996 2304
rect 481048 2252 481054 2304
rect 496446 2252 496452 2304
rect 496504 2252 496510 2304
rect 527358 2252 527364 2304
rect 527416 2252 527422 2304
rect 542814 2252 542820 2304
rect 542872 2252 542878 2304
rect 547846 2292 547874 2332
rect 558273 2295 558331 2301
rect 558273 2292 558285 2295
rect 547846 2264 558285 2292
rect 558273 2261 558285 2264
rect 558319 2261 558331 2295
rect 558273 2255 558331 2261
rect 573726 2252 573732 2304
rect 573784 2252 573790 2304
rect 589182 2252 589188 2304
rect 589240 2252 589246 2304
rect 618254 2252 618260 2304
rect 618312 2292 618318 2304
rect 620097 2295 620155 2301
rect 620097 2292 620109 2295
rect 618312 2264 620109 2292
rect 618312 2252 618318 2264
rect 620097 2261 620109 2264
rect 620143 2261 620155 2295
rect 620097 2255 620155 2261
rect 633434 2252 633440 2304
rect 633492 2292 633498 2304
rect 635553 2295 635611 2301
rect 635553 2292 635565 2295
rect 633492 2264 635565 2292
rect 633492 2252 633498 2264
rect 635553 2261 635565 2264
rect 635599 2261 635611 2295
rect 635553 2255 635611 2261
rect 1104 2202 648876 2224
rect 1104 2150 82581 2202
rect 82633 2150 82645 2202
rect 82697 2150 82709 2202
rect 82761 2150 82773 2202
rect 82825 2150 82837 2202
rect 82889 2150 244524 2202
rect 244576 2150 244588 2202
rect 244640 2150 244652 2202
rect 244704 2150 244716 2202
rect 244768 2150 244780 2202
rect 244832 2150 406467 2202
rect 406519 2150 406531 2202
rect 406583 2150 406595 2202
rect 406647 2150 406659 2202
rect 406711 2150 406723 2202
rect 406775 2150 568410 2202
rect 568462 2150 568474 2202
rect 568526 2150 568538 2202
rect 568590 2150 568602 2202
rect 568654 2150 568666 2202
rect 568718 2150 648876 2202
rect 1104 2128 648876 2150
rect 74 796 130 800
rect 1578 796 1584 808
rect 74 768 1584 796
rect 74 0 130 768
rect 1578 756 1584 768
rect 1636 756 1642 808
rect 15374 796 15430 800
rect 15930 796 15936 808
rect 15374 768 15936 796
rect 15374 0 15430 768
rect 15930 756 15936 768
rect 15988 756 15994 808
rect 30674 796 30730 800
rect 31662 796 31668 808
rect 30674 768 31668 796
rect 30674 0 30730 768
rect 31662 756 31668 768
rect 31720 756 31726 808
rect 45974 796 46030 800
rect 47946 796 47952 808
rect 45974 768 47952 796
rect 45974 0 46030 768
rect 47946 756 47952 768
rect 48004 756 48010 808
rect 61274 796 61330 800
rect 62022 796 62028 808
rect 61274 768 62028 796
rect 61274 0 61330 768
rect 62022 756 62028 768
rect 62080 756 62086 808
rect 76574 796 76630 800
rect 77202 796 77208 808
rect 76574 768 77208 796
rect 76574 0 76630 768
rect 77202 756 77208 768
rect 77260 756 77266 808
rect 91874 796 91930 800
rect 94314 796 94320 808
rect 91874 768 94320 796
rect 91874 0 91930 768
rect 94314 756 94320 768
rect 94372 756 94378 808
rect 107174 796 107230 800
rect 107562 796 107568 808
rect 107174 768 107568 796
rect 107174 0 107230 768
rect 107562 756 107568 768
rect 107620 756 107626 808
rect 122474 796 122530 800
rect 122650 796 122656 808
rect 122474 768 122656 796
rect 122474 0 122530 768
rect 122650 756 122656 768
rect 122708 756 122714 808
rect 137774 796 137830 800
rect 141050 796 141056 808
rect 137774 768 141056 796
rect 137774 0 137830 768
rect 141050 756 141056 768
rect 141108 756 141114 808
rect 153074 796 153130 800
rect 156414 796 156420 808
rect 153074 768 156420 796
rect 153074 0 153130 768
rect 156414 756 156420 768
rect 156472 756 156478 808
rect 168374 796 168430 800
rect 169662 796 169668 808
rect 168374 768 169668 796
rect 168374 0 168430 768
rect 169662 756 169668 768
rect 169720 756 169726 808
rect 183674 796 183730 800
rect 186866 796 186872 808
rect 183674 768 186872 796
rect 183674 0 183730 768
rect 186866 756 186872 768
rect 186924 756 186930 808
rect 198974 796 199030 800
rect 199470 796 199476 808
rect 198974 768 199476 796
rect 198974 0 199030 768
rect 199470 756 199476 768
rect 199528 756 199534 808
rect 214274 796 214330 800
rect 218238 796 218244 808
rect 214274 768 218244 796
rect 214274 0 214330 768
rect 218238 756 218244 768
rect 218296 756 218302 808
rect 229574 796 229630 800
rect 233786 796 233792 808
rect 229574 768 233792 796
rect 229574 0 229630 768
rect 233786 756 233792 768
rect 233844 756 233850 808
rect 244874 796 244930 800
rect 249150 796 249156 808
rect 244874 768 249156 796
rect 244874 0 244930 768
rect 249150 756 249156 768
rect 249208 756 249214 808
rect 260174 796 260230 800
rect 264606 796 264612 808
rect 260174 768 264612 796
rect 260174 0 260230 768
rect 264606 756 264612 768
rect 264664 756 264670 808
rect 275474 796 275530 800
rect 279602 796 279608 808
rect 275474 768 279608 796
rect 275474 0 275530 768
rect 279602 756 279608 768
rect 279660 756 279666 808
rect 290774 796 290830 800
rect 293954 796 293960 808
rect 290774 768 293960 796
rect 290774 0 290830 768
rect 293954 756 293960 768
rect 294012 756 294018 808
rect 306074 48 306130 800
rect 321374 796 321430 800
rect 326522 796 326528 808
rect 321374 768 326528 796
rect 309134 48 309140 60
rect 306074 20 309140 48
rect 306074 0 306130 20
rect 309134 8 309140 20
rect 309192 8 309198 60
rect 321374 0 321430 768
rect 326522 756 326528 768
rect 326580 756 326586 808
rect 336674 796 336730 800
rect 339494 796 339500 808
rect 336674 768 339500 796
rect 336674 0 336730 768
rect 339494 756 339500 768
rect 339552 756 339558 808
rect 351974 796 352030 800
rect 357342 796 357348 808
rect 351974 768 357348 796
rect 351974 0 352030 768
rect 357342 756 357348 768
rect 357400 756 357406 808
rect 367274 796 367330 800
rect 372614 796 372620 808
rect 367274 768 372620 796
rect 367274 0 367330 768
rect 372614 756 372620 768
rect 372672 756 372678 808
rect 382574 48 382630 800
rect 397874 796 397930 800
rect 402698 796 402704 808
rect 397874 768 402704 796
rect 386414 48 386420 60
rect 382574 20 386420 48
rect 382574 0 382630 20
rect 386414 8 386420 20
rect 386472 8 386478 60
rect 397874 0 397930 768
rect 402698 756 402704 768
rect 402756 756 402762 808
rect 413174 796 413230 800
rect 418062 796 418068 808
rect 413174 768 418068 796
rect 413174 0 413230 768
rect 418062 756 418068 768
rect 418120 756 418126 808
rect 428474 796 428530 800
rect 432782 796 432788 808
rect 428474 768 432788 796
rect 428474 0 428530 768
rect 432782 756 432788 768
rect 432840 756 432846 808
rect 443774 796 443830 800
rect 450078 796 450084 808
rect 443774 768 450084 796
rect 443774 0 443830 768
rect 450078 756 450084 768
rect 450136 756 450142 808
rect 459074 48 459130 800
rect 474374 796 474430 800
rect 480990 796 480996 808
rect 474374 768 480996 796
rect 465258 48 465264 60
rect 459074 20 465264 48
rect 459074 0 459130 20
rect 465258 8 465264 20
rect 465316 8 465322 60
rect 474374 0 474430 768
rect 480990 756 480996 768
rect 481048 756 481054 808
rect 489674 48 489730 800
rect 504974 796 505030 800
rect 511902 796 511908 808
rect 504974 768 511908 796
rect 496446 48 496452 60
rect 489674 20 496452 48
rect 489674 0 489730 20
rect 496446 8 496452 20
rect 496504 8 496510 60
rect 504974 0 505030 768
rect 511902 756 511908 768
rect 511960 756 511966 808
rect 520274 796 520330 800
rect 527358 796 527364 808
rect 520274 768 527364 796
rect 520274 0 520330 768
rect 527358 756 527364 768
rect 527416 756 527422 808
rect 535574 48 535630 800
rect 550874 796 550930 800
rect 557994 796 558000 808
rect 550874 768 558000 796
rect 542814 48 542820 60
rect 535574 20 542820 48
rect 535574 0 535630 20
rect 542814 8 542820 20
rect 542872 8 542878 60
rect 550874 0 550930 768
rect 557994 756 558000 768
rect 558052 756 558058 808
rect 566174 48 566230 800
rect 581474 796 581530 800
rect 589182 796 589188 808
rect 581474 768 589188 796
rect 573726 48 573732 60
rect 566174 20 573732 48
rect 566174 0 566230 20
rect 573726 8 573732 20
rect 573784 8 573790 60
rect 581474 0 581530 768
rect 589182 756 589188 768
rect 589240 756 589246 808
rect 596774 796 596830 800
rect 604362 796 604368 808
rect 596774 768 604368 796
rect 596774 0 596830 768
rect 604362 756 604368 768
rect 604420 756 604426 808
rect 612074 48 612130 800
rect 627374 796 627430 800
rect 633434 796 633440 808
rect 627374 768 633440 796
rect 618254 48 618260 60
rect 612074 20 618260 48
rect 612074 0 612130 20
rect 618254 8 618260 20
rect 618312 8 618318 60
rect 627374 0 627430 768
rect 633434 756 633440 768
rect 633492 756 633498 808
<< via1 >>
rect 19708 9188 19760 9240
rect 20168 9188 20220 9240
rect 20996 9188 21048 9240
rect 21272 9188 21324 9240
rect 22928 9188 22980 9240
rect 23204 9188 23256 9240
rect 23756 9188 23808 9240
rect 20628 8848 20680 8900
rect 21824 8916 21876 8968
rect 22008 8916 22060 8968
rect 21916 8848 21968 8900
rect 23388 9120 23440 9172
rect 24308 9188 24360 9240
rect 24584 9188 24636 9240
rect 25136 9188 25188 9240
rect 23296 8916 23348 8968
rect 24768 9120 24820 9172
rect 25688 9188 25740 9240
rect 25964 9188 26016 9240
rect 26148 9188 26200 9240
rect 26700 9188 26752 9240
rect 27252 9188 27304 9240
rect 27528 9188 27580 9240
rect 27804 9188 27856 9240
rect 28080 9188 28132 9240
rect 28356 9188 28408 9240
rect 28908 9188 28960 9240
rect 29184 9188 29236 9240
rect 29460 9188 29512 9240
rect 29736 9188 29788 9240
rect 30012 9188 30064 9240
rect 30104 9120 30156 9172
rect 30472 9120 30524 9172
rect 30840 9188 30892 9240
rect 31116 9188 31168 9240
rect 31484 9188 31536 9240
rect 118976 9120 119028 9172
rect 30288 9052 30340 9104
rect 110144 9052 110196 9104
rect 108488 8984 108540 9036
rect 30380 8916 30432 8968
rect 107292 8916 107344 8968
rect 30472 8848 30524 8900
rect 104624 8848 104676 8900
rect 78036 8780 78088 8832
rect 29736 8712 29788 8764
rect 74080 8712 74132 8764
rect 30288 8644 30340 8696
rect 30380 8644 30432 8696
rect 62580 8644 62632 8696
rect 26148 8508 26200 8560
rect 30196 8508 30248 8560
rect 35256 8576 35308 8628
rect 30656 8508 30708 8560
rect 36820 8576 36872 8628
rect 25688 8440 25740 8492
rect 32680 8440 32732 8492
rect 27252 8372 27304 8424
rect 123852 8372 123904 8424
rect 30656 8236 30708 8288
rect 57336 8236 57388 8288
rect 151176 8236 151228 8288
rect 74908 8168 74960 8220
rect 168196 8168 168248 8220
rect 22928 8100 22980 8152
rect 65892 8100 65944 8152
rect 72792 8100 72844 8152
rect 166448 8100 166500 8152
rect 28080 8032 28132 8084
rect 76104 8032 76156 8084
rect 24768 7964 24820 8016
rect 79968 7964 80020 8016
rect 31116 7896 31168 7948
rect 56600 7896 56652 7948
rect 76932 7896 76984 7948
rect 170128 7896 170180 7948
rect 33508 7828 33560 7880
rect 125324 7828 125376 7880
rect 27804 7760 27856 7812
rect 60924 7760 60976 7812
rect 107844 7760 107896 7812
rect 200120 7760 200172 7812
rect 31484 7692 31536 7744
rect 71964 7692 72016 7744
rect 105820 7692 105872 7744
rect 197912 7692 197964 7744
rect 82581 7590 82633 7642
rect 82645 7590 82697 7642
rect 82709 7590 82761 7642
rect 82773 7590 82825 7642
rect 82837 7590 82889 7642
rect 244524 7590 244576 7642
rect 244588 7590 244640 7642
rect 244652 7590 244704 7642
rect 244716 7590 244768 7642
rect 244780 7590 244832 7642
rect 406467 7590 406519 7642
rect 406531 7590 406583 7642
rect 406595 7590 406647 7642
rect 406659 7590 406711 7642
rect 406723 7590 406775 7642
rect 568410 7590 568462 7642
rect 568474 7590 568526 7642
rect 568538 7590 568590 7642
rect 568602 7590 568654 7642
rect 568666 7590 568718 7642
rect 25136 7488 25188 7540
rect 25964 7420 26016 7472
rect 32680 7395 32732 7404
rect 32680 7361 32689 7395
rect 32689 7361 32723 7395
rect 32723 7361 32732 7395
rect 32680 7352 32732 7361
rect 33508 7395 33560 7404
rect 33508 7361 33517 7395
rect 33517 7361 33551 7395
rect 33551 7361 33560 7395
rect 33508 7352 33560 7361
rect 35256 7395 35308 7404
rect 35256 7361 35265 7395
rect 35265 7361 35299 7395
rect 35299 7361 35308 7395
rect 35256 7352 35308 7361
rect 36820 7395 36872 7404
rect 36820 7361 36829 7395
rect 36829 7361 36863 7395
rect 36863 7361 36872 7395
rect 36820 7352 36872 7361
rect 56600 7395 56652 7404
rect 56600 7361 56609 7395
rect 56609 7361 56643 7395
rect 56643 7361 56652 7395
rect 56600 7352 56652 7361
rect 57336 7395 57388 7404
rect 57336 7361 57345 7395
rect 57345 7361 57379 7395
rect 57379 7361 57388 7395
rect 57336 7352 57388 7361
rect 35532 7327 35584 7336
rect 35532 7293 35541 7327
rect 35541 7293 35575 7327
rect 35575 7293 35584 7327
rect 35532 7284 35584 7293
rect 37740 7327 37792 7336
rect 37740 7293 37749 7327
rect 37749 7293 37783 7327
rect 37783 7293 37792 7327
rect 37740 7284 37792 7293
rect 29460 7216 29512 7268
rect 60924 7395 60976 7404
rect 60924 7361 60933 7395
rect 60933 7361 60967 7395
rect 60967 7361 60976 7395
rect 60924 7352 60976 7361
rect 62580 7352 62632 7404
rect 63040 7352 63092 7404
rect 64788 7395 64840 7404
rect 64788 7361 64797 7395
rect 64797 7361 64831 7395
rect 64831 7361 64840 7395
rect 64788 7352 64840 7361
rect 65892 7395 65944 7404
rect 65892 7361 65901 7395
rect 65901 7361 65935 7395
rect 65935 7361 65944 7395
rect 65892 7352 65944 7361
rect 71964 7395 72016 7404
rect 71964 7361 71973 7395
rect 71973 7361 72007 7395
rect 72007 7361 72016 7395
rect 71964 7352 72016 7361
rect 72792 7395 72844 7404
rect 72792 7361 72801 7395
rect 72801 7361 72835 7395
rect 72835 7361 72844 7395
rect 72792 7352 72844 7361
rect 74080 7395 74132 7404
rect 74080 7361 74089 7395
rect 74089 7361 74123 7395
rect 74123 7361 74132 7395
rect 74080 7352 74132 7361
rect 74908 7395 74960 7404
rect 74908 7361 74917 7395
rect 74917 7361 74951 7395
rect 74951 7361 74960 7395
rect 74908 7352 74960 7361
rect 76104 7395 76156 7404
rect 76104 7361 76113 7395
rect 76113 7361 76147 7395
rect 76147 7361 76156 7395
rect 76104 7352 76156 7361
rect 76932 7395 76984 7404
rect 76932 7361 76941 7395
rect 76941 7361 76975 7395
rect 76975 7361 76984 7395
rect 76932 7352 76984 7361
rect 78036 7395 78088 7404
rect 78036 7361 78045 7395
rect 78045 7361 78079 7395
rect 78079 7361 78088 7395
rect 78036 7352 78088 7361
rect 79600 7352 79652 7404
rect 79968 7352 80020 7404
rect 104624 7395 104676 7404
rect 104624 7361 104633 7395
rect 104633 7361 104667 7395
rect 104667 7361 104676 7395
rect 104624 7352 104676 7361
rect 105820 7395 105872 7404
rect 105820 7361 105829 7395
rect 105829 7361 105863 7395
rect 105863 7361 105872 7395
rect 105820 7352 105872 7361
rect 107292 7395 107344 7404
rect 107292 7361 107301 7395
rect 107301 7361 107335 7395
rect 107335 7361 107344 7395
rect 107292 7352 107344 7361
rect 107844 7463 107896 7472
rect 107844 7429 107853 7463
rect 107853 7429 107887 7463
rect 107887 7429 107896 7463
rect 107844 7420 107896 7429
rect 123208 7488 123260 7540
rect 110144 7395 110196 7404
rect 110144 7361 110153 7395
rect 110153 7361 110187 7395
rect 110187 7361 110196 7395
rect 110144 7352 110196 7361
rect 59636 7327 59688 7336
rect 59636 7293 59645 7327
rect 59645 7293 59679 7327
rect 59679 7293 59688 7327
rect 59636 7284 59688 7293
rect 63776 7327 63828 7336
rect 63776 7293 63785 7327
rect 63785 7293 63819 7327
rect 63819 7293 63828 7327
rect 63776 7284 63828 7293
rect 65064 7327 65116 7336
rect 65064 7293 65073 7327
rect 65073 7293 65107 7327
rect 65107 7293 65116 7327
rect 65064 7284 65116 7293
rect 66720 7327 66772 7336
rect 66720 7293 66729 7327
rect 66729 7293 66763 7327
rect 66763 7293 66772 7327
rect 66720 7284 66772 7293
rect 79324 7327 79376 7336
rect 79324 7293 79333 7327
rect 79333 7293 79367 7327
rect 79367 7293 79376 7327
rect 79324 7284 79376 7293
rect 80612 7327 80664 7336
rect 80612 7293 80621 7327
rect 80621 7293 80655 7327
rect 80655 7293 80664 7327
rect 80612 7284 80664 7293
rect 111340 7327 111392 7336
rect 111340 7293 111349 7327
rect 111349 7293 111383 7327
rect 111383 7293 111392 7327
rect 111340 7284 111392 7293
rect 117964 7352 118016 7404
rect 119344 7352 119396 7404
rect 118976 7284 119028 7336
rect 121460 7395 121512 7404
rect 121460 7361 121469 7395
rect 121469 7361 121503 7395
rect 121503 7361 121512 7395
rect 121460 7352 121512 7361
rect 121828 7395 121880 7404
rect 121828 7361 121837 7395
rect 121837 7361 121871 7395
rect 121871 7361 121880 7395
rect 121828 7352 121880 7361
rect 122840 7395 122892 7404
rect 122840 7361 122849 7395
rect 122849 7361 122883 7395
rect 122883 7361 122892 7395
rect 122840 7352 122892 7361
rect 123208 7395 123260 7404
rect 123208 7361 123217 7395
rect 123217 7361 123251 7395
rect 123251 7361 123260 7395
rect 123208 7352 123260 7361
rect 123852 7395 123904 7404
rect 123852 7361 123861 7395
rect 123861 7361 123895 7395
rect 123895 7361 123904 7395
rect 123852 7352 123904 7361
rect 125324 7395 125376 7404
rect 125324 7361 125333 7395
rect 125333 7361 125367 7395
rect 125367 7361 125376 7395
rect 125324 7352 125376 7361
rect 151176 7395 151228 7404
rect 151176 7361 151185 7395
rect 151185 7361 151219 7395
rect 151219 7361 151228 7395
rect 151176 7352 151228 7361
rect 152740 7352 152792 7404
rect 125508 7284 125560 7336
rect 126520 7327 126572 7336
rect 126520 7293 126529 7327
rect 126529 7293 126563 7327
rect 126563 7293 126572 7327
rect 126520 7284 126572 7293
rect 151728 7327 151780 7336
rect 151728 7293 151737 7327
rect 151737 7293 151771 7327
rect 151771 7293 151780 7327
rect 151728 7284 151780 7293
rect 154488 7284 154540 7336
rect 166448 7395 166500 7404
rect 166448 7361 166457 7395
rect 166457 7361 166491 7395
rect 166491 7361 166500 7395
rect 166448 7352 166500 7361
rect 168196 7395 168248 7404
rect 168196 7361 168205 7395
rect 168205 7361 168239 7395
rect 168239 7361 168248 7395
rect 168196 7352 168248 7361
rect 170128 7395 170180 7404
rect 170128 7361 170137 7395
rect 170137 7361 170171 7395
rect 170171 7361 170180 7395
rect 170128 7352 170180 7361
rect 197912 7395 197964 7404
rect 197912 7361 197921 7395
rect 197921 7361 197955 7395
rect 197955 7361 197964 7395
rect 197912 7352 197964 7361
rect 200120 7395 200172 7404
rect 200120 7361 200129 7395
rect 200129 7361 200163 7395
rect 200163 7361 200172 7395
rect 200120 7352 200172 7361
rect 217876 7352 217928 7404
rect 220452 7352 220504 7404
rect 244372 7395 244424 7404
rect 244372 7361 244381 7395
rect 244381 7361 244415 7395
rect 244415 7361 244424 7395
rect 244372 7352 244424 7361
rect 157340 7284 157392 7336
rect 154580 7216 154632 7268
rect 169484 7327 169536 7336
rect 169484 7293 169493 7327
rect 169493 7293 169527 7327
rect 169527 7293 169536 7327
rect 169484 7284 169536 7293
rect 170680 7327 170732 7336
rect 170680 7293 170689 7327
rect 170689 7293 170723 7327
rect 170723 7293 170732 7327
rect 170680 7284 170732 7293
rect 199108 7327 199160 7336
rect 199108 7293 199117 7327
rect 199117 7293 199151 7327
rect 199151 7293 199160 7327
rect 199108 7284 199160 7293
rect 201316 7327 201368 7336
rect 201316 7293 201325 7327
rect 201325 7293 201359 7327
rect 201359 7293 201368 7327
rect 201316 7284 201368 7293
rect 214564 7327 214616 7336
rect 214564 7293 214573 7327
rect 214573 7293 214607 7327
rect 214607 7293 214616 7327
rect 214564 7284 214616 7293
rect 214748 7284 214800 7336
rect 245476 7327 245528 7336
rect 245476 7293 245485 7327
rect 245485 7293 245519 7327
rect 245519 7293 245528 7327
rect 245476 7284 245528 7293
rect 260748 7327 260800 7336
rect 260748 7293 260757 7327
rect 260757 7293 260791 7327
rect 260791 7293 260800 7327
rect 260748 7284 260800 7293
rect 152740 7191 152792 7200
rect 152740 7157 152749 7191
rect 152749 7157 152783 7191
rect 152783 7157 152792 7191
rect 152740 7148 152792 7157
rect 217876 7191 217928 7200
rect 217876 7157 217885 7191
rect 217885 7157 217919 7191
rect 217919 7157 217928 7191
rect 217876 7148 217928 7157
rect 220452 7191 220504 7200
rect 220452 7157 220461 7191
rect 220461 7157 220495 7191
rect 220495 7157 220504 7191
rect 220452 7148 220504 7157
rect 81921 7046 81973 7098
rect 81985 7046 82037 7098
rect 82049 7046 82101 7098
rect 82113 7046 82165 7098
rect 82177 7046 82229 7098
rect 243864 7046 243916 7098
rect 243928 7046 243980 7098
rect 243992 7046 244044 7098
rect 244056 7046 244108 7098
rect 244120 7046 244172 7098
rect 405807 7046 405859 7098
rect 405871 7046 405923 7098
rect 405935 7046 405987 7098
rect 405999 7046 406051 7098
rect 406063 7046 406115 7098
rect 567750 7046 567802 7098
rect 567814 7046 567866 7098
rect 567878 7046 567930 7098
rect 567942 7046 567994 7098
rect 568006 7046 568058 7098
rect 24584 6944 24636 6996
rect 35256 6876 35308 6928
rect 59636 6944 59688 6996
rect 152740 6944 152792 6996
rect 64788 6876 64840 6928
rect 107292 6876 107344 6928
rect 118976 6919 119028 6928
rect 118976 6885 118985 6919
rect 118985 6885 119019 6919
rect 119019 6885 119028 6919
rect 118976 6876 119028 6885
rect 123208 6876 123260 6928
rect 151176 6876 151228 6928
rect 151728 6876 151780 6928
rect 154580 6919 154632 6928
rect 154580 6885 154589 6919
rect 154589 6885 154623 6919
rect 154623 6885 154632 6919
rect 154580 6876 154632 6885
rect 166448 6944 166500 6996
rect 170128 6944 170180 6996
rect 170220 6944 170272 6996
rect 172336 6944 172388 6996
rect 215300 6944 215352 6996
rect 218796 6944 218848 6996
rect 215852 6876 215904 6928
rect 216036 6876 216088 6928
rect 244372 6876 244424 6928
rect 17868 6808 17920 6860
rect 19708 6808 19760 6860
rect 26700 6808 26752 6860
rect 18052 6740 18104 6792
rect 20168 6740 20220 6792
rect 63040 6740 63092 6792
rect 79600 6740 79652 6792
rect 81532 6783 81584 6792
rect 81532 6749 81541 6783
rect 81541 6749 81575 6783
rect 81575 6749 81584 6783
rect 81532 6740 81584 6749
rect 30012 6672 30064 6724
rect 82452 6672 82504 6724
rect 108488 6783 108540 6792
rect 108488 6749 108497 6783
rect 108497 6749 108531 6783
rect 108531 6749 108540 6783
rect 108488 6740 108540 6749
rect 116124 6715 116176 6724
rect 116124 6681 116133 6715
rect 116133 6681 116167 6715
rect 116167 6681 116176 6715
rect 116124 6672 116176 6681
rect 117044 6740 117096 6792
rect 120448 6740 120500 6792
rect 121460 6740 121512 6792
rect 124036 6783 124088 6792
rect 124036 6749 124045 6783
rect 124045 6749 124079 6783
rect 124079 6749 124088 6783
rect 124036 6740 124088 6749
rect 117412 6647 117464 6656
rect 117412 6613 117421 6647
rect 117421 6613 117455 6647
rect 117455 6613 117464 6647
rect 117412 6604 117464 6613
rect 117964 6647 118016 6656
rect 117964 6613 117973 6647
rect 117973 6613 118007 6647
rect 118007 6613 118016 6647
rect 117964 6604 118016 6613
rect 120816 6715 120868 6724
rect 120816 6681 120825 6715
rect 120825 6681 120859 6715
rect 120859 6681 120868 6715
rect 120816 6672 120868 6681
rect 124680 6715 124732 6724
rect 124680 6681 124689 6715
rect 124689 6681 124723 6715
rect 124723 6681 124732 6715
rect 124680 6672 124732 6681
rect 155776 6740 155828 6792
rect 155776 6647 155828 6656
rect 155776 6613 155785 6647
rect 155785 6613 155819 6647
rect 155819 6613 155828 6647
rect 155776 6604 155828 6613
rect 156972 6715 157024 6724
rect 156972 6681 156981 6715
rect 156981 6681 157015 6715
rect 157015 6681 157024 6715
rect 156972 6672 157024 6681
rect 170220 6808 170272 6860
rect 170680 6808 170732 6860
rect 215760 6808 215812 6860
rect 216220 6808 216272 6860
rect 262956 6808 263008 6860
rect 171048 6740 171100 6792
rect 173072 6740 173124 6792
rect 215300 6740 215352 6792
rect 171048 6647 171100 6656
rect 171048 6613 171057 6647
rect 171057 6613 171091 6647
rect 171091 6613 171100 6647
rect 171048 6604 171100 6613
rect 172244 6715 172296 6724
rect 172244 6681 172253 6715
rect 172253 6681 172287 6715
rect 172287 6681 172296 6715
rect 172244 6672 172296 6681
rect 172336 6672 172388 6724
rect 214748 6672 214800 6724
rect 190552 6604 190604 6656
rect 190644 6604 190696 6656
rect 213276 6604 213328 6656
rect 213368 6604 213420 6656
rect 216588 6715 216640 6724
rect 216588 6681 216597 6715
rect 216597 6681 216631 6715
rect 216631 6681 216640 6715
rect 216588 6672 216640 6681
rect 217508 6715 217560 6724
rect 217508 6681 217517 6715
rect 217517 6681 217551 6715
rect 217551 6681 217560 6715
rect 217508 6672 217560 6681
rect 218796 6740 218848 6792
rect 246764 6783 246816 6792
rect 246764 6749 246773 6783
rect 246773 6749 246807 6783
rect 246807 6749 246816 6783
rect 246764 6740 246816 6749
rect 261760 6740 261812 6792
rect 246120 6647 246172 6656
rect 246120 6613 246129 6647
rect 246129 6613 246163 6647
rect 246163 6613 246172 6647
rect 246120 6604 246172 6613
rect 247316 6715 247368 6724
rect 247316 6681 247325 6715
rect 247325 6681 247359 6715
rect 247359 6681 247368 6715
rect 247316 6672 247368 6681
rect 262588 6715 262640 6724
rect 262588 6681 262597 6715
rect 262597 6681 262631 6715
rect 262631 6681 262640 6715
rect 262588 6672 262640 6681
rect 310888 6604 310940 6656
rect 82581 6502 82633 6554
rect 82645 6502 82697 6554
rect 82709 6502 82761 6554
rect 82773 6502 82825 6554
rect 82837 6502 82889 6554
rect 244524 6502 244576 6554
rect 244588 6502 244640 6554
rect 244652 6502 244704 6554
rect 244716 6502 244768 6554
rect 244780 6502 244832 6554
rect 406467 6502 406519 6554
rect 406531 6502 406583 6554
rect 406595 6502 406647 6554
rect 406659 6502 406711 6554
rect 406723 6502 406775 6554
rect 568410 6502 568462 6554
rect 568474 6502 568526 6554
rect 568538 6502 568590 6554
rect 568602 6502 568654 6554
rect 568666 6502 568718 6554
rect 63776 6400 63828 6452
rect 155776 6400 155828 6452
rect 157340 6400 157392 6452
rect 167184 6400 167236 6452
rect 169484 6400 169536 6452
rect 173072 6400 173124 6452
rect 173164 6400 173216 6452
rect 190644 6400 190696 6452
rect 190736 6400 190788 6452
rect 200580 6400 200632 6452
rect 23756 6332 23808 6384
rect 27528 6264 27580 6316
rect 123852 6332 123904 6384
rect 124036 6332 124088 6384
rect 214564 6400 214616 6452
rect 120816 6264 120868 6316
rect 122564 6307 122616 6316
rect 122564 6273 122573 6307
rect 122573 6273 122607 6307
rect 122607 6273 122616 6307
rect 122564 6264 122616 6273
rect 112352 6239 112404 6248
rect 112352 6205 112361 6239
rect 112361 6205 112395 6239
rect 112395 6205 112404 6239
rect 112352 6196 112404 6205
rect 126888 6264 126940 6316
rect 127532 6239 127584 6248
rect 127532 6205 127541 6239
rect 127541 6205 127575 6239
rect 127575 6205 127584 6239
rect 127532 6196 127584 6205
rect 127624 6196 127676 6248
rect 20628 6128 20680 6180
rect 32496 6128 32548 6180
rect 35532 6128 35584 6180
rect 126888 6128 126940 6180
rect 126980 6128 127032 6180
rect 171048 6128 171100 6180
rect 200580 6196 200632 6248
rect 217508 6332 217560 6384
rect 260748 6332 260800 6384
rect 213368 6264 213420 6316
rect 213644 6264 213696 6316
rect 202788 6239 202840 6248
rect 202788 6205 202797 6239
rect 202797 6205 202831 6239
rect 202831 6205 202840 6239
rect 202788 6196 202840 6205
rect 211528 6196 211580 6248
rect 212908 6239 212960 6248
rect 212908 6205 212917 6239
rect 212917 6205 212951 6239
rect 212951 6205 212960 6239
rect 212908 6196 212960 6205
rect 213276 6196 213328 6248
rect 214104 6239 214156 6248
rect 214104 6205 214113 6239
rect 214113 6205 214147 6239
rect 214147 6205 214156 6239
rect 214104 6196 214156 6205
rect 214932 6264 214984 6316
rect 215116 6196 215168 6248
rect 216496 6264 216548 6316
rect 220452 6264 220504 6316
rect 292580 6264 292632 6316
rect 292764 6307 292816 6316
rect 292764 6273 292773 6307
rect 292773 6273 292807 6307
rect 292807 6273 292816 6307
rect 292764 6264 292816 6273
rect 218428 6239 218480 6248
rect 218428 6205 218437 6239
rect 218437 6205 218471 6239
rect 218471 6205 218480 6239
rect 218428 6196 218480 6205
rect 261760 6239 261812 6248
rect 261760 6205 261769 6239
rect 261769 6205 261803 6239
rect 261803 6205 261812 6239
rect 261760 6196 261812 6205
rect 293316 6239 293368 6248
rect 293316 6205 293325 6239
rect 293325 6205 293359 6239
rect 293359 6205 293368 6239
rect 293316 6196 293368 6205
rect 310888 6307 310940 6316
rect 310888 6273 310897 6307
rect 310897 6273 310931 6307
rect 310931 6273 310940 6307
rect 310888 6264 310940 6273
rect 311900 6264 311952 6316
rect 313740 6264 313792 6316
rect 308680 6239 308732 6248
rect 308680 6205 308689 6239
rect 308689 6205 308723 6239
rect 308723 6205 308732 6239
rect 308680 6196 308732 6205
rect 23204 6060 23256 6112
rect 81532 6060 81584 6112
rect 119344 6103 119396 6112
rect 119344 6069 119353 6103
rect 119353 6069 119387 6103
rect 119387 6069 119396 6103
rect 119344 6060 119396 6069
rect 120448 6103 120500 6112
rect 120448 6069 120457 6103
rect 120457 6069 120491 6103
rect 120491 6069 120500 6103
rect 120448 6060 120500 6069
rect 121460 6103 121512 6112
rect 121460 6069 121469 6103
rect 121469 6069 121503 6103
rect 121503 6069 121512 6103
rect 121460 6060 121512 6069
rect 121828 6060 121880 6112
rect 203156 6128 203208 6180
rect 214932 6060 214984 6112
rect 216496 6103 216548 6112
rect 216496 6069 216505 6103
rect 216505 6069 216539 6103
rect 216539 6069 216548 6103
rect 216496 6060 216548 6069
rect 292672 6128 292724 6180
rect 339408 6239 339460 6248
rect 339408 6205 339417 6239
rect 339417 6205 339451 6239
rect 339451 6205 339460 6239
rect 339408 6196 339460 6205
rect 354588 6239 354640 6248
rect 354588 6205 354597 6239
rect 354597 6205 354631 6239
rect 354631 6205 354640 6239
rect 354588 6196 354640 6205
rect 292764 6060 292816 6112
rect 313740 6103 313792 6112
rect 313740 6069 313749 6103
rect 313749 6069 313783 6103
rect 313783 6069 313792 6103
rect 313740 6060 313792 6069
rect 338212 6103 338264 6112
rect 338212 6069 338221 6103
rect 338221 6069 338255 6103
rect 338255 6069 338264 6103
rect 338212 6060 338264 6069
rect 81921 5958 81973 6010
rect 81985 5958 82037 6010
rect 82049 5958 82101 6010
rect 82113 5958 82165 6010
rect 82177 5958 82229 6010
rect 243864 5958 243916 6010
rect 243928 5958 243980 6010
rect 243992 5958 244044 6010
rect 244056 5958 244108 6010
rect 244120 5958 244172 6010
rect 405807 5958 405859 6010
rect 405871 5958 405923 6010
rect 405935 5958 405987 6010
rect 405999 5958 406051 6010
rect 406063 5958 406115 6010
rect 567750 5958 567802 6010
rect 567814 5958 567866 6010
rect 567878 5958 567930 6010
rect 567942 5958 567994 6010
rect 568006 5958 568058 6010
rect 24308 5856 24360 5908
rect 116124 5856 116176 5908
rect 120448 5856 120500 5908
rect 212908 5856 212960 5908
rect 245476 5856 245528 5908
rect 338212 5856 338264 5908
rect 121460 5788 121512 5840
rect 214104 5788 214156 5840
rect 217876 5788 217928 5840
rect 80612 5720 80664 5772
rect 65064 5652 65116 5704
rect 23388 5584 23440 5636
rect 115664 5695 115716 5704
rect 115664 5661 115673 5695
rect 115673 5661 115707 5695
rect 115707 5661 115716 5695
rect 115664 5652 115716 5661
rect 199108 5720 199160 5772
rect 203156 5720 203208 5772
rect 201316 5652 201368 5704
rect 211528 5695 211580 5704
rect 211528 5661 211537 5695
rect 211537 5661 211571 5695
rect 211571 5661 211580 5695
rect 211528 5652 211580 5661
rect 119344 5584 119396 5636
rect 127624 5584 127676 5636
rect 157892 5627 157944 5636
rect 157892 5593 157901 5627
rect 157901 5593 157935 5627
rect 157935 5593 157944 5627
rect 157892 5584 157944 5593
rect 167000 5584 167052 5636
rect 173164 5584 173216 5636
rect 173256 5627 173308 5636
rect 173256 5593 173265 5627
rect 173265 5593 173299 5627
rect 173299 5593 173308 5627
rect 173256 5584 173308 5593
rect 247592 5695 247644 5704
rect 247592 5661 247601 5695
rect 247601 5661 247635 5695
rect 247635 5661 247644 5695
rect 247592 5652 247644 5661
rect 262956 5695 263008 5704
rect 262956 5661 262965 5695
rect 262965 5661 262999 5695
rect 262999 5661 263008 5695
rect 262956 5652 263008 5661
rect 311072 5652 311124 5704
rect 248972 5627 249024 5636
rect 248972 5593 248981 5627
rect 248981 5593 249015 5627
rect 249015 5593 249024 5627
rect 248972 5584 249024 5593
rect 264336 5627 264388 5636
rect 264336 5593 264345 5627
rect 264345 5593 264379 5627
rect 264379 5593 264388 5627
rect 264336 5584 264388 5593
rect 295064 5627 295116 5636
rect 295064 5593 295073 5627
rect 295073 5593 295107 5627
rect 295107 5593 295116 5627
rect 295064 5584 295116 5593
rect 28908 5516 28960 5568
rect 122564 5516 122616 5568
rect 212724 5559 212776 5568
rect 212724 5525 212733 5559
rect 212733 5525 212767 5559
rect 212767 5525 212776 5559
rect 212724 5516 212776 5525
rect 213736 5559 213788 5568
rect 213736 5525 213745 5559
rect 213745 5525 213779 5559
rect 213779 5525 213788 5559
rect 213736 5516 213788 5525
rect 215300 5559 215352 5568
rect 215300 5525 215309 5559
rect 215309 5525 215343 5559
rect 215343 5525 215352 5559
rect 215300 5516 215352 5525
rect 311900 5559 311952 5568
rect 311900 5525 311909 5559
rect 311909 5525 311943 5559
rect 311943 5525 311952 5559
rect 311900 5516 311952 5525
rect 82581 5414 82633 5466
rect 82645 5414 82697 5466
rect 82709 5414 82761 5466
rect 82773 5414 82825 5466
rect 82837 5414 82889 5466
rect 244524 5414 244576 5466
rect 244588 5414 244640 5466
rect 244652 5414 244704 5466
rect 244716 5414 244768 5466
rect 244780 5414 244832 5466
rect 406467 5414 406519 5466
rect 406531 5414 406583 5466
rect 406595 5414 406647 5466
rect 406659 5414 406711 5466
rect 406723 5414 406775 5466
rect 568410 5414 568462 5466
rect 568474 5414 568526 5466
rect 568538 5414 568590 5466
rect 568602 5414 568654 5466
rect 568666 5414 568718 5466
rect 308680 5312 308732 5364
rect 216496 5244 216548 5296
rect 111340 5040 111392 5092
rect 203892 5151 203944 5160
rect 203892 5117 203901 5151
rect 203901 5117 203935 5151
rect 203935 5117 203944 5151
rect 203892 5108 203944 5117
rect 126520 4972 126572 5024
rect 219164 5151 219216 5160
rect 219164 5117 219173 5151
rect 219173 5117 219207 5151
rect 219207 5117 219216 5151
rect 219164 5108 219216 5117
rect 262588 5244 262640 5296
rect 339868 5219 339920 5228
rect 339868 5185 339877 5219
rect 339877 5185 339911 5219
rect 339911 5185 339920 5219
rect 339868 5176 339920 5185
rect 309968 5151 310020 5160
rect 309968 5117 309977 5151
rect 309977 5117 310011 5151
rect 310011 5117 310020 5151
rect 309968 5108 310020 5117
rect 311072 5151 311124 5160
rect 311072 5117 311081 5151
rect 311081 5117 311115 5151
rect 311115 5117 311124 5151
rect 311072 5108 311124 5117
rect 293316 5040 293368 5092
rect 340696 5151 340748 5160
rect 340696 5117 340705 5151
rect 340705 5117 340739 5151
rect 340739 5117 340748 5151
rect 340696 5108 340748 5117
rect 355968 5151 356020 5160
rect 355968 5117 355977 5151
rect 355977 5117 356011 5151
rect 356011 5117 356020 5151
rect 355968 5108 356020 5117
rect 387064 5151 387116 5160
rect 387064 5117 387073 5151
rect 387073 5117 387107 5151
rect 387107 5117 387116 5151
rect 387064 5108 387116 5117
rect 402520 5151 402572 5160
rect 402520 5117 402529 5151
rect 402529 5117 402563 5151
rect 402563 5117 402572 5151
rect 402520 5108 402572 5117
rect 404544 5108 404596 5160
rect 432144 5219 432196 5228
rect 432144 5185 432153 5219
rect 432153 5185 432187 5219
rect 432187 5185 432196 5219
rect 432144 5176 432196 5185
rect 433248 5151 433300 5160
rect 433248 5117 433257 5151
rect 433257 5117 433291 5151
rect 433291 5117 433300 5151
rect 433248 5108 433300 5117
rect 448796 5151 448848 5160
rect 448796 5117 448805 5151
rect 448805 5117 448839 5151
rect 448839 5117 448848 5151
rect 448796 5108 448848 5117
rect 247316 4972 247368 5024
rect 339868 4972 339920 5024
rect 407304 5015 407356 5024
rect 407304 4981 407313 5015
rect 407313 4981 407347 5015
rect 407347 4981 407356 5015
rect 407304 4972 407356 4981
rect 447416 5015 447468 5024
rect 447416 4981 447425 5015
rect 447425 4981 447459 5015
rect 447459 4981 447468 5015
rect 447416 4972 447468 4981
rect 81921 4870 81973 4922
rect 81985 4870 82037 4922
rect 82049 4870 82101 4922
rect 82113 4870 82165 4922
rect 82177 4870 82229 4922
rect 243864 4870 243916 4922
rect 243928 4870 243980 4922
rect 243992 4870 244044 4922
rect 244056 4870 244108 4922
rect 244120 4870 244172 4922
rect 405807 4870 405859 4922
rect 405871 4870 405923 4922
rect 405935 4870 405987 4922
rect 405999 4870 406051 4922
rect 406063 4870 406115 4922
rect 567750 4870 567802 4922
rect 567814 4870 567866 4922
rect 567878 4870 567930 4922
rect 567942 4870 567994 4922
rect 568006 4870 568058 4922
rect 233884 4768 233936 4820
rect 249340 4768 249392 4820
rect 172244 4700 172296 4752
rect 239312 4700 239364 4752
rect 239496 4700 239548 4752
rect 264704 4768 264756 4820
rect 156972 4632 157024 4684
rect 233884 4632 233936 4684
rect 114468 4564 114520 4616
rect 211344 4564 211396 4616
rect 216588 4564 216640 4616
rect 23296 4496 23348 4548
rect 117964 4496 118016 4548
rect 202788 4428 202840 4480
rect 211344 4471 211396 4480
rect 211344 4437 211353 4471
rect 211353 4437 211387 4471
rect 211387 4437 211396 4471
rect 211344 4428 211396 4437
rect 215300 4496 215352 4548
rect 239404 4496 239456 4548
rect 239588 4428 239640 4480
rect 248788 4428 248840 4480
rect 249340 4607 249392 4616
rect 249340 4573 249349 4607
rect 249349 4573 249383 4607
rect 249383 4573 249392 4607
rect 249340 4564 249392 4573
rect 249708 4539 249760 4548
rect 249708 4505 249717 4539
rect 249717 4505 249751 4539
rect 249751 4505 249760 4539
rect 249708 4496 249760 4505
rect 249800 4496 249852 4548
rect 264704 4607 264756 4616
rect 264704 4573 264713 4607
rect 264713 4573 264747 4607
rect 264747 4573 264756 4607
rect 264704 4564 264756 4573
rect 265256 4539 265308 4548
rect 265256 4505 265265 4539
rect 265265 4505 265299 4539
rect 265299 4505 265308 4539
rect 265256 4496 265308 4505
rect 407304 4768 407356 4820
rect 499948 4768 500000 4820
rect 339408 4700 339460 4752
rect 432144 4700 432196 4752
rect 309324 4632 309376 4684
rect 295984 4539 296036 4548
rect 295984 4505 295993 4539
rect 295993 4505 296027 4539
rect 296027 4505 296036 4539
rect 295984 4496 296036 4505
rect 308864 4564 308916 4616
rect 354588 4632 354640 4684
rect 447416 4632 447468 4684
rect 310796 4564 310848 4616
rect 310336 4539 310388 4548
rect 310336 4505 310345 4539
rect 310345 4505 310379 4539
rect 310379 4505 310388 4539
rect 310336 4496 310388 4505
rect 311624 4539 311676 4548
rect 311624 4505 311633 4539
rect 311633 4505 311667 4539
rect 311667 4505 311676 4539
rect 311624 4496 311676 4505
rect 311900 4496 311952 4548
rect 313740 4428 313792 4480
rect 404544 4428 404596 4480
rect 406200 4428 406252 4480
rect 82581 4326 82633 4378
rect 82645 4326 82697 4378
rect 82709 4326 82761 4378
rect 82773 4326 82825 4378
rect 82837 4326 82889 4378
rect 244524 4326 244576 4378
rect 244588 4326 244640 4378
rect 244652 4326 244704 4378
rect 244716 4326 244768 4378
rect 244780 4326 244832 4378
rect 406467 4326 406519 4378
rect 406531 4326 406583 4378
rect 406595 4326 406647 4378
rect 406659 4326 406711 4378
rect 406723 4326 406775 4378
rect 568410 4326 568462 4378
rect 568474 4326 568526 4378
rect 568538 4326 568590 4378
rect 568602 4326 568654 4378
rect 568666 4326 568718 4378
rect 248788 4224 248840 4276
rect 249800 4224 249852 4276
rect 309324 4267 309376 4276
rect 309324 4233 309333 4267
rect 309333 4233 309367 4267
rect 309367 4233 309376 4267
rect 309324 4224 309376 4233
rect 218428 4156 218480 4208
rect 310796 4199 310848 4208
rect 310796 4165 310805 4199
rect 310805 4165 310839 4199
rect 310839 4165 310848 4199
rect 310796 4156 310848 4165
rect 248972 4088 249024 4140
rect 264336 4020 264388 4072
rect 213736 3952 213788 4004
rect 296720 4020 296772 4072
rect 306472 4131 306524 4140
rect 306472 4097 306481 4131
rect 306481 4097 306515 4131
rect 306515 4097 306524 4131
rect 306472 4088 306524 4097
rect 341340 4088 341392 4140
rect 307024 3952 307076 4004
rect 340696 4020 340748 4072
rect 342076 4020 342128 4072
rect 342720 4063 342772 4072
rect 342720 4029 342729 4063
rect 342729 4029 342763 4063
rect 342763 4029 342772 4063
rect 342720 4020 342772 4029
rect 355968 4088 356020 4140
rect 358084 4063 358136 4072
rect 358084 4029 358093 4063
rect 358093 4029 358127 4063
rect 358127 4029 358136 4063
rect 358084 4020 358136 4029
rect 387800 4131 387852 4140
rect 387800 4097 387809 4131
rect 387809 4097 387843 4131
rect 387843 4097 387852 4131
rect 387800 4088 387852 4097
rect 388996 4063 389048 4072
rect 388996 4029 389005 4063
rect 389005 4029 389039 4063
rect 389039 4029 389048 4063
rect 388996 4020 389048 4029
rect 402612 4088 402664 4140
rect 499948 4199 500000 4208
rect 499948 4165 499957 4199
rect 499957 4165 499991 4199
rect 499991 4165 500000 4199
rect 499948 4156 500000 4165
rect 404452 4063 404504 4072
rect 404452 4029 404461 4063
rect 404461 4029 404495 4063
rect 404495 4029 404504 4063
rect 404452 4020 404504 4029
rect 296720 3884 296772 3936
rect 306472 3884 306524 3936
rect 307116 3927 307168 3936
rect 307116 3893 307125 3927
rect 307125 3893 307159 3927
rect 307159 3893 307168 3927
rect 307116 3884 307168 3893
rect 308864 3927 308916 3936
rect 308864 3893 308873 3927
rect 308873 3893 308907 3927
rect 308907 3893 308916 3927
rect 308864 3884 308916 3893
rect 342260 3952 342312 4004
rect 479892 4088 479944 4140
rect 435364 4063 435416 4072
rect 435364 4029 435373 4063
rect 435373 4029 435407 4063
rect 435407 4029 435416 4063
rect 435364 4020 435416 4029
rect 450820 4063 450872 4072
rect 450820 4029 450829 4063
rect 450829 4029 450863 4063
rect 450863 4029 450872 4063
rect 450820 4020 450872 4029
rect 495440 4088 495492 4140
rect 497188 4063 497240 4072
rect 497188 4029 497197 4063
rect 497197 4029 497231 4063
rect 497231 4029 497240 4063
rect 497188 4020 497240 4029
rect 500500 4131 500552 4140
rect 500500 4097 500509 4131
rect 500509 4097 500543 4131
rect 500543 4097 500552 4131
rect 500500 4088 500552 4097
rect 619824 4020 619876 4072
rect 387800 3884 387852 3936
rect 402612 3927 402664 3936
rect 402612 3893 402621 3927
rect 402621 3893 402655 3927
rect 402655 3893 402664 3927
rect 402612 3884 402664 3893
rect 433248 3884 433300 3936
rect 573456 3952 573508 4004
rect 479892 3927 479944 3936
rect 479892 3893 479901 3927
rect 479901 3893 479935 3927
rect 479935 3893 479944 3927
rect 479892 3884 479944 3893
rect 495440 3927 495492 3936
rect 495440 3893 495449 3927
rect 495449 3893 495483 3927
rect 495483 3893 495492 3927
rect 495440 3884 495492 3893
rect 500500 3884 500552 3936
rect 594064 3884 594116 3936
rect 81921 3782 81973 3834
rect 81985 3782 82037 3834
rect 82049 3782 82101 3834
rect 82113 3782 82165 3834
rect 82177 3782 82229 3834
rect 243864 3782 243916 3834
rect 243928 3782 243980 3834
rect 243992 3782 244044 3834
rect 244056 3782 244108 3834
rect 244120 3782 244172 3834
rect 405807 3782 405859 3834
rect 405871 3782 405923 3834
rect 405935 3782 405987 3834
rect 405999 3782 406051 3834
rect 406063 3782 406115 3834
rect 567750 3782 567802 3834
rect 567814 3782 567866 3834
rect 567878 3782 567930 3834
rect 567942 3782 567994 3834
rect 568006 3782 568058 3834
rect 295064 3680 295116 3732
rect 307024 3680 307076 3732
rect 310336 3680 310388 3732
rect 402612 3680 402664 3732
rect 404452 3680 404504 3732
rect 496176 3680 496228 3732
rect 497188 3680 497240 3732
rect 588912 3680 588964 3732
rect 295984 3612 296036 3664
rect 387984 3612 388036 3664
rect 341340 3587 341392 3596
rect 341340 3553 341349 3587
rect 341349 3553 341383 3587
rect 341383 3553 341392 3587
rect 341340 3544 341392 3553
rect 387064 3544 387116 3596
rect 479892 3544 479944 3596
rect 233608 3476 233660 3528
rect 311072 3476 311124 3528
rect 117412 3408 117464 3460
rect 309968 3408 310020 3460
rect 403348 3476 403400 3528
rect 497280 3476 497332 3528
rect 499856 3476 499908 3528
rect 342720 3340 342772 3392
rect 406200 3408 406252 3460
rect 434352 3340 434404 3392
rect 448796 3340 448848 3392
rect 499856 3383 499908 3392
rect 499856 3349 499865 3383
rect 499865 3349 499899 3383
rect 499899 3349 499908 3383
rect 499856 3340 499908 3349
rect 635280 3408 635332 3460
rect 82581 3238 82633 3290
rect 82645 3238 82697 3290
rect 82709 3238 82761 3290
rect 82773 3238 82825 3290
rect 82837 3238 82889 3290
rect 244524 3238 244576 3290
rect 244588 3238 244640 3290
rect 244652 3238 244704 3290
rect 244716 3238 244768 3290
rect 244780 3238 244832 3290
rect 406467 3238 406519 3290
rect 406531 3238 406583 3290
rect 406595 3238 406647 3290
rect 406659 3238 406711 3290
rect 406723 3238 406775 3290
rect 568410 3238 568462 3290
rect 568474 3238 568526 3290
rect 568538 3238 568590 3290
rect 568602 3238 568654 3290
rect 568666 3238 568718 3290
rect 32496 3179 32548 3188
rect 32496 3145 32505 3179
rect 32505 3145 32539 3179
rect 32539 3145 32548 3179
rect 32496 3136 32548 3145
rect 112352 3136 112404 3188
rect 202512 3179 202564 3188
rect 202512 3145 202521 3179
rect 202521 3145 202555 3179
rect 202555 3145 202564 3179
rect 202512 3136 202564 3145
rect 203892 3136 203944 3188
rect 295708 3136 295760 3188
rect 22008 3068 22060 3120
rect 110236 3068 110288 3120
rect 173256 3068 173308 3120
rect 264796 3068 264848 3120
rect 265256 3068 265308 3120
rect 304816 3136 304868 3188
rect 326344 3136 326396 3188
rect 358084 3136 358136 3188
rect 450268 3136 450320 3188
rect 450820 3136 450872 3188
rect 543004 3136 543056 3188
rect 573456 3179 573508 3188
rect 573456 3145 573465 3179
rect 573465 3145 573499 3179
rect 573499 3145 573508 3179
rect 573456 3136 573508 3145
rect 588912 3179 588964 3188
rect 588912 3145 588921 3179
rect 588921 3145 588955 3179
rect 588955 3145 588964 3179
rect 588912 3136 588964 3145
rect 619824 3179 619876 3188
rect 619824 3145 619833 3179
rect 619833 3145 619867 3179
rect 619867 3145 619876 3179
rect 619824 3136 619876 3145
rect 635280 3179 635332 3188
rect 635280 3145 635289 3179
rect 635289 3145 635323 3179
rect 635323 3145 635332 3179
rect 635280 3136 635332 3145
rect 357072 3111 357124 3120
rect 37740 3000 37792 3052
rect 125232 3043 125284 3052
rect 125232 3009 125241 3043
rect 125241 3009 125275 3043
rect 125275 3009 125284 3043
rect 125232 3000 125284 3009
rect 127532 3000 127584 3052
rect 218428 3000 218480 3052
rect 219164 3000 219216 3052
rect 21916 2932 21968 2984
rect 79324 2932 79376 2984
rect 82452 2932 82504 2984
rect 172060 2932 172112 2984
rect 212724 2932 212776 2984
rect 304816 3000 304868 3052
rect 357072 3077 357081 3111
rect 357081 3077 357115 3111
rect 357115 3077 357124 3111
rect 357072 3068 357124 3077
rect 387984 3111 388036 3120
rect 387984 3077 387993 3111
rect 387993 3077 388027 3111
rect 388027 3077 388036 3111
rect 387984 3068 388036 3077
rect 308864 3000 308916 3052
rect 311164 2932 311216 2984
rect 21272 2864 21324 2916
rect 63868 2864 63920 2916
rect 66720 2864 66772 2916
rect 156604 2864 156656 2916
rect 157892 2864 157944 2916
rect 1584 2839 1636 2848
rect 1584 2805 1593 2839
rect 1593 2805 1627 2839
rect 1627 2805 1636 2839
rect 1584 2796 1636 2805
rect 47952 2839 48004 2848
rect 47952 2805 47961 2839
rect 47961 2805 47995 2839
rect 47995 2805 48004 2839
rect 47952 2796 48004 2805
rect 94320 2839 94372 2848
rect 94320 2805 94329 2839
rect 94329 2805 94363 2839
rect 94363 2805 94372 2839
rect 94320 2796 94372 2805
rect 141056 2796 141108 2848
rect 186872 2839 186924 2848
rect 186872 2805 186881 2839
rect 186881 2805 186915 2839
rect 186915 2805 186924 2839
rect 186872 2796 186924 2805
rect 233792 2796 233844 2848
rect 249708 2864 249760 2916
rect 248972 2796 249024 2848
rect 279608 2839 279660 2848
rect 279608 2805 279617 2839
rect 279617 2805 279651 2839
rect 279651 2805 279660 2839
rect 279608 2796 279660 2805
rect 326528 2796 326580 2848
rect 388996 2864 389048 2916
rect 342076 2796 342128 2848
rect 372620 2839 372672 2848
rect 372620 2805 372629 2839
rect 372629 2805 372663 2839
rect 372663 2805 372672 2839
rect 372620 2796 372672 2805
rect 434352 3111 434404 3120
rect 434352 3077 434361 3111
rect 434361 3077 434395 3111
rect 434395 3077 434404 3111
rect 434352 3068 434404 3077
rect 435364 3068 435416 3120
rect 527548 3068 527600 3120
rect 594064 3111 594116 3120
rect 594064 3077 594073 3111
rect 594073 3077 594107 3111
rect 594107 3077 594116 3111
rect 594064 3068 594116 3077
rect 402520 3000 402572 3052
rect 495440 3000 495492 3052
rect 496176 3043 496228 3052
rect 496176 3009 496185 3043
rect 496185 3009 496219 3043
rect 496219 3009 496228 3043
rect 496176 3000 496228 3009
rect 497280 3043 497332 3052
rect 497280 3009 497289 3043
rect 497289 3009 497323 3043
rect 497323 3009 497332 3043
rect 497280 3000 497332 3009
rect 510528 3000 510580 3052
rect 602896 3000 602948 3052
rect 403348 2975 403400 2984
rect 403348 2941 403357 2975
rect 403357 2941 403391 2975
rect 403391 2941 403400 2975
rect 403348 2932 403400 2941
rect 415308 2796 415360 2848
rect 465264 2839 465316 2848
rect 465264 2805 465273 2839
rect 465273 2805 465307 2839
rect 465307 2805 465316 2839
rect 465264 2796 465316 2805
rect 480812 2796 480864 2848
rect 558000 2839 558052 2848
rect 558000 2805 558009 2839
rect 558009 2805 558043 2839
rect 558043 2805 558052 2839
rect 558000 2796 558052 2805
rect 81921 2694 81973 2746
rect 81985 2694 82037 2746
rect 82049 2694 82101 2746
rect 82113 2694 82165 2746
rect 82177 2694 82229 2746
rect 243864 2694 243916 2746
rect 243928 2694 243980 2746
rect 243992 2694 244044 2746
rect 244056 2694 244108 2746
rect 244120 2694 244172 2746
rect 405807 2694 405859 2746
rect 405871 2694 405923 2746
rect 405935 2694 405987 2746
rect 405999 2694 406051 2746
rect 406063 2694 406115 2746
rect 567750 2694 567802 2746
rect 567814 2694 567866 2746
rect 567878 2694 567930 2746
rect 567942 2694 567994 2746
rect 568006 2694 568058 2746
rect 18052 2635 18104 2644
rect 18052 2601 18061 2635
rect 18061 2601 18095 2635
rect 18095 2601 18104 2635
rect 18052 2592 18104 2601
rect 415308 2592 415360 2644
rect 510528 2592 510580 2644
rect 602896 2592 602948 2644
rect 21824 2456 21876 2508
rect 233608 2567 233660 2576
rect 233608 2533 233617 2567
rect 233617 2533 233651 2567
rect 233651 2533 233660 2567
rect 233608 2524 233660 2533
rect 326344 2567 326396 2576
rect 326344 2533 326353 2567
rect 326353 2533 326387 2567
rect 326387 2533 326396 2567
rect 326344 2524 326396 2533
rect 115664 2456 115716 2508
rect 211344 2456 211396 2508
rect 311624 2456 311676 2508
rect 1584 2388 1636 2440
rect 18052 2388 18104 2440
rect 32496 2388 32548 2440
rect 47952 2388 48004 2440
rect 63868 2431 63920 2440
rect 63868 2397 63877 2431
rect 63877 2397 63911 2431
rect 63911 2397 63920 2431
rect 63868 2388 63920 2397
rect 79324 2431 79376 2440
rect 79324 2397 79333 2431
rect 79333 2397 79367 2431
rect 79367 2397 79376 2431
rect 79324 2388 79376 2397
rect 94320 2388 94372 2440
rect 110236 2431 110288 2440
rect 110236 2397 110245 2431
rect 110245 2397 110279 2431
rect 110279 2397 110288 2431
rect 110236 2388 110288 2397
rect 125232 2388 125284 2440
rect 156604 2431 156656 2440
rect 156604 2397 156613 2431
rect 156613 2397 156647 2431
rect 156647 2397 156656 2431
rect 156604 2388 156656 2397
rect 172060 2431 172112 2440
rect 172060 2397 172069 2431
rect 172069 2397 172103 2431
rect 172103 2397 172112 2431
rect 172060 2388 172112 2397
rect 202512 2388 202564 2440
rect 218428 2431 218480 2440
rect 218428 2397 218437 2431
rect 218437 2397 218471 2431
rect 218471 2397 218480 2431
rect 218428 2388 218480 2397
rect 248972 2388 249024 2440
rect 264796 2431 264848 2440
rect 264796 2397 264805 2431
rect 264805 2397 264839 2431
rect 264839 2397 264848 2431
rect 264796 2388 264848 2397
rect 295708 2431 295760 2440
rect 295708 2397 295717 2431
rect 295717 2397 295751 2431
rect 295751 2397 295760 2431
rect 295708 2388 295760 2397
rect 311164 2431 311216 2440
rect 311164 2397 311173 2431
rect 311173 2397 311207 2431
rect 311207 2397 311216 2431
rect 311164 2388 311216 2397
rect 17868 2320 17920 2372
rect 20996 2320 21048 2372
rect 15936 2252 15988 2304
rect 31668 2252 31720 2304
rect 114468 2320 114520 2372
rect 141056 2363 141108 2372
rect 141056 2329 141065 2363
rect 141065 2329 141099 2363
rect 141099 2329 141108 2363
rect 141056 2320 141108 2329
rect 186872 2320 186924 2372
rect 233792 2363 233844 2372
rect 233792 2329 233801 2363
rect 233801 2329 233835 2363
rect 233835 2329 233844 2363
rect 233792 2320 233844 2329
rect 279608 2320 279660 2372
rect 307116 2320 307168 2372
rect 326528 2363 326580 2372
rect 326528 2329 326537 2363
rect 326537 2329 326571 2363
rect 326571 2329 326580 2363
rect 326528 2320 326580 2329
rect 342076 2431 342128 2440
rect 342076 2397 342085 2431
rect 342085 2397 342119 2431
rect 342119 2397 342128 2431
rect 342076 2388 342128 2397
rect 357072 2388 357124 2440
rect 372620 2388 372672 2440
rect 387984 2388 388036 2440
rect 418068 2388 418120 2440
rect 434352 2388 434404 2440
rect 450268 2431 450320 2440
rect 450268 2397 450277 2431
rect 450277 2397 450311 2431
rect 450311 2397 450320 2431
rect 450268 2388 450320 2397
rect 465264 2388 465316 2440
rect 480812 2388 480864 2440
rect 496176 2388 496228 2440
rect 511908 2431 511960 2440
rect 511908 2397 511917 2431
rect 511917 2397 511951 2431
rect 511951 2397 511960 2431
rect 511908 2388 511960 2397
rect 527548 2431 527600 2440
rect 527548 2397 527557 2431
rect 527557 2397 527591 2431
rect 527591 2397 527600 2431
rect 527548 2388 527600 2397
rect 543004 2431 543056 2440
rect 543004 2397 543013 2431
rect 543013 2397 543047 2431
rect 543047 2397 543056 2431
rect 543004 2388 543056 2397
rect 558000 2388 558052 2440
rect 573456 2388 573508 2440
rect 588912 2388 588964 2440
rect 604368 2388 604420 2440
rect 619824 2388 619876 2440
rect 635280 2388 635332 2440
rect 62028 2252 62080 2304
rect 77208 2252 77260 2304
rect 107568 2252 107620 2304
rect 122656 2252 122708 2304
rect 156420 2295 156472 2304
rect 156420 2261 156429 2295
rect 156429 2261 156463 2295
rect 156463 2261 156472 2295
rect 156420 2252 156472 2261
rect 169668 2252 169720 2304
rect 199476 2252 199528 2304
rect 218244 2295 218296 2304
rect 218244 2261 218253 2295
rect 218253 2261 218287 2295
rect 218287 2261 218296 2295
rect 218244 2252 218296 2261
rect 249156 2295 249208 2304
rect 249156 2261 249165 2295
rect 249165 2261 249199 2295
rect 249199 2261 249208 2295
rect 249156 2252 249208 2261
rect 264612 2295 264664 2304
rect 264612 2261 264621 2295
rect 264621 2261 264655 2295
rect 264655 2261 264664 2295
rect 264612 2252 264664 2261
rect 293960 2252 294012 2304
rect 309140 2252 309192 2304
rect 339500 2252 339552 2304
rect 357348 2295 357400 2304
rect 357348 2261 357357 2295
rect 357357 2261 357391 2295
rect 357391 2261 357400 2295
rect 357348 2252 357400 2261
rect 403348 2320 403400 2372
rect 386420 2252 386472 2304
rect 402704 2252 402756 2304
rect 432788 2252 432840 2304
rect 450084 2295 450136 2304
rect 450084 2261 450093 2295
rect 450093 2261 450127 2295
rect 450127 2261 450136 2295
rect 450084 2252 450136 2261
rect 499856 2320 499908 2372
rect 480996 2295 481048 2304
rect 480996 2261 481005 2295
rect 481005 2261 481039 2295
rect 481039 2261 481048 2295
rect 480996 2252 481048 2261
rect 496452 2295 496504 2304
rect 496452 2261 496461 2295
rect 496461 2261 496495 2295
rect 496495 2261 496504 2295
rect 496452 2252 496504 2261
rect 527364 2295 527416 2304
rect 527364 2261 527373 2295
rect 527373 2261 527407 2295
rect 527407 2261 527416 2295
rect 527364 2252 527416 2261
rect 542820 2295 542872 2304
rect 542820 2261 542829 2295
rect 542829 2261 542863 2295
rect 542863 2261 542872 2295
rect 542820 2252 542872 2261
rect 573732 2295 573784 2304
rect 573732 2261 573741 2295
rect 573741 2261 573775 2295
rect 573775 2261 573784 2295
rect 573732 2252 573784 2261
rect 589188 2295 589240 2304
rect 589188 2261 589197 2295
rect 589197 2261 589231 2295
rect 589231 2261 589240 2295
rect 589188 2252 589240 2261
rect 618260 2252 618312 2304
rect 633440 2252 633492 2304
rect 82581 2150 82633 2202
rect 82645 2150 82697 2202
rect 82709 2150 82761 2202
rect 82773 2150 82825 2202
rect 82837 2150 82889 2202
rect 244524 2150 244576 2202
rect 244588 2150 244640 2202
rect 244652 2150 244704 2202
rect 244716 2150 244768 2202
rect 244780 2150 244832 2202
rect 406467 2150 406519 2202
rect 406531 2150 406583 2202
rect 406595 2150 406647 2202
rect 406659 2150 406711 2202
rect 406723 2150 406775 2202
rect 568410 2150 568462 2202
rect 568474 2150 568526 2202
rect 568538 2150 568590 2202
rect 568602 2150 568654 2202
rect 568666 2150 568718 2202
rect 1584 756 1636 808
rect 15936 756 15988 808
rect 31668 756 31720 808
rect 47952 756 48004 808
rect 62028 756 62080 808
rect 77208 756 77260 808
rect 94320 756 94372 808
rect 107568 756 107620 808
rect 122656 756 122708 808
rect 141056 756 141108 808
rect 156420 756 156472 808
rect 169668 756 169720 808
rect 186872 756 186924 808
rect 199476 756 199528 808
rect 218244 756 218296 808
rect 233792 756 233844 808
rect 249156 756 249208 808
rect 264612 756 264664 808
rect 279608 756 279660 808
rect 293960 756 294012 808
rect 309140 8 309192 60
rect 326528 756 326580 808
rect 339500 756 339552 808
rect 357348 756 357400 808
rect 372620 756 372672 808
rect 386420 8 386472 60
rect 402704 756 402756 808
rect 418068 756 418120 808
rect 432788 756 432840 808
rect 450084 756 450136 808
rect 465264 8 465316 60
rect 480996 756 481048 808
rect 496452 8 496504 60
rect 511908 756 511960 808
rect 527364 756 527416 808
rect 542820 8 542872 60
rect 558000 756 558052 808
rect 573732 8 573784 60
rect 589188 756 589240 808
rect 604368 756 604420 808
rect 618260 8 618312 60
rect 633440 756 633492 808
<< metal2 >>
rect -1076 9784 -756 9796
rect -1076 9728 -1064 9784
rect -1008 9728 -984 9784
rect -928 9728 -904 9784
rect -848 9728 -824 9784
rect -768 9728 -756 9784
rect -1076 9704 -756 9728
rect -1076 9648 -1064 9704
rect -1008 9648 -984 9704
rect -928 9648 -904 9704
rect -848 9648 -824 9704
rect -768 9648 -756 9704
rect -1076 9624 -756 9648
rect -1076 9568 -1064 9624
rect -1008 9568 -984 9624
rect -928 9568 -904 9624
rect -848 9568 -824 9624
rect -768 9568 -756 9624
rect -1076 9544 -756 9568
rect -1076 9488 -1064 9544
rect -1008 9488 -984 9544
rect -928 9488 -904 9544
rect -848 9488 -824 9544
rect -768 9488 -756 9544
rect -1076 7740 -756 9488
rect 30116 9302 30420 9330
rect 19708 9240 19760 9246
rect 19708 9182 19760 9188
rect 20168 9240 20220 9246
rect 20168 9182 20220 9188
rect 20996 9240 21048 9246
rect 20996 9182 21048 9188
rect 21272 9240 21324 9246
rect 21272 9182 21324 9188
rect 22928 9240 22980 9246
rect 22928 9182 22980 9188
rect 23204 9240 23256 9246
rect 23204 9182 23256 9188
rect 23756 9240 23808 9246
rect 23756 9182 23808 9188
rect 24308 9240 24360 9246
rect 24308 9182 24360 9188
rect 24584 9240 24636 9246
rect 24584 9182 24636 9188
rect 25136 9240 25188 9246
rect 25136 9182 25188 9188
rect 25688 9240 25740 9246
rect 25688 9182 25740 9188
rect 25964 9240 26016 9246
rect 25964 9182 26016 9188
rect 26148 9240 26200 9246
rect 26148 9182 26200 9188
rect 26700 9240 26752 9246
rect 26700 9182 26752 9188
rect 27252 9240 27304 9246
rect 27252 9182 27304 9188
rect 27528 9240 27580 9246
rect 27528 9182 27580 9188
rect 27804 9240 27856 9246
rect 27804 9182 27856 9188
rect 28080 9240 28132 9246
rect 28080 9182 28132 9188
rect 28356 9240 28408 9246
rect 28356 9182 28408 9188
rect 28908 9240 28960 9246
rect 28908 9182 28960 9188
rect 29184 9240 29236 9246
rect 29184 9182 29236 9188
rect 29460 9240 29512 9246
rect 29460 9182 29512 9188
rect 29736 9240 29788 9246
rect 29736 9182 29788 9188
rect 30012 9240 30064 9246
rect 30012 9182 30064 9188
rect -1076 7684 -1064 7740
rect -1008 7684 -984 7740
rect -928 7684 -904 7740
rect -848 7684 -824 7740
rect -768 7684 -756 7740
rect -1076 7660 -756 7684
rect -1076 7604 -1064 7660
rect -1008 7604 -984 7660
rect -928 7604 -904 7660
rect -848 7604 -824 7660
rect -768 7604 -756 7660
rect -1076 7580 -756 7604
rect -1076 7524 -1064 7580
rect -1008 7524 -984 7580
rect -928 7524 -904 7580
rect -848 7524 -824 7580
rect -768 7524 -756 7580
rect -1076 7500 -756 7524
rect -1076 7444 -1064 7500
rect -1008 7444 -984 7500
rect -928 7444 -904 7500
rect -848 7444 -824 7500
rect -768 7444 -756 7500
rect -1076 6381 -756 7444
rect -1076 6325 -1064 6381
rect -1008 6325 -984 6381
rect -928 6325 -904 6381
rect -848 6325 -824 6381
rect -768 6325 -756 6381
rect -1076 6301 -756 6325
rect -1076 6245 -1064 6301
rect -1008 6245 -984 6301
rect -928 6245 -904 6301
rect -848 6245 -824 6301
rect -768 6245 -756 6301
rect -1076 6221 -756 6245
rect -1076 6165 -1064 6221
rect -1008 6165 -984 6221
rect -928 6165 -904 6221
rect -848 6165 -824 6221
rect -768 6165 -756 6221
rect -1076 6141 -756 6165
rect -1076 6085 -1064 6141
rect -1008 6085 -984 6141
rect -928 6085 -904 6141
rect -848 6085 -824 6141
rect -768 6085 -756 6141
rect -1076 5022 -756 6085
rect -1076 4966 -1064 5022
rect -1008 4966 -984 5022
rect -928 4966 -904 5022
rect -848 4966 -824 5022
rect -768 4966 -756 5022
rect -1076 4942 -756 4966
rect -1076 4886 -1064 4942
rect -1008 4886 -984 4942
rect -928 4886 -904 4942
rect -848 4886 -824 4942
rect -768 4886 -756 4942
rect -1076 4862 -756 4886
rect -1076 4806 -1064 4862
rect -1008 4806 -984 4862
rect -928 4806 -904 4862
rect -848 4806 -824 4862
rect -768 4806 -756 4862
rect -1076 4782 -756 4806
rect -1076 4726 -1064 4782
rect -1008 4726 -984 4782
rect -928 4726 -904 4782
rect -848 4726 -824 4782
rect -768 4726 -756 4782
rect -1076 3663 -756 4726
rect -1076 3607 -1064 3663
rect -1008 3607 -984 3663
rect -928 3607 -904 3663
rect -848 3607 -824 3663
rect -768 3607 -756 3663
rect -1076 3583 -756 3607
rect -1076 3527 -1064 3583
rect -1008 3527 -984 3583
rect -928 3527 -904 3583
rect -848 3527 -824 3583
rect -768 3527 -756 3583
rect -1076 3503 -756 3527
rect -1076 3447 -1064 3503
rect -1008 3447 -984 3503
rect -928 3447 -904 3503
rect -848 3447 -824 3503
rect -768 3447 -756 3503
rect -1076 3423 -756 3447
rect -1076 3367 -1064 3423
rect -1008 3367 -984 3423
rect -928 3367 -904 3423
rect -848 3367 -824 3423
rect -768 3367 -756 3423
rect -1076 304 -756 3367
rect -416 9124 -96 9136
rect -416 9068 -404 9124
rect -348 9068 -324 9124
rect -268 9068 -244 9124
rect -188 9068 -164 9124
rect -108 9068 -96 9124
rect -416 9044 -96 9068
rect -416 8988 -404 9044
rect -348 8988 -324 9044
rect -268 8988 -244 9044
rect -188 8988 -164 9044
rect -108 8988 -96 9044
rect -416 8964 -96 8988
rect -416 8908 -404 8964
rect -348 8908 -324 8964
rect -268 8908 -244 8964
rect -188 8908 -164 8964
rect -108 8908 -96 8964
rect -416 8884 -96 8908
rect -416 8828 -404 8884
rect -348 8828 -324 8884
rect -268 8828 -244 8884
rect -188 8828 -164 8884
rect -108 8828 -96 8884
rect -416 7080 -96 8828
rect -416 7024 -404 7080
rect -348 7024 -324 7080
rect -268 7024 -244 7080
rect -188 7024 -164 7080
rect -108 7024 -96 7080
rect -416 7000 -96 7024
rect -416 6944 -404 7000
rect -348 6944 -324 7000
rect -268 6944 -244 7000
rect -188 6944 -164 7000
rect -108 6944 -96 7000
rect -416 6920 -96 6944
rect -416 6864 -404 6920
rect -348 6864 -324 6920
rect -268 6864 -244 6920
rect -188 6864 -164 6920
rect -108 6864 -96 6920
rect 19720 6866 19748 9182
rect -416 6840 -96 6864
rect -416 6784 -404 6840
rect -348 6784 -324 6840
rect -268 6784 -244 6840
rect -188 6784 -164 6840
rect -108 6784 -96 6840
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 19708 6860 19760 6866
rect 19708 6802 19760 6808
rect -416 5721 -96 6784
rect -416 5665 -404 5721
rect -348 5665 -324 5721
rect -268 5665 -244 5721
rect -188 5665 -164 5721
rect -108 5665 -96 5721
rect -416 5641 -96 5665
rect -416 5585 -404 5641
rect -348 5585 -324 5641
rect -268 5585 -244 5641
rect -188 5585 -164 5641
rect -108 5585 -96 5641
rect -416 5561 -96 5585
rect -416 5505 -404 5561
rect -348 5505 -324 5561
rect -268 5505 -244 5561
rect -188 5505 -164 5561
rect -108 5505 -96 5561
rect -416 5481 -96 5505
rect -416 5425 -404 5481
rect -348 5425 -324 5481
rect -268 5425 -244 5481
rect -188 5425 -164 5481
rect -108 5425 -96 5481
rect -416 4362 -96 5425
rect -416 4306 -404 4362
rect -348 4306 -324 4362
rect -268 4306 -244 4362
rect -188 4306 -164 4362
rect -108 4306 -96 4362
rect -416 4282 -96 4306
rect -416 4226 -404 4282
rect -348 4226 -324 4282
rect -268 4226 -244 4282
rect -188 4226 -164 4282
rect -108 4226 -96 4282
rect -416 4202 -96 4226
rect -416 4146 -404 4202
rect -348 4146 -324 4202
rect -268 4146 -244 4202
rect -188 4146 -164 4202
rect -108 4146 -96 4202
rect -416 4122 -96 4146
rect -416 4066 -404 4122
rect -348 4066 -324 4122
rect -268 4066 -244 4122
rect -188 4066 -164 4122
rect -108 4066 -96 4122
rect -416 3003 -96 4066
rect -416 2947 -404 3003
rect -348 2947 -324 3003
rect -268 2947 -244 3003
rect -188 2947 -164 3003
rect -108 2947 -96 3003
rect -416 2923 -96 2947
rect -416 2867 -404 2923
rect -348 2867 -324 2923
rect -268 2867 -244 2923
rect -188 2867 -164 2923
rect -108 2867 -96 2923
rect -416 2843 -96 2867
rect -416 2787 -404 2843
rect -348 2787 -324 2843
rect -268 2787 -244 2843
rect -188 2787 -164 2843
rect -108 2787 -96 2843
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect -416 2763 -96 2787
rect -416 2707 -404 2763
rect -348 2707 -324 2763
rect -268 2707 -244 2763
rect -188 2707 -164 2763
rect -108 2707 -96 2763
rect -416 964 -96 2707
rect 1596 2446 1624 2790
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect -416 908 -404 964
rect -348 908 -324 964
rect -268 908 -244 964
rect -188 908 -164 964
rect -108 908 -96 964
rect -416 884 -96 908
rect -416 828 -404 884
rect -348 828 -324 884
rect -268 828 -244 884
rect -188 828 -164 884
rect -108 828 -96 884
rect -416 804 -96 828
rect 1596 814 1624 2382
rect 17880 2378 17908 6802
rect 20180 6798 20208 9182
rect 20628 8900 20680 8906
rect 20628 8842 20680 8848
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 18064 2650 18092 6734
rect 20640 6186 20668 8842
rect 20628 6180 20680 6186
rect 20628 6122 20680 6128
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 18064 2446 18092 2586
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 21008 2378 21036 9182
rect 21284 2922 21312 9182
rect 21824 8968 21876 8974
rect 21824 8910 21876 8916
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 21272 2916 21324 2922
rect 21272 2858 21324 2864
rect 21836 2514 21864 8910
rect 21916 8900 21968 8906
rect 21916 8842 21968 8848
rect 21928 2990 21956 8842
rect 22020 3126 22048 8910
rect 22940 8158 22968 9182
rect 22928 8152 22980 8158
rect 22928 8094 22980 8100
rect 23216 6118 23244 9182
rect 23388 9172 23440 9178
rect 23388 9114 23440 9120
rect 23296 8968 23348 8974
rect 23296 8910 23348 8916
rect 23204 6112 23256 6118
rect 23204 6054 23256 6060
rect 23308 4554 23336 8910
rect 23400 5642 23428 9114
rect 23768 6390 23796 9182
rect 23756 6384 23808 6390
rect 23756 6326 23808 6332
rect 24320 5914 24348 9182
rect 24596 7002 24624 9182
rect 24768 9172 24820 9178
rect 24768 9114 24820 9120
rect 24780 8022 24808 9114
rect 24768 8016 24820 8022
rect 24768 7958 24820 7964
rect 25148 7546 25176 9182
rect 25700 8498 25728 9182
rect 25688 8492 25740 8498
rect 25688 8434 25740 8440
rect 25136 7540 25188 7546
rect 25136 7482 25188 7488
rect 25976 7478 26004 9182
rect 26160 8566 26188 9182
rect 26148 8560 26200 8566
rect 26148 8502 26200 8508
rect 25964 7472 26016 7478
rect 25964 7414 26016 7420
rect 24584 6996 24636 7002
rect 24584 6938 24636 6944
rect 26712 6866 26740 9182
rect 27264 8430 27292 9182
rect 27252 8424 27304 8430
rect 27252 8366 27304 8372
rect 26700 6860 26752 6866
rect 26700 6802 26752 6808
rect 27540 6322 27568 9182
rect 27816 7818 27844 9182
rect 28092 8090 28120 9182
rect 28368 8129 28396 9182
rect 28354 8120 28410 8129
rect 28080 8084 28132 8090
rect 28354 8055 28410 8064
rect 28080 8026 28132 8032
rect 27804 7812 27856 7818
rect 27804 7754 27856 7760
rect 27528 6316 27580 6322
rect 27528 6258 27580 6264
rect 24308 5908 24360 5914
rect 24308 5850 24360 5856
rect 23388 5636 23440 5642
rect 23388 5578 23440 5584
rect 28920 5574 28948 9182
rect 29196 7993 29224 9182
rect 29182 7984 29238 7993
rect 29182 7919 29238 7928
rect 29472 7274 29500 9182
rect 29748 8770 29776 9182
rect 29736 8764 29788 8770
rect 29736 8706 29788 8712
rect 29460 7268 29512 7274
rect 29460 7210 29512 7216
rect 30024 6730 30052 9182
rect 30116 9178 30144 9302
rect 30104 9172 30156 9178
rect 30104 9114 30156 9120
rect 30288 9104 30340 9110
rect 30288 9046 30340 9052
rect 30300 8702 30328 9046
rect 30392 8974 30420 9302
rect 30840 9240 30892 9246
rect 30840 9182 30892 9188
rect 31116 9240 31168 9246
rect 31116 9182 31168 9188
rect 31484 9240 31536 9246
rect 31484 9182 31536 9188
rect 30472 9172 30524 9178
rect 30472 9114 30524 9120
rect 30380 8968 30432 8974
rect 30380 8910 30432 8916
rect 30484 8906 30512 9114
rect 30472 8900 30524 8906
rect 30472 8842 30524 8848
rect 30288 8696 30340 8702
rect 30288 8638 30340 8644
rect 30380 8696 30432 8702
rect 30380 8638 30432 8644
rect 30196 8560 30248 8566
rect 30392 8514 30420 8638
rect 30248 8508 30420 8514
rect 30196 8502 30420 8508
rect 30656 8560 30708 8566
rect 30656 8502 30708 8508
rect 30208 8486 30420 8502
rect 30668 8294 30696 8502
rect 30656 8288 30708 8294
rect 30656 8230 30708 8236
rect 30012 6724 30064 6730
rect 30012 6666 30064 6672
rect 30852 6633 30880 9182
rect 31128 7954 31156 9182
rect 31116 7948 31168 7954
rect 31116 7890 31168 7896
rect 31496 7750 31524 9182
rect 81915 9124 82235 9796
rect 81915 9068 81927 9124
rect 81983 9068 82007 9124
rect 82063 9068 82087 9124
rect 82143 9068 82167 9124
rect 82223 9068 82235 9124
rect 81915 9044 82235 9068
rect 81915 8988 81927 9044
rect 81983 8988 82007 9044
rect 82063 8988 82087 9044
rect 82143 8988 82167 9044
rect 82223 8988 82235 9044
rect 81915 8964 82235 8988
rect 81915 8908 81927 8964
rect 81983 8908 82007 8964
rect 82063 8908 82087 8964
rect 82143 8908 82167 8964
rect 82223 8908 82235 8964
rect 81915 8884 82235 8908
rect 78036 8832 78088 8838
rect 78036 8774 78088 8780
rect 81915 8828 81927 8884
rect 81983 8828 82007 8884
rect 82063 8828 82087 8884
rect 82143 8828 82167 8884
rect 82223 8828 82235 8884
rect 74080 8764 74132 8770
rect 74080 8706 74132 8712
rect 62580 8696 62632 8702
rect 62580 8638 62632 8644
rect 35256 8628 35308 8634
rect 35256 8570 35308 8576
rect 36820 8628 36872 8634
rect 36820 8570 36872 8576
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 31484 7744 31536 7750
rect 31484 7686 31536 7692
rect 32692 7410 32720 8434
rect 33508 7880 33560 7886
rect 33508 7822 33560 7828
rect 33520 7410 33548 7822
rect 35268 7410 35296 8570
rect 36832 7410 36860 8570
rect 57336 8288 57388 8294
rect 57336 8230 57388 8236
rect 56600 7948 56652 7954
rect 56600 7890 56652 7896
rect 56612 7410 56640 7890
rect 57348 7410 57376 8230
rect 60924 7812 60976 7818
rect 60924 7754 60976 7760
rect 60936 7410 60964 7754
rect 62592 7410 62620 8638
rect 65892 8152 65944 8158
rect 65892 8094 65944 8100
rect 72792 8152 72844 8158
rect 72792 8094 72844 8100
rect 65904 7410 65932 8094
rect 71964 7744 72016 7750
rect 71964 7686 72016 7692
rect 71976 7410 72004 7686
rect 72804 7410 72832 8094
rect 74092 7410 74120 8706
rect 74908 8220 74960 8226
rect 74908 8162 74960 8168
rect 74920 7410 74948 8162
rect 76104 8084 76156 8090
rect 76104 8026 76156 8032
rect 76116 7410 76144 8026
rect 76932 7948 76984 7954
rect 76932 7890 76984 7896
rect 76944 7410 76972 7890
rect 78048 7410 78076 8774
rect 79968 8016 80020 8022
rect 79968 7958 80020 7964
rect 79980 7410 80008 7958
rect 32680 7404 32732 7410
rect 32680 7346 32732 7352
rect 33508 7404 33560 7410
rect 33508 7346 33560 7352
rect 35256 7404 35308 7410
rect 35256 7346 35308 7352
rect 36820 7404 36872 7410
rect 36820 7346 36872 7352
rect 56600 7404 56652 7410
rect 56600 7346 56652 7352
rect 57336 7404 57388 7410
rect 57336 7346 57388 7352
rect 60924 7404 60976 7410
rect 60924 7346 60976 7352
rect 62580 7404 62632 7410
rect 62580 7346 62632 7352
rect 63040 7404 63092 7410
rect 63040 7346 63092 7352
rect 64788 7404 64840 7410
rect 64788 7346 64840 7352
rect 65892 7404 65944 7410
rect 65892 7346 65944 7352
rect 71964 7404 72016 7410
rect 71964 7346 72016 7352
rect 72792 7404 72844 7410
rect 72792 7346 72844 7352
rect 74080 7404 74132 7410
rect 74080 7346 74132 7352
rect 74908 7404 74960 7410
rect 74908 7346 74960 7352
rect 76104 7404 76156 7410
rect 76104 7346 76156 7352
rect 76932 7404 76984 7410
rect 76932 7346 76984 7352
rect 78036 7404 78088 7410
rect 78036 7346 78088 7352
rect 79600 7404 79652 7410
rect 79600 7346 79652 7352
rect 79968 7404 80020 7410
rect 79968 7346 80020 7352
rect 35268 6934 35296 7346
rect 35532 7336 35584 7342
rect 35532 7278 35584 7284
rect 37740 7336 37792 7342
rect 37740 7278 37792 7284
rect 59636 7336 59688 7342
rect 59636 7278 59688 7284
rect 35256 6928 35308 6934
rect 35256 6870 35308 6876
rect 30838 6624 30894 6633
rect 30838 6559 30894 6568
rect 35544 6186 35572 7278
rect 32496 6180 32548 6186
rect 32496 6122 32548 6128
rect 35532 6180 35584 6186
rect 35532 6122 35584 6128
rect 28908 5568 28960 5574
rect 28908 5510 28960 5516
rect 23296 4548 23348 4554
rect 23296 4490 23348 4496
rect 32508 3194 32536 6122
rect 32496 3188 32548 3194
rect 32496 3130 32548 3136
rect 22008 3120 22060 3126
rect 22008 3062 22060 3068
rect 21916 2984 21968 2990
rect 21916 2926 21968 2932
rect 21824 2508 21876 2514
rect 21824 2450 21876 2456
rect 32508 2446 32536 3130
rect 37752 3058 37780 7278
rect 59648 7002 59676 7278
rect 59636 6996 59688 7002
rect 59636 6938 59688 6944
rect 63052 6798 63080 7346
rect 63776 7336 63828 7342
rect 63776 7278 63828 7284
rect 63040 6792 63092 6798
rect 63040 6734 63092 6740
rect 63788 6458 63816 7278
rect 64800 6934 64828 7346
rect 65064 7336 65116 7342
rect 65064 7278 65116 7284
rect 66720 7336 66772 7342
rect 66720 7278 66772 7284
rect 79324 7336 79376 7342
rect 79324 7278 79376 7284
rect 64788 6928 64840 6934
rect 64788 6870 64840 6876
rect 63776 6452 63828 6458
rect 63776 6394 63828 6400
rect 65076 5710 65104 7278
rect 65064 5704 65116 5710
rect 65064 5646 65116 5652
rect 37740 3052 37792 3058
rect 37740 2994 37792 3000
rect 66732 2922 66760 7278
rect 79336 5953 79364 7278
rect 79612 6798 79640 7346
rect 80612 7336 80664 7342
rect 80612 7278 80664 7284
rect 79600 6792 79652 6798
rect 79600 6734 79652 6740
rect 79322 5944 79378 5953
rect 79322 5879 79378 5888
rect 80624 5778 80652 7278
rect 81915 7098 82235 8828
rect 81915 7046 81921 7098
rect 81973 7080 81985 7098
rect 82037 7080 82049 7098
rect 82101 7080 82113 7098
rect 82165 7080 82177 7098
rect 81983 7046 81985 7080
rect 82165 7046 82167 7080
rect 82229 7046 82235 7098
rect 81915 7024 81927 7046
rect 81983 7024 82007 7046
rect 82063 7024 82087 7046
rect 82143 7024 82167 7046
rect 82223 7024 82235 7046
rect 81915 7000 82235 7024
rect 81915 6944 81927 7000
rect 81983 6944 82007 7000
rect 82063 6944 82087 7000
rect 82143 6944 82167 7000
rect 82223 6944 82235 7000
rect 81915 6920 82235 6944
rect 81915 6864 81927 6920
rect 81983 6864 82007 6920
rect 82063 6864 82087 6920
rect 82143 6864 82167 6920
rect 82223 6864 82235 6920
rect 81915 6840 82235 6864
rect 81532 6792 81584 6798
rect 81532 6734 81584 6740
rect 81915 6784 81927 6840
rect 81983 6784 82007 6840
rect 82063 6784 82087 6840
rect 82143 6784 82167 6840
rect 82223 6784 82235 6840
rect 81544 6118 81572 6734
rect 81532 6112 81584 6118
rect 81532 6054 81584 6060
rect 81915 6010 82235 6784
rect 82575 9784 82895 9796
rect 82575 9728 82587 9784
rect 82643 9728 82667 9784
rect 82723 9728 82747 9784
rect 82803 9728 82827 9784
rect 82883 9728 82895 9784
rect 82575 9704 82895 9728
rect 82575 9648 82587 9704
rect 82643 9648 82667 9704
rect 82723 9648 82747 9704
rect 82803 9648 82827 9704
rect 82883 9648 82895 9704
rect 82575 9624 82895 9648
rect 82575 9568 82587 9624
rect 82643 9568 82667 9624
rect 82723 9568 82747 9624
rect 82803 9568 82827 9624
rect 82883 9568 82895 9624
rect 82575 9544 82895 9568
rect 82575 9488 82587 9544
rect 82643 9488 82667 9544
rect 82723 9488 82747 9544
rect 82803 9488 82827 9544
rect 82883 9488 82895 9544
rect 82575 7740 82895 9488
rect 118976 9172 119028 9178
rect 118976 9114 119028 9120
rect 243858 9124 244178 9796
rect 110144 9104 110196 9110
rect 110144 9046 110196 9052
rect 108488 9036 108540 9042
rect 108488 8978 108540 8984
rect 107292 8968 107344 8974
rect 107292 8910 107344 8916
rect 104624 8900 104676 8906
rect 104624 8842 104676 8848
rect 82575 7684 82587 7740
rect 82643 7684 82667 7740
rect 82723 7684 82747 7740
rect 82803 7684 82827 7740
rect 82883 7684 82895 7740
rect 82575 7660 82895 7684
rect 82575 7642 82587 7660
rect 82643 7642 82667 7660
rect 82723 7642 82747 7660
rect 82803 7642 82827 7660
rect 82883 7642 82895 7660
rect 82575 7590 82581 7642
rect 82643 7604 82645 7642
rect 82825 7604 82827 7642
rect 82633 7590 82645 7604
rect 82697 7590 82709 7604
rect 82761 7590 82773 7604
rect 82825 7590 82837 7604
rect 82889 7590 82895 7642
rect 82575 7580 82895 7590
rect 82575 7524 82587 7580
rect 82643 7524 82667 7580
rect 82723 7524 82747 7580
rect 82803 7524 82827 7580
rect 82883 7524 82895 7580
rect 82575 7500 82895 7524
rect 82575 7444 82587 7500
rect 82643 7444 82667 7500
rect 82723 7444 82747 7500
rect 82803 7444 82827 7500
rect 82883 7444 82895 7500
rect 82452 6724 82504 6730
rect 82452 6666 82504 6672
rect 81915 5958 81921 6010
rect 81973 5958 81985 6010
rect 82037 5958 82049 6010
rect 82101 5958 82113 6010
rect 82165 5958 82177 6010
rect 82229 5958 82235 6010
rect 80612 5772 80664 5778
rect 80612 5714 80664 5720
rect 81915 5721 82235 5958
rect 81915 5665 81927 5721
rect 81983 5665 82007 5721
rect 82063 5665 82087 5721
rect 82143 5665 82167 5721
rect 82223 5665 82235 5721
rect 81915 5641 82235 5665
rect 81915 5585 81927 5641
rect 81983 5585 82007 5641
rect 82063 5585 82087 5641
rect 82143 5585 82167 5641
rect 82223 5585 82235 5641
rect 81915 5561 82235 5585
rect 81915 5505 81927 5561
rect 81983 5505 82007 5561
rect 82063 5505 82087 5561
rect 82143 5505 82167 5561
rect 82223 5505 82235 5561
rect 81915 5481 82235 5505
rect 81915 5425 81927 5481
rect 81983 5425 82007 5481
rect 82063 5425 82087 5481
rect 82143 5425 82167 5481
rect 82223 5425 82235 5481
rect 81915 4922 82235 5425
rect 81915 4870 81921 4922
rect 81973 4870 81985 4922
rect 82037 4870 82049 4922
rect 82101 4870 82113 4922
rect 82165 4870 82177 4922
rect 82229 4870 82235 4922
rect 81915 4362 82235 4870
rect 81915 4306 81927 4362
rect 81983 4306 82007 4362
rect 82063 4306 82087 4362
rect 82143 4306 82167 4362
rect 82223 4306 82235 4362
rect 81915 4282 82235 4306
rect 81915 4226 81927 4282
rect 81983 4226 82007 4282
rect 82063 4226 82087 4282
rect 82143 4226 82167 4282
rect 82223 4226 82235 4282
rect 81915 4202 82235 4226
rect 81915 4146 81927 4202
rect 81983 4146 82007 4202
rect 82063 4146 82087 4202
rect 82143 4146 82167 4202
rect 82223 4146 82235 4202
rect 81915 4122 82235 4146
rect 81915 4066 81927 4122
rect 81983 4066 82007 4122
rect 82063 4066 82087 4122
rect 82143 4066 82167 4122
rect 82223 4066 82235 4122
rect 81915 3834 82235 4066
rect 81915 3782 81921 3834
rect 81973 3782 81985 3834
rect 82037 3782 82049 3834
rect 82101 3782 82113 3834
rect 82165 3782 82177 3834
rect 82229 3782 82235 3834
rect 81915 3003 82235 3782
rect 79324 2984 79376 2990
rect 79324 2926 79376 2932
rect 81915 2947 81927 3003
rect 81983 2947 82007 3003
rect 82063 2947 82087 3003
rect 82143 2947 82167 3003
rect 82223 2947 82235 3003
rect 82464 2990 82492 6666
rect 82575 6554 82895 7444
rect 104636 7410 104664 8842
rect 105820 7744 105872 7750
rect 105820 7686 105872 7692
rect 105832 7410 105860 7686
rect 107304 7410 107332 8910
rect 107844 7812 107896 7818
rect 107844 7754 107896 7760
rect 107856 7478 107884 7754
rect 107844 7472 107896 7478
rect 107844 7414 107896 7420
rect 104624 7404 104676 7410
rect 104624 7346 104676 7352
rect 105820 7404 105872 7410
rect 105820 7346 105872 7352
rect 107292 7404 107344 7410
rect 107292 7346 107344 7352
rect 107304 6934 107332 7346
rect 107292 6928 107344 6934
rect 107292 6870 107344 6876
rect 108500 6798 108528 8978
rect 110156 7410 110184 9046
rect 110144 7404 110196 7410
rect 110144 7346 110196 7352
rect 117964 7404 118016 7410
rect 117964 7346 118016 7352
rect 111340 7336 111392 7342
rect 111340 7278 111392 7284
rect 108488 6792 108540 6798
rect 108488 6734 108540 6740
rect 82575 6502 82581 6554
rect 82633 6502 82645 6554
rect 82697 6502 82709 6554
rect 82761 6502 82773 6554
rect 82825 6502 82837 6554
rect 82889 6502 82895 6554
rect 82575 6381 82895 6502
rect 82575 6325 82587 6381
rect 82643 6325 82667 6381
rect 82723 6325 82747 6381
rect 82803 6325 82827 6381
rect 82883 6325 82895 6381
rect 82575 6301 82895 6325
rect 82575 6245 82587 6301
rect 82643 6245 82667 6301
rect 82723 6245 82747 6301
rect 82803 6245 82827 6301
rect 82883 6245 82895 6301
rect 82575 6221 82895 6245
rect 82575 6165 82587 6221
rect 82643 6165 82667 6221
rect 82723 6165 82747 6221
rect 82803 6165 82827 6221
rect 82883 6165 82895 6221
rect 82575 6141 82895 6165
rect 82575 6085 82587 6141
rect 82643 6085 82667 6141
rect 82723 6085 82747 6141
rect 82803 6085 82827 6141
rect 82883 6085 82895 6141
rect 82575 5466 82895 6085
rect 82575 5414 82581 5466
rect 82633 5414 82645 5466
rect 82697 5414 82709 5466
rect 82761 5414 82773 5466
rect 82825 5414 82837 5466
rect 82889 5414 82895 5466
rect 82575 5022 82895 5414
rect 111352 5098 111380 7278
rect 117044 6792 117096 6798
rect 117096 6740 117452 6746
rect 117044 6734 117452 6740
rect 116124 6724 116176 6730
rect 117056 6718 117452 6734
rect 116124 6666 116176 6672
rect 112352 6248 112404 6254
rect 112352 6190 112404 6196
rect 111340 5092 111392 5098
rect 111340 5034 111392 5040
rect 82575 4966 82587 5022
rect 82643 4966 82667 5022
rect 82723 4966 82747 5022
rect 82803 4966 82827 5022
rect 82883 4966 82895 5022
rect 82575 4942 82895 4966
rect 82575 4886 82587 4942
rect 82643 4886 82667 4942
rect 82723 4886 82747 4942
rect 82803 4886 82827 4942
rect 82883 4886 82895 4942
rect 82575 4862 82895 4886
rect 82575 4806 82587 4862
rect 82643 4806 82667 4862
rect 82723 4806 82747 4862
rect 82803 4806 82827 4862
rect 82883 4806 82895 4862
rect 82575 4782 82895 4806
rect 82575 4726 82587 4782
rect 82643 4726 82667 4782
rect 82723 4726 82747 4782
rect 82803 4726 82827 4782
rect 82883 4726 82895 4782
rect 82575 4378 82895 4726
rect 82575 4326 82581 4378
rect 82633 4326 82645 4378
rect 82697 4326 82709 4378
rect 82761 4326 82773 4378
rect 82825 4326 82837 4378
rect 82889 4326 82895 4378
rect 82575 3663 82895 4326
rect 82575 3607 82587 3663
rect 82643 3607 82667 3663
rect 82723 3607 82747 3663
rect 82803 3607 82827 3663
rect 82883 3607 82895 3663
rect 82575 3583 82895 3607
rect 82575 3527 82587 3583
rect 82643 3527 82667 3583
rect 82723 3527 82747 3583
rect 82803 3527 82827 3583
rect 82883 3527 82895 3583
rect 82575 3503 82895 3527
rect 82575 3447 82587 3503
rect 82643 3447 82667 3503
rect 82723 3447 82747 3503
rect 82803 3447 82827 3503
rect 82883 3447 82895 3503
rect 82575 3423 82895 3447
rect 82575 3367 82587 3423
rect 82643 3367 82667 3423
rect 82723 3367 82747 3423
rect 82803 3367 82827 3423
rect 82883 3367 82895 3423
rect 82575 3290 82895 3367
rect 82575 3238 82581 3290
rect 82633 3238 82645 3290
rect 82697 3238 82709 3290
rect 82761 3238 82773 3290
rect 82825 3238 82837 3290
rect 82889 3238 82895 3290
rect 63868 2916 63920 2922
rect 63868 2858 63920 2864
rect 66720 2916 66772 2922
rect 66720 2858 66772 2864
rect 47952 2848 48004 2854
rect 47952 2790 48004 2796
rect 47964 2446 47992 2790
rect 63880 2446 63908 2858
rect 79336 2446 79364 2926
rect 81915 2923 82235 2947
rect 82452 2984 82504 2990
rect 82452 2926 82504 2932
rect 81915 2867 81927 2923
rect 81983 2867 82007 2923
rect 82063 2867 82087 2923
rect 82143 2867 82167 2923
rect 82223 2867 82235 2923
rect 81915 2843 82235 2867
rect 81915 2787 81927 2843
rect 81983 2787 82007 2843
rect 82063 2787 82087 2843
rect 82143 2787 82167 2843
rect 82223 2787 82235 2843
rect 81915 2763 82235 2787
rect 81915 2746 81927 2763
rect 81983 2746 82007 2763
rect 82063 2746 82087 2763
rect 82143 2746 82167 2763
rect 82223 2746 82235 2763
rect 81915 2694 81921 2746
rect 81983 2707 81985 2746
rect 82165 2707 82167 2746
rect 81973 2694 81985 2707
rect 82037 2694 82049 2707
rect 82101 2694 82113 2707
rect 82165 2694 82177 2707
rect 82229 2694 82235 2746
rect 32496 2440 32548 2446
rect 32496 2382 32548 2388
rect 47952 2440 48004 2446
rect 47952 2382 48004 2388
rect 63868 2440 63920 2446
rect 63868 2382 63920 2388
rect 79324 2440 79376 2446
rect 79324 2382 79376 2388
rect 17868 2372 17920 2378
rect 17868 2314 17920 2320
rect 20996 2372 21048 2378
rect 20996 2314 21048 2320
rect 15936 2304 15988 2310
rect 15936 2246 15988 2252
rect 31668 2304 31720 2310
rect 31668 2246 31720 2252
rect 15948 814 15976 2246
rect 31680 814 31708 2246
rect 47964 814 47992 2382
rect 62028 2304 62080 2310
rect 62028 2246 62080 2252
rect 77208 2304 77260 2310
rect 77208 2246 77260 2252
rect 62040 814 62068 2246
rect 77220 814 77248 2246
rect 81915 964 82235 2694
rect 81915 908 81927 964
rect 81983 908 82007 964
rect 82063 908 82087 964
rect 82143 908 82167 964
rect 82223 908 82235 964
rect 81915 884 82235 908
rect 81915 828 81927 884
rect 81983 828 82007 884
rect 82063 828 82087 884
rect 82143 828 82167 884
rect 82223 828 82235 884
rect -416 748 -404 804
rect -348 748 -324 804
rect -268 748 -244 804
rect -188 748 -164 804
rect -108 748 -96 804
rect 1584 808 1636 814
rect 1584 750 1636 756
rect 15936 808 15988 814
rect 15936 750 15988 756
rect 31668 808 31720 814
rect 31668 750 31720 756
rect 47952 808 48004 814
rect 47952 750 48004 756
rect 62028 808 62080 814
rect 62028 750 62080 756
rect 77208 808 77260 814
rect 77208 750 77260 756
rect 81915 804 82235 828
rect -416 724 -96 748
rect -416 668 -404 724
rect -348 668 -324 724
rect -268 668 -244 724
rect -188 668 -164 724
rect -108 668 -96 724
rect -416 656 -96 668
rect 81915 748 81927 804
rect 81983 748 82007 804
rect 82063 748 82087 804
rect 82143 748 82167 804
rect 82223 748 82235 804
rect 81915 724 82235 748
rect 81915 668 81927 724
rect 81983 668 82007 724
rect 82063 668 82087 724
rect 82143 668 82167 724
rect 82223 668 82235 724
rect -1076 248 -1064 304
rect -1008 248 -984 304
rect -928 248 -904 304
rect -848 248 -824 304
rect -768 248 -756 304
rect -1076 224 -756 248
rect -1076 168 -1064 224
rect -1008 168 -984 224
rect -928 168 -904 224
rect -848 168 -824 224
rect -768 168 -756 224
rect -1076 144 -756 168
rect -1076 88 -1064 144
rect -1008 88 -984 144
rect -928 88 -904 144
rect -848 88 -824 144
rect -768 88 -756 144
rect -1076 64 -756 88
rect -1076 8 -1064 64
rect -1008 8 -984 64
rect -928 8 -904 64
rect -848 8 -824 64
rect -768 8 -756 64
rect -1076 -4 -756 8
rect 81915 -4 82235 668
rect 82575 2202 82895 3238
rect 112364 3194 112392 6190
rect 116136 5914 116164 6666
rect 117424 6662 117452 6718
rect 117976 6662 118004 7346
rect 118988 7342 119016 9114
rect 243858 9068 243870 9124
rect 243926 9068 243950 9124
rect 244006 9068 244030 9124
rect 244086 9068 244110 9124
rect 244166 9068 244178 9124
rect 243858 9044 244178 9068
rect 243858 8988 243870 9044
rect 243926 8988 243950 9044
rect 244006 8988 244030 9044
rect 244086 8988 244110 9044
rect 244166 8988 244178 9044
rect 243858 8964 244178 8988
rect 243858 8908 243870 8964
rect 243926 8908 243950 8964
rect 244006 8908 244030 8964
rect 244086 8908 244110 8964
rect 244166 8908 244178 8964
rect 243858 8884 244178 8908
rect 243858 8828 243870 8884
rect 243926 8828 243950 8884
rect 244006 8828 244030 8884
rect 244086 8828 244110 8884
rect 244166 8828 244178 8884
rect 123852 8424 123904 8430
rect 123852 8366 123904 8372
rect 121458 8120 121514 8129
rect 121458 8055 121514 8064
rect 121472 7410 121500 8055
rect 122838 7984 122894 7993
rect 122838 7919 122894 7928
rect 122852 7410 122880 7919
rect 123208 7540 123260 7546
rect 123208 7482 123260 7488
rect 123220 7410 123248 7482
rect 123864 7410 123892 8366
rect 151176 8288 151228 8294
rect 151176 8230 151228 8236
rect 125324 7880 125376 7886
rect 125324 7822 125376 7828
rect 125336 7410 125364 7822
rect 151188 7410 151216 8230
rect 168196 8220 168248 8226
rect 168196 8162 168248 8168
rect 166448 8152 166500 8158
rect 166448 8094 166500 8100
rect 166460 7410 166488 8094
rect 168208 7410 168236 8162
rect 170128 7948 170180 7954
rect 170128 7890 170180 7896
rect 170140 7410 170168 7890
rect 200120 7812 200172 7818
rect 200120 7754 200172 7760
rect 197912 7744 197964 7750
rect 197912 7686 197964 7692
rect 197924 7410 197952 7686
rect 200132 7410 200160 7754
rect 119344 7404 119396 7410
rect 119344 7346 119396 7352
rect 121460 7404 121512 7410
rect 121460 7346 121512 7352
rect 121828 7404 121880 7410
rect 121828 7346 121880 7352
rect 122840 7404 122892 7410
rect 122840 7346 122892 7352
rect 123208 7404 123260 7410
rect 123208 7346 123260 7352
rect 123852 7404 123904 7410
rect 123852 7346 123904 7352
rect 125324 7404 125376 7410
rect 125324 7346 125376 7352
rect 151176 7404 151228 7410
rect 151176 7346 151228 7352
rect 152740 7404 152792 7410
rect 152740 7346 152792 7352
rect 166448 7404 166500 7410
rect 166448 7346 166500 7352
rect 168196 7404 168248 7410
rect 168196 7346 168248 7352
rect 170128 7404 170180 7410
rect 170128 7346 170180 7352
rect 197912 7404 197964 7410
rect 197912 7346 197964 7352
rect 200120 7404 200172 7410
rect 200120 7346 200172 7352
rect 217876 7404 217928 7410
rect 217876 7346 217928 7352
rect 220452 7404 220504 7410
rect 220452 7346 220504 7352
rect 118976 7336 119028 7342
rect 118976 7278 119028 7284
rect 118988 6934 119016 7278
rect 118976 6928 119028 6934
rect 118976 6870 119028 6876
rect 117412 6656 117464 6662
rect 117412 6598 117464 6604
rect 117964 6656 118016 6662
rect 117964 6598 118016 6604
rect 116124 5908 116176 5914
rect 116124 5850 116176 5856
rect 115664 5704 115716 5710
rect 115664 5646 115716 5652
rect 114468 4616 114520 4622
rect 114468 4558 114520 4564
rect 112352 3188 112404 3194
rect 112352 3130 112404 3136
rect 110236 3120 110288 3126
rect 110236 3062 110288 3068
rect 94320 2848 94372 2854
rect 94320 2790 94372 2796
rect 94332 2446 94360 2790
rect 110248 2446 110276 3062
rect 94320 2440 94372 2446
rect 94320 2382 94372 2388
rect 110236 2440 110288 2446
rect 110236 2382 110288 2388
rect 82575 2150 82581 2202
rect 82633 2150 82645 2202
rect 82697 2150 82709 2202
rect 82761 2150 82773 2202
rect 82825 2150 82837 2202
rect 82889 2150 82895 2202
rect 82575 304 82895 2150
rect 94332 814 94360 2382
rect 114480 2378 114508 4558
rect 115676 2514 115704 5646
rect 117424 3466 117452 6598
rect 117976 4554 118004 6598
rect 119356 6118 119384 7346
rect 120448 6792 120500 6798
rect 120448 6734 120500 6740
rect 121460 6792 121512 6798
rect 121460 6734 121512 6740
rect 120460 6118 120488 6734
rect 120816 6724 120868 6730
rect 120816 6666 120868 6672
rect 120828 6322 120856 6666
rect 120816 6316 120868 6322
rect 120816 6258 120868 6264
rect 121472 6118 121500 6734
rect 121840 6118 121868 7346
rect 123220 6934 123248 7346
rect 123208 6928 123260 6934
rect 123208 6870 123260 6876
rect 123864 6390 123892 7346
rect 125508 7336 125560 7342
rect 125508 7278 125560 7284
rect 126520 7336 126572 7342
rect 126520 7278 126572 7284
rect 124036 6792 124088 6798
rect 124036 6734 124088 6740
rect 124048 6390 124076 6734
rect 124680 6724 124732 6730
rect 124680 6666 124732 6672
rect 124692 6633 124720 6666
rect 125520 6633 125548 7278
rect 124678 6624 124734 6633
rect 124678 6559 124734 6568
rect 125506 6624 125562 6633
rect 125506 6559 125562 6568
rect 123852 6384 123904 6390
rect 123852 6326 123904 6332
rect 124036 6384 124088 6390
rect 124036 6326 124088 6332
rect 122564 6316 122616 6322
rect 122564 6258 122616 6264
rect 119344 6112 119396 6118
rect 119344 6054 119396 6060
rect 120448 6112 120500 6118
rect 120448 6054 120500 6060
rect 121460 6112 121512 6118
rect 121460 6054 121512 6060
rect 121828 6112 121880 6118
rect 121828 6054 121880 6060
rect 119356 5642 119384 6054
rect 120460 5914 120488 6054
rect 120448 5908 120500 5914
rect 120448 5850 120500 5856
rect 121472 5846 121500 6054
rect 121460 5840 121512 5846
rect 121460 5782 121512 5788
rect 119344 5636 119396 5642
rect 119344 5578 119396 5584
rect 122576 5574 122604 6258
rect 122564 5568 122616 5574
rect 122564 5510 122616 5516
rect 126532 5030 126560 7278
rect 151188 6934 151216 7346
rect 151728 7336 151780 7342
rect 151728 7278 151780 7284
rect 151740 6934 151768 7278
rect 152752 7206 152780 7346
rect 154488 7336 154540 7342
rect 154488 7278 154540 7284
rect 157340 7336 157392 7342
rect 157340 7278 157392 7284
rect 152740 7200 152792 7206
rect 152740 7142 152792 7148
rect 152752 7002 152780 7142
rect 152740 6996 152792 7002
rect 152740 6938 152792 6944
rect 151176 6928 151228 6934
rect 151176 6870 151228 6876
rect 151728 6928 151780 6934
rect 151728 6870 151780 6876
rect 154500 6633 154528 7278
rect 154580 7268 154632 7274
rect 154580 7210 154632 7216
rect 154592 6934 154620 7210
rect 154580 6928 154632 6934
rect 154580 6870 154632 6876
rect 155776 6792 155828 6798
rect 155776 6734 155828 6740
rect 155788 6662 155816 6734
rect 156972 6724 157024 6730
rect 156972 6666 157024 6672
rect 155776 6656 155828 6662
rect 154302 6624 154358 6633
rect 154302 6559 154358 6568
rect 154486 6624 154542 6633
rect 155776 6598 155828 6604
rect 154486 6559 154542 6568
rect 126888 6316 126940 6322
rect 126888 6258 126940 6264
rect 126900 6186 126928 6258
rect 127532 6248 127584 6254
rect 127532 6190 127584 6196
rect 127624 6248 127676 6254
rect 127624 6190 127676 6196
rect 126888 6180 126940 6186
rect 126888 6122 126940 6128
rect 126980 6180 127032 6186
rect 126980 6122 127032 6128
rect 126992 5953 127020 6122
rect 126978 5944 127034 5953
rect 126978 5879 127034 5888
rect 126520 5024 126572 5030
rect 126520 4966 126572 4972
rect 117964 4548 118016 4554
rect 117964 4490 118016 4496
rect 117412 3460 117464 3466
rect 117412 3402 117464 3408
rect 127544 3058 127572 6190
rect 127636 5642 127664 6190
rect 154316 5953 154344 6559
rect 155788 6458 155816 6598
rect 155776 6452 155828 6458
rect 155776 6394 155828 6400
rect 154302 5944 154358 5953
rect 154302 5879 154358 5888
rect 127624 5636 127676 5642
rect 127624 5578 127676 5584
rect 156984 4690 157012 6666
rect 157352 6458 157380 7278
rect 166460 7002 166488 7346
rect 169484 7336 169536 7342
rect 169484 7278 169536 7284
rect 166448 6996 166500 7002
rect 166448 6938 166500 6944
rect 169496 6458 169524 7278
rect 170140 7002 170168 7346
rect 170680 7336 170732 7342
rect 170680 7278 170732 7284
rect 199108 7336 199160 7342
rect 199108 7278 199160 7284
rect 201316 7336 201368 7342
rect 201316 7278 201368 7284
rect 214564 7336 214616 7342
rect 214564 7278 214616 7284
rect 214748 7336 214800 7342
rect 214748 7278 214800 7284
rect 170128 6996 170180 7002
rect 170128 6938 170180 6944
rect 170220 6996 170272 7002
rect 170220 6938 170272 6944
rect 170232 6866 170260 6938
rect 170692 6866 170720 7278
rect 172336 6996 172388 7002
rect 172336 6938 172388 6944
rect 170220 6860 170272 6866
rect 170220 6802 170272 6808
rect 170680 6860 170732 6866
rect 170680 6802 170732 6808
rect 171048 6792 171100 6798
rect 171048 6734 171100 6740
rect 171060 6662 171088 6734
rect 172348 6730 172376 6938
rect 173072 6792 173124 6798
rect 173072 6734 173124 6740
rect 172244 6724 172296 6730
rect 172244 6666 172296 6672
rect 172336 6724 172388 6730
rect 172336 6666 172388 6672
rect 171048 6656 171100 6662
rect 171048 6598 171100 6604
rect 157340 6452 157392 6458
rect 157340 6394 157392 6400
rect 167184 6452 167236 6458
rect 167184 6394 167236 6400
rect 169484 6452 169536 6458
rect 169484 6394 169536 6400
rect 167196 5953 167224 6394
rect 171060 6186 171088 6598
rect 171048 6180 171100 6186
rect 171048 6122 171100 6128
rect 166998 5944 167054 5953
rect 166998 5879 167054 5888
rect 167182 5944 167238 5953
rect 167182 5879 167238 5888
rect 167012 5642 167040 5879
rect 157892 5636 157944 5642
rect 157892 5578 157944 5584
rect 167000 5636 167052 5642
rect 167000 5578 167052 5584
rect 156972 4684 157024 4690
rect 156972 4626 157024 4632
rect 125232 3052 125284 3058
rect 125232 2994 125284 3000
rect 127532 3052 127584 3058
rect 127532 2994 127584 3000
rect 115664 2508 115716 2514
rect 115664 2450 115716 2456
rect 125244 2446 125272 2994
rect 157904 2922 157932 5578
rect 172256 4758 172284 6666
rect 173084 6458 173112 6734
rect 190552 6656 190604 6662
rect 190552 6598 190604 6604
rect 190644 6656 190696 6662
rect 190644 6598 190696 6604
rect 173072 6452 173124 6458
rect 173072 6394 173124 6400
rect 173164 6452 173216 6458
rect 173164 6394 173216 6400
rect 173176 5642 173204 6394
rect 190564 6338 190592 6598
rect 190656 6458 190684 6598
rect 190644 6452 190696 6458
rect 190644 6394 190696 6400
rect 190736 6452 190788 6458
rect 190736 6394 190788 6400
rect 190748 6338 190776 6394
rect 190564 6310 190776 6338
rect 199120 5778 199148 7278
rect 200580 6452 200632 6458
rect 200580 6394 200632 6400
rect 200592 6254 200620 6394
rect 200580 6248 200632 6254
rect 200580 6190 200632 6196
rect 199108 5772 199160 5778
rect 199108 5714 199160 5720
rect 201328 5710 201356 7278
rect 213276 6656 213328 6662
rect 213276 6598 213328 6604
rect 213368 6656 213420 6662
rect 213368 6598 213420 6604
rect 213288 6254 213316 6598
rect 213380 6322 213408 6598
rect 214576 6458 214604 7278
rect 214760 6730 214788 7278
rect 217888 7206 217916 7346
rect 220464 7206 220492 7346
rect 217876 7200 217928 7206
rect 217876 7142 217928 7148
rect 220452 7200 220504 7206
rect 220452 7142 220504 7148
rect 215300 6996 215352 7002
rect 215300 6938 215352 6944
rect 215772 6990 216260 7018
rect 215312 6798 215340 6938
rect 215772 6866 215800 6990
rect 215852 6928 215904 6934
rect 216036 6928 216088 6934
rect 215904 6876 216036 6882
rect 215852 6870 216088 6876
rect 215760 6860 215812 6866
rect 215864 6854 216076 6870
rect 216232 6866 216260 6990
rect 216220 6860 216272 6866
rect 215760 6802 215812 6808
rect 216220 6802 216272 6808
rect 215300 6792 215352 6798
rect 215300 6734 215352 6740
rect 214748 6724 214800 6730
rect 214748 6666 214800 6672
rect 216588 6724 216640 6730
rect 216588 6666 216640 6672
rect 217508 6724 217560 6730
rect 217508 6666 217560 6672
rect 214564 6452 214616 6458
rect 214564 6394 214616 6400
rect 214944 6322 215340 6338
rect 213368 6316 213420 6322
rect 213368 6258 213420 6264
rect 213644 6316 213696 6322
rect 213644 6258 213696 6264
rect 214932 6316 215340 6322
rect 214984 6310 215340 6316
rect 214932 6258 214984 6264
rect 202788 6248 202840 6254
rect 202788 6190 202840 6196
rect 211528 6248 211580 6254
rect 211528 6190 211580 6196
rect 212908 6248 212960 6254
rect 212908 6190 212960 6196
rect 213276 6248 213328 6254
rect 213276 6190 213328 6196
rect 213656 6202 213684 6258
rect 214104 6248 214156 6254
rect 201316 5704 201368 5710
rect 201316 5646 201368 5652
rect 173164 5636 173216 5642
rect 173164 5578 173216 5584
rect 173256 5636 173308 5642
rect 173256 5578 173308 5584
rect 172244 4752 172296 4758
rect 172244 4694 172296 4700
rect 173268 3126 173296 5578
rect 202800 4486 202828 6190
rect 203156 6180 203208 6186
rect 203156 6122 203208 6128
rect 203168 5778 203196 6122
rect 203156 5772 203208 5778
rect 203156 5714 203208 5720
rect 211540 5710 211568 6190
rect 212920 5914 212948 6190
rect 213656 6174 213776 6202
rect 215116 6248 215168 6254
rect 214104 6190 214156 6196
rect 214944 6196 215116 6202
rect 214944 6190 215168 6196
rect 212908 5908 212960 5914
rect 212908 5850 212960 5856
rect 211528 5704 211580 5710
rect 211528 5646 211580 5652
rect 213748 5574 213776 6174
rect 214116 5846 214144 6190
rect 214944 6174 215156 6190
rect 214944 6118 214972 6174
rect 214932 6112 214984 6118
rect 214932 6054 214984 6060
rect 214104 5840 214156 5846
rect 214104 5782 214156 5788
rect 215312 5574 215340 6310
rect 216496 6316 216548 6322
rect 216496 6258 216548 6264
rect 216508 6118 216536 6258
rect 216496 6112 216548 6118
rect 216496 6054 216548 6060
rect 212724 5568 212776 5574
rect 212724 5510 212776 5516
rect 213736 5568 213788 5574
rect 213736 5510 213788 5516
rect 215300 5568 215352 5574
rect 215300 5510 215352 5516
rect 203892 5160 203944 5166
rect 203892 5102 203944 5108
rect 202788 4480 202840 4486
rect 202788 4422 202840 4428
rect 203904 3194 203932 5102
rect 211344 4616 211396 4622
rect 211344 4558 211396 4564
rect 211356 4486 211384 4558
rect 211344 4480 211396 4486
rect 211344 4422 211396 4428
rect 202512 3188 202564 3194
rect 202512 3130 202564 3136
rect 203892 3188 203944 3194
rect 203892 3130 203944 3136
rect 173256 3120 173308 3126
rect 173256 3062 173308 3068
rect 172060 2984 172112 2990
rect 172060 2926 172112 2932
rect 156604 2916 156656 2922
rect 156604 2858 156656 2864
rect 157892 2916 157944 2922
rect 157892 2858 157944 2864
rect 141056 2848 141108 2854
rect 141056 2790 141108 2796
rect 125232 2440 125284 2446
rect 125232 2382 125284 2388
rect 141068 2378 141096 2790
rect 156616 2446 156644 2858
rect 172072 2446 172100 2926
rect 186872 2848 186924 2854
rect 186872 2790 186924 2796
rect 156604 2440 156656 2446
rect 156604 2382 156656 2388
rect 172060 2440 172112 2446
rect 172060 2382 172112 2388
rect 186884 2378 186912 2790
rect 202524 2446 202552 3130
rect 211356 2514 211384 4422
rect 212736 2990 212764 5510
rect 213748 4010 213776 5510
rect 215312 4554 215340 5510
rect 216508 5302 216536 6054
rect 216496 5296 216548 5302
rect 216496 5238 216548 5244
rect 216600 4622 216628 6666
rect 217520 6390 217548 6666
rect 217508 6384 217560 6390
rect 217508 6326 217560 6332
rect 217888 5846 217916 7142
rect 218796 6996 218848 7002
rect 218796 6938 218848 6944
rect 218808 6798 218836 6938
rect 218796 6792 218848 6798
rect 218796 6734 218848 6740
rect 220464 6322 220492 7142
rect 243858 7098 244178 8828
rect 244518 9784 244838 9796
rect 244518 9728 244530 9784
rect 244586 9728 244610 9784
rect 244666 9728 244690 9784
rect 244746 9728 244770 9784
rect 244826 9728 244838 9784
rect 244518 9704 244838 9728
rect 244518 9648 244530 9704
rect 244586 9648 244610 9704
rect 244666 9648 244690 9704
rect 244746 9648 244770 9704
rect 244826 9648 244838 9704
rect 244518 9624 244838 9648
rect 244518 9568 244530 9624
rect 244586 9568 244610 9624
rect 244666 9568 244690 9624
rect 244746 9568 244770 9624
rect 244826 9568 244838 9624
rect 244518 9544 244838 9568
rect 244518 9488 244530 9544
rect 244586 9488 244610 9544
rect 244666 9488 244690 9544
rect 244746 9488 244770 9544
rect 244826 9488 244838 9544
rect 244518 7740 244838 9488
rect 244518 7684 244530 7740
rect 244586 7684 244610 7740
rect 244666 7684 244690 7740
rect 244746 7684 244770 7740
rect 244826 7684 244838 7740
rect 244518 7660 244838 7684
rect 244518 7642 244530 7660
rect 244586 7642 244610 7660
rect 244666 7642 244690 7660
rect 244746 7642 244770 7660
rect 244826 7642 244838 7660
rect 244518 7590 244524 7642
rect 244586 7604 244588 7642
rect 244768 7604 244770 7642
rect 244576 7590 244588 7604
rect 244640 7590 244652 7604
rect 244704 7590 244716 7604
rect 244768 7590 244780 7604
rect 244832 7590 244838 7642
rect 244518 7580 244838 7590
rect 244518 7524 244530 7580
rect 244586 7524 244610 7580
rect 244666 7524 244690 7580
rect 244746 7524 244770 7580
rect 244826 7524 244838 7580
rect 244518 7500 244838 7524
rect 244518 7444 244530 7500
rect 244586 7444 244610 7500
rect 244666 7444 244690 7500
rect 244746 7444 244770 7500
rect 244826 7444 244838 7500
rect 244372 7404 244424 7410
rect 244372 7346 244424 7352
rect 243858 7046 243864 7098
rect 243916 7080 243928 7098
rect 243980 7080 243992 7098
rect 244044 7080 244056 7098
rect 244108 7080 244120 7098
rect 243926 7046 243928 7080
rect 244108 7046 244110 7080
rect 244172 7046 244178 7098
rect 243858 7024 243870 7046
rect 243926 7024 243950 7046
rect 244006 7024 244030 7046
rect 244086 7024 244110 7046
rect 244166 7024 244178 7046
rect 243858 7000 244178 7024
rect 243858 6944 243870 7000
rect 243926 6944 243950 7000
rect 244006 6944 244030 7000
rect 244086 6944 244110 7000
rect 244166 6944 244178 7000
rect 243858 6920 244178 6944
rect 244384 6934 244412 7346
rect 243858 6864 243870 6920
rect 243926 6864 243950 6920
rect 244006 6864 244030 6920
rect 244086 6864 244110 6920
rect 244166 6864 244178 6920
rect 244372 6928 244424 6934
rect 244372 6870 244424 6876
rect 243858 6840 244178 6864
rect 243858 6784 243870 6840
rect 243926 6784 243950 6840
rect 244006 6784 244030 6840
rect 244086 6784 244110 6840
rect 244166 6784 244178 6840
rect 220452 6316 220504 6322
rect 220452 6258 220504 6264
rect 218428 6248 218480 6254
rect 218428 6190 218480 6196
rect 217876 5840 217928 5846
rect 217876 5782 217928 5788
rect 216588 4616 216640 4622
rect 216588 4558 216640 4564
rect 215300 4548 215352 4554
rect 215300 4490 215352 4496
rect 218440 4214 218468 6190
rect 243858 6010 244178 6784
rect 243858 5958 243864 6010
rect 243916 5958 243928 6010
rect 243980 5958 243992 6010
rect 244044 5958 244056 6010
rect 244108 5958 244120 6010
rect 244172 5958 244178 6010
rect 243858 5721 244178 5958
rect 243858 5665 243870 5721
rect 243926 5665 243950 5721
rect 244006 5665 244030 5721
rect 244086 5665 244110 5721
rect 244166 5665 244178 5721
rect 243858 5641 244178 5665
rect 243858 5585 243870 5641
rect 243926 5585 243950 5641
rect 244006 5585 244030 5641
rect 244086 5585 244110 5641
rect 244166 5585 244178 5641
rect 243858 5561 244178 5585
rect 243858 5505 243870 5561
rect 243926 5505 243950 5561
rect 244006 5505 244030 5561
rect 244086 5505 244110 5561
rect 244166 5505 244178 5561
rect 243858 5481 244178 5505
rect 243858 5425 243870 5481
rect 243926 5425 243950 5481
rect 244006 5425 244030 5481
rect 244086 5425 244110 5481
rect 244166 5425 244178 5481
rect 219164 5160 219216 5166
rect 219164 5102 219216 5108
rect 218428 4208 218480 4214
rect 218428 4150 218480 4156
rect 213736 4004 213788 4010
rect 213736 3946 213788 3952
rect 219176 3058 219204 5102
rect 243858 4922 244178 5425
rect 243858 4870 243864 4922
rect 243916 4870 243928 4922
rect 243980 4870 243992 4922
rect 244044 4870 244056 4922
rect 244108 4870 244120 4922
rect 244172 4870 244178 4922
rect 233884 4820 233936 4826
rect 233884 4762 233936 4768
rect 233896 4690 233924 4762
rect 239312 4752 239364 4758
rect 239496 4752 239548 4758
rect 239364 4700 239496 4706
rect 239312 4694 239548 4700
rect 233884 4684 233936 4690
rect 239324 4678 239536 4694
rect 233884 4626 233936 4632
rect 239404 4548 239456 4554
rect 239404 4490 239456 4496
rect 239416 4434 239444 4490
rect 239588 4480 239640 4486
rect 239416 4428 239588 4434
rect 239416 4422 239640 4428
rect 239416 4406 239628 4422
rect 243858 4362 244178 4870
rect 243858 4306 243870 4362
rect 243926 4306 243950 4362
rect 244006 4306 244030 4362
rect 244086 4306 244110 4362
rect 244166 4306 244178 4362
rect 243858 4282 244178 4306
rect 243858 4226 243870 4282
rect 243926 4226 243950 4282
rect 244006 4226 244030 4282
rect 244086 4226 244110 4282
rect 244166 4226 244178 4282
rect 243858 4202 244178 4226
rect 243858 4146 243870 4202
rect 243926 4146 243950 4202
rect 244006 4146 244030 4202
rect 244086 4146 244110 4202
rect 244166 4146 244178 4202
rect 243858 4122 244178 4146
rect 243858 4066 243870 4122
rect 243926 4066 243950 4122
rect 244006 4066 244030 4122
rect 244086 4066 244110 4122
rect 244166 4066 244178 4122
rect 243858 3834 244178 4066
rect 243858 3782 243864 3834
rect 243916 3782 243928 3834
rect 243980 3782 243992 3834
rect 244044 3782 244056 3834
rect 244108 3782 244120 3834
rect 244172 3782 244178 3834
rect 233608 3528 233660 3534
rect 233608 3470 233660 3476
rect 218428 3052 218480 3058
rect 218428 2994 218480 3000
rect 219164 3052 219216 3058
rect 219164 2994 219216 3000
rect 212724 2984 212776 2990
rect 212724 2926 212776 2932
rect 211344 2508 211396 2514
rect 211344 2450 211396 2456
rect 218440 2446 218468 2994
rect 233620 2582 233648 3470
rect 243858 3003 244178 3782
rect 243858 2947 243870 3003
rect 243926 2947 243950 3003
rect 244006 2947 244030 3003
rect 244086 2947 244110 3003
rect 244166 2947 244178 3003
rect 243858 2923 244178 2947
rect 243858 2867 243870 2923
rect 243926 2867 243950 2923
rect 244006 2867 244030 2923
rect 244086 2867 244110 2923
rect 244166 2867 244178 2923
rect 233792 2848 233844 2854
rect 233792 2790 233844 2796
rect 243858 2843 244178 2867
rect 233608 2576 233660 2582
rect 233608 2518 233660 2524
rect 202512 2440 202564 2446
rect 202512 2382 202564 2388
rect 218428 2440 218480 2446
rect 218428 2382 218480 2388
rect 233804 2378 233832 2790
rect 243858 2787 243870 2843
rect 243926 2787 243950 2843
rect 244006 2787 244030 2843
rect 244086 2787 244110 2843
rect 244166 2787 244178 2843
rect 243858 2763 244178 2787
rect 243858 2746 243870 2763
rect 243926 2746 243950 2763
rect 244006 2746 244030 2763
rect 244086 2746 244110 2763
rect 244166 2746 244178 2763
rect 243858 2694 243864 2746
rect 243926 2707 243928 2746
rect 244108 2707 244110 2746
rect 243916 2694 243928 2707
rect 243980 2694 243992 2707
rect 244044 2694 244056 2707
rect 244108 2694 244120 2707
rect 244172 2694 244178 2746
rect 114468 2372 114520 2378
rect 114468 2314 114520 2320
rect 141056 2372 141108 2378
rect 141056 2314 141108 2320
rect 186872 2372 186924 2378
rect 186872 2314 186924 2320
rect 233792 2372 233844 2378
rect 233792 2314 233844 2320
rect 107568 2304 107620 2310
rect 107568 2246 107620 2252
rect 122656 2304 122708 2310
rect 122656 2246 122708 2252
rect 107580 814 107608 2246
rect 122668 814 122696 2246
rect 141068 814 141096 2314
rect 156420 2304 156472 2310
rect 156420 2246 156472 2252
rect 169668 2304 169720 2310
rect 169668 2246 169720 2252
rect 156432 814 156460 2246
rect 169680 814 169708 2246
rect 186884 814 186912 2314
rect 199476 2304 199528 2310
rect 199476 2246 199528 2252
rect 218244 2304 218296 2310
rect 218244 2246 218296 2252
rect 199488 814 199516 2246
rect 218256 814 218284 2246
rect 233804 814 233832 2314
rect 243858 964 244178 2694
rect 243858 908 243870 964
rect 243926 908 243950 964
rect 244006 908 244030 964
rect 244086 908 244110 964
rect 244166 908 244178 964
rect 243858 884 244178 908
rect 243858 828 243870 884
rect 243926 828 243950 884
rect 244006 828 244030 884
rect 244086 828 244110 884
rect 244166 828 244178 884
rect 94320 808 94372 814
rect 94320 750 94372 756
rect 107568 808 107620 814
rect 107568 750 107620 756
rect 122656 808 122708 814
rect 122656 750 122708 756
rect 141056 808 141108 814
rect 141056 750 141108 756
rect 156420 808 156472 814
rect 156420 750 156472 756
rect 169668 808 169720 814
rect 169668 750 169720 756
rect 186872 808 186924 814
rect 186872 750 186924 756
rect 199476 808 199528 814
rect 199476 750 199528 756
rect 218244 808 218296 814
rect 218244 750 218296 756
rect 233792 808 233844 814
rect 233792 750 233844 756
rect 243858 804 244178 828
rect 82575 248 82587 304
rect 82643 248 82667 304
rect 82723 248 82747 304
rect 82803 248 82827 304
rect 82883 248 82895 304
rect 82575 224 82895 248
rect 82575 168 82587 224
rect 82643 168 82667 224
rect 82723 168 82747 224
rect 82803 168 82827 224
rect 82883 168 82895 224
rect 82575 144 82895 168
rect 82575 88 82587 144
rect 82643 88 82667 144
rect 82723 88 82747 144
rect 82803 88 82827 144
rect 82883 88 82895 144
rect 82575 64 82895 88
rect 82575 8 82587 64
rect 82643 8 82667 64
rect 82723 8 82747 64
rect 82803 8 82827 64
rect 82883 8 82895 64
rect 82575 -4 82895 8
rect 243858 748 243870 804
rect 243926 748 243950 804
rect 244006 748 244030 804
rect 244086 748 244110 804
rect 244166 748 244178 804
rect 243858 724 244178 748
rect 243858 668 243870 724
rect 243926 668 243950 724
rect 244006 668 244030 724
rect 244086 668 244110 724
rect 244166 668 244178 724
rect 243858 -4 244178 668
rect 244518 6554 244838 7444
rect 405801 9124 406121 9796
rect 405801 9068 405813 9124
rect 405869 9068 405893 9124
rect 405949 9068 405973 9124
rect 406029 9068 406053 9124
rect 406109 9068 406121 9124
rect 405801 9044 406121 9068
rect 405801 8988 405813 9044
rect 405869 8988 405893 9044
rect 405949 8988 405973 9044
rect 406029 8988 406053 9044
rect 406109 8988 406121 9044
rect 405801 8964 406121 8988
rect 405801 8908 405813 8964
rect 405869 8908 405893 8964
rect 405949 8908 405973 8964
rect 406029 8908 406053 8964
rect 406109 8908 406121 8964
rect 405801 8884 406121 8908
rect 405801 8828 405813 8884
rect 405869 8828 405893 8884
rect 405949 8828 405973 8884
rect 406029 8828 406053 8884
rect 406109 8828 406121 8884
rect 245476 7336 245528 7342
rect 245476 7278 245528 7284
rect 260748 7336 260800 7342
rect 260748 7278 260800 7284
rect 244518 6502 244524 6554
rect 244576 6502 244588 6554
rect 244640 6502 244652 6554
rect 244704 6502 244716 6554
rect 244768 6502 244780 6554
rect 244832 6502 244838 6554
rect 244518 6381 244838 6502
rect 244518 6325 244530 6381
rect 244586 6325 244610 6381
rect 244666 6325 244690 6381
rect 244746 6325 244770 6381
rect 244826 6325 244838 6381
rect 244518 6301 244838 6325
rect 244518 6245 244530 6301
rect 244586 6245 244610 6301
rect 244666 6245 244690 6301
rect 244746 6245 244770 6301
rect 244826 6245 244838 6301
rect 244518 6221 244838 6245
rect 244518 6165 244530 6221
rect 244586 6165 244610 6221
rect 244666 6165 244690 6221
rect 244746 6165 244770 6221
rect 244826 6165 244838 6221
rect 244518 6141 244838 6165
rect 244518 6085 244530 6141
rect 244586 6085 244610 6141
rect 244666 6085 244690 6141
rect 244746 6085 244770 6141
rect 244826 6085 244838 6141
rect 244518 5466 244838 6085
rect 245488 5914 245516 7278
rect 246764 6792 246816 6798
rect 246764 6734 246816 6740
rect 246120 6656 246172 6662
rect 246118 6624 246120 6633
rect 246776 6633 246804 6734
rect 247316 6724 247368 6730
rect 247316 6666 247368 6672
rect 246172 6624 246174 6633
rect 246118 6559 246174 6568
rect 246762 6624 246818 6633
rect 246762 6559 246818 6568
rect 245476 5908 245528 5914
rect 245476 5850 245528 5856
rect 244518 5414 244524 5466
rect 244576 5414 244588 5466
rect 244640 5414 244652 5466
rect 244704 5414 244716 5466
rect 244768 5414 244780 5466
rect 244832 5414 244838 5466
rect 244518 5022 244838 5414
rect 247328 5030 247356 6666
rect 260760 6390 260788 7278
rect 405801 7098 406121 8828
rect 405801 7046 405807 7098
rect 405859 7080 405871 7098
rect 405923 7080 405935 7098
rect 405987 7080 405999 7098
rect 406051 7080 406063 7098
rect 405869 7046 405871 7080
rect 406051 7046 406053 7080
rect 406115 7046 406121 7098
rect 405801 7024 405813 7046
rect 405869 7024 405893 7046
rect 405949 7024 405973 7046
rect 406029 7024 406053 7046
rect 406109 7024 406121 7046
rect 405801 7000 406121 7024
rect 405801 6944 405813 7000
rect 405869 6944 405893 7000
rect 405949 6944 405973 7000
rect 406029 6944 406053 7000
rect 406109 6944 406121 7000
rect 405801 6920 406121 6944
rect 262956 6860 263008 6866
rect 262956 6802 263008 6808
rect 405801 6864 405813 6920
rect 405869 6864 405893 6920
rect 405949 6864 405973 6920
rect 406029 6864 406053 6920
rect 406109 6864 406121 6920
rect 405801 6840 406121 6864
rect 261760 6792 261812 6798
rect 261760 6734 261812 6740
rect 260748 6384 260800 6390
rect 260748 6326 260800 6332
rect 261772 6254 261800 6734
rect 262588 6724 262640 6730
rect 262588 6666 262640 6672
rect 261760 6248 261812 6254
rect 261760 6190 261812 6196
rect 247590 5944 247646 5953
rect 247590 5879 247646 5888
rect 247604 5710 247632 5879
rect 247592 5704 247644 5710
rect 247592 5646 247644 5652
rect 248972 5636 249024 5642
rect 248972 5578 249024 5584
rect 244518 4966 244530 5022
rect 244586 4966 244610 5022
rect 244666 4966 244690 5022
rect 244746 4966 244770 5022
rect 244826 4966 244838 5022
rect 247316 5024 247368 5030
rect 247316 4966 247368 4972
rect 244518 4942 244838 4966
rect 244518 4886 244530 4942
rect 244586 4886 244610 4942
rect 244666 4886 244690 4942
rect 244746 4886 244770 4942
rect 244826 4886 244838 4942
rect 244518 4862 244838 4886
rect 244518 4806 244530 4862
rect 244586 4806 244610 4862
rect 244666 4806 244690 4862
rect 244746 4806 244770 4862
rect 244826 4806 244838 4862
rect 244518 4782 244838 4806
rect 244518 4726 244530 4782
rect 244586 4726 244610 4782
rect 244666 4726 244690 4782
rect 244746 4726 244770 4782
rect 244826 4726 244838 4782
rect 244518 4378 244838 4726
rect 248788 4480 248840 4486
rect 248788 4422 248840 4428
rect 244518 4326 244524 4378
rect 244576 4326 244588 4378
rect 244640 4326 244652 4378
rect 244704 4326 244716 4378
rect 244768 4326 244780 4378
rect 244832 4326 244838 4378
rect 244518 3663 244838 4326
rect 248800 4282 248828 4422
rect 248788 4276 248840 4282
rect 248788 4218 248840 4224
rect 248984 4146 249012 5578
rect 262600 5302 262628 6666
rect 262968 5710 262996 6802
rect 405801 6784 405813 6840
rect 405869 6784 405893 6840
rect 405949 6784 405973 6840
rect 406029 6784 406053 6840
rect 406109 6784 406121 6840
rect 310888 6656 310940 6662
rect 310888 6598 310940 6604
rect 310900 6322 310928 6598
rect 292580 6316 292632 6322
rect 292580 6258 292632 6264
rect 292764 6316 292816 6322
rect 292764 6258 292816 6264
rect 310888 6316 310940 6322
rect 310888 6258 310940 6264
rect 311900 6316 311952 6322
rect 311900 6258 311952 6264
rect 313740 6316 313792 6322
rect 313740 6258 313792 6264
rect 292592 6202 292620 6258
rect 292592 6186 292712 6202
rect 292592 6180 292724 6186
rect 292592 6174 292672 6180
rect 292672 6122 292724 6128
rect 292776 6118 292804 6258
rect 293316 6248 293368 6254
rect 293316 6190 293368 6196
rect 308680 6248 308732 6254
rect 308680 6190 308732 6196
rect 292764 6112 292816 6118
rect 292764 6054 292816 6060
rect 262956 5704 263008 5710
rect 262956 5646 263008 5652
rect 264336 5636 264388 5642
rect 264336 5578 264388 5584
rect 262588 5296 262640 5302
rect 262588 5238 262640 5244
rect 249340 4820 249392 4826
rect 249340 4762 249392 4768
rect 249352 4622 249380 4762
rect 249340 4616 249392 4622
rect 249340 4558 249392 4564
rect 249708 4548 249760 4554
rect 249708 4490 249760 4496
rect 249800 4548 249852 4554
rect 249800 4490 249852 4496
rect 248972 4140 249024 4146
rect 248972 4082 249024 4088
rect 244518 3607 244530 3663
rect 244586 3607 244610 3663
rect 244666 3607 244690 3663
rect 244746 3607 244770 3663
rect 244826 3607 244838 3663
rect 244518 3583 244838 3607
rect 244518 3527 244530 3583
rect 244586 3527 244610 3583
rect 244666 3527 244690 3583
rect 244746 3527 244770 3583
rect 244826 3527 244838 3583
rect 244518 3503 244838 3527
rect 244518 3447 244530 3503
rect 244586 3447 244610 3503
rect 244666 3447 244690 3503
rect 244746 3447 244770 3503
rect 244826 3447 244838 3503
rect 244518 3423 244838 3447
rect 244518 3367 244530 3423
rect 244586 3367 244610 3423
rect 244666 3367 244690 3423
rect 244746 3367 244770 3423
rect 244826 3367 244838 3423
rect 244518 3290 244838 3367
rect 244518 3238 244524 3290
rect 244576 3238 244588 3290
rect 244640 3238 244652 3290
rect 244704 3238 244716 3290
rect 244768 3238 244780 3290
rect 244832 3238 244838 3290
rect 244518 2202 244838 3238
rect 249720 2922 249748 4490
rect 249812 4282 249840 4490
rect 249800 4276 249852 4282
rect 249800 4218 249852 4224
rect 264348 4078 264376 5578
rect 293328 5098 293356 6190
rect 295064 5636 295116 5642
rect 295064 5578 295116 5584
rect 293316 5092 293368 5098
rect 293316 5034 293368 5040
rect 264704 4820 264756 4826
rect 264704 4762 264756 4768
rect 264716 4622 264744 4762
rect 264704 4616 264756 4622
rect 264704 4558 264756 4564
rect 265256 4548 265308 4554
rect 265256 4490 265308 4496
rect 264336 4072 264388 4078
rect 264336 4014 264388 4020
rect 265268 3126 265296 4490
rect 295076 3738 295104 5578
rect 308692 5370 308720 6190
rect 311072 5704 311124 5710
rect 311072 5646 311124 5652
rect 308680 5364 308732 5370
rect 308680 5306 308732 5312
rect 311084 5166 311112 5646
rect 311912 5574 311940 6258
rect 313752 6118 313780 6258
rect 339408 6248 339460 6254
rect 339408 6190 339460 6196
rect 354588 6248 354640 6254
rect 354588 6190 354640 6196
rect 313740 6112 313792 6118
rect 313740 6054 313792 6060
rect 338212 6112 338264 6118
rect 338212 6054 338264 6060
rect 311900 5568 311952 5574
rect 311900 5510 311952 5516
rect 309968 5160 310020 5166
rect 309968 5102 310020 5108
rect 311072 5160 311124 5166
rect 311072 5102 311124 5108
rect 309324 4684 309376 4690
rect 309324 4626 309376 4632
rect 308864 4616 308916 4622
rect 308864 4558 308916 4564
rect 295984 4548 296036 4554
rect 295984 4490 296036 4496
rect 295064 3732 295116 3738
rect 295064 3674 295116 3680
rect 295996 3670 296024 4490
rect 306472 4140 306524 4146
rect 306472 4082 306524 4088
rect 296720 4072 296772 4078
rect 296720 4014 296772 4020
rect 296732 3942 296760 4014
rect 306484 3942 306512 4082
rect 307024 4004 307076 4010
rect 307024 3946 307076 3952
rect 296720 3936 296772 3942
rect 296720 3878 296772 3884
rect 306472 3936 306524 3942
rect 306472 3878 306524 3884
rect 307036 3738 307064 3946
rect 308876 3942 308904 4558
rect 309336 4282 309364 4626
rect 309324 4276 309376 4282
rect 309324 4218 309376 4224
rect 307116 3936 307168 3942
rect 307116 3878 307168 3884
rect 308864 3936 308916 3942
rect 308864 3878 308916 3884
rect 307024 3732 307076 3738
rect 307024 3674 307076 3680
rect 295984 3664 296036 3670
rect 295984 3606 296036 3612
rect 295708 3188 295760 3194
rect 295708 3130 295760 3136
rect 304816 3188 304868 3194
rect 304816 3130 304868 3136
rect 264796 3120 264848 3126
rect 264796 3062 264848 3068
rect 265256 3120 265308 3126
rect 265256 3062 265308 3068
rect 249708 2916 249760 2922
rect 249708 2858 249760 2864
rect 248972 2848 249024 2854
rect 248972 2790 249024 2796
rect 248984 2446 249012 2790
rect 264808 2446 264836 3062
rect 279608 2848 279660 2854
rect 279608 2790 279660 2796
rect 248972 2440 249024 2446
rect 248972 2382 249024 2388
rect 264796 2440 264848 2446
rect 264796 2382 264848 2388
rect 279620 2378 279648 2790
rect 295720 2446 295748 3130
rect 304828 3058 304856 3130
rect 304816 3052 304868 3058
rect 304816 2994 304868 3000
rect 295708 2440 295760 2446
rect 295708 2382 295760 2388
rect 307128 2378 307156 3878
rect 308876 3058 308904 3878
rect 309980 3466 310008 5102
rect 310796 4616 310848 4622
rect 310796 4558 310848 4564
rect 310336 4548 310388 4554
rect 310336 4490 310388 4496
rect 310348 3738 310376 4490
rect 310808 4214 310836 4558
rect 310796 4208 310848 4214
rect 310796 4150 310848 4156
rect 310336 3732 310388 3738
rect 310336 3674 310388 3680
rect 311084 3534 311112 5102
rect 311912 4554 311940 5510
rect 311624 4548 311676 4554
rect 311624 4490 311676 4496
rect 311900 4548 311952 4554
rect 311900 4490 311952 4496
rect 311072 3528 311124 3534
rect 311072 3470 311124 3476
rect 309968 3460 310020 3466
rect 309968 3402 310020 3408
rect 308864 3052 308916 3058
rect 308864 2994 308916 3000
rect 311164 2984 311216 2990
rect 311164 2926 311216 2932
rect 311176 2446 311204 2926
rect 311636 2514 311664 4490
rect 313752 4486 313780 6054
rect 338224 5914 338252 6054
rect 338212 5908 338264 5914
rect 338212 5850 338264 5856
rect 339420 4758 339448 6190
rect 339868 5228 339920 5234
rect 339868 5170 339920 5176
rect 339880 5030 339908 5170
rect 340696 5160 340748 5166
rect 340696 5102 340748 5108
rect 339868 5024 339920 5030
rect 339868 4966 339920 4972
rect 339408 4752 339460 4758
rect 339408 4694 339460 4700
rect 313740 4480 313792 4486
rect 313740 4422 313792 4428
rect 340708 4078 340736 5102
rect 354600 4690 354628 6190
rect 405801 6010 406121 6784
rect 405801 5958 405807 6010
rect 405859 5958 405871 6010
rect 405923 5958 405935 6010
rect 405987 5958 405999 6010
rect 406051 5958 406063 6010
rect 406115 5958 406121 6010
rect 405801 5721 406121 5958
rect 405801 5665 405813 5721
rect 405869 5665 405893 5721
rect 405949 5665 405973 5721
rect 406029 5665 406053 5721
rect 406109 5665 406121 5721
rect 405801 5641 406121 5665
rect 405801 5585 405813 5641
rect 405869 5585 405893 5641
rect 405949 5585 405973 5641
rect 406029 5585 406053 5641
rect 406109 5585 406121 5641
rect 405801 5561 406121 5585
rect 405801 5505 405813 5561
rect 405869 5505 405893 5561
rect 405949 5505 405973 5561
rect 406029 5505 406053 5561
rect 406109 5505 406121 5561
rect 405801 5481 406121 5505
rect 405801 5425 405813 5481
rect 405869 5425 405893 5481
rect 405949 5425 405973 5481
rect 406029 5425 406053 5481
rect 406109 5425 406121 5481
rect 355968 5160 356020 5166
rect 355968 5102 356020 5108
rect 387064 5160 387116 5166
rect 387064 5102 387116 5108
rect 402520 5160 402572 5166
rect 402520 5102 402572 5108
rect 404544 5160 404596 5166
rect 404544 5102 404596 5108
rect 354588 4684 354640 4690
rect 354588 4626 354640 4632
rect 355980 4146 356008 5102
rect 341340 4140 341392 4146
rect 341340 4082 341392 4088
rect 355968 4140 356020 4146
rect 355968 4082 356020 4088
rect 340696 4072 340748 4078
rect 340696 4014 340748 4020
rect 341352 3602 341380 4082
rect 342076 4072 342128 4078
rect 342720 4072 342772 4078
rect 342128 4020 342300 4026
rect 342076 4014 342300 4020
rect 342720 4014 342772 4020
rect 358084 4072 358136 4078
rect 358084 4014 358136 4020
rect 342088 4010 342300 4014
rect 342088 4004 342312 4010
rect 342088 3998 342260 4004
rect 342260 3946 342312 3952
rect 341340 3596 341392 3602
rect 341340 3538 341392 3544
rect 342732 3398 342760 4014
rect 342720 3392 342772 3398
rect 342720 3334 342772 3340
rect 358096 3194 358124 4014
rect 387076 3602 387104 5102
rect 387800 4140 387852 4146
rect 387800 4082 387852 4088
rect 387812 3942 387840 4082
rect 388996 4072 389048 4078
rect 388996 4014 389048 4020
rect 387800 3936 387852 3942
rect 387800 3878 387852 3884
rect 387984 3664 388036 3670
rect 387984 3606 388036 3612
rect 387064 3596 387116 3602
rect 387064 3538 387116 3544
rect 326344 3188 326396 3194
rect 326344 3130 326396 3136
rect 358084 3188 358136 3194
rect 358084 3130 358136 3136
rect 326356 2582 326384 3130
rect 387996 3126 388024 3606
rect 357072 3120 357124 3126
rect 357072 3062 357124 3068
rect 387984 3120 388036 3126
rect 387984 3062 388036 3068
rect 326528 2848 326580 2854
rect 326528 2790 326580 2796
rect 342076 2848 342128 2854
rect 342076 2790 342128 2796
rect 326344 2576 326396 2582
rect 326344 2518 326396 2524
rect 311624 2508 311676 2514
rect 311624 2450 311676 2456
rect 311164 2440 311216 2446
rect 311164 2382 311216 2388
rect 326540 2378 326568 2790
rect 342088 2446 342116 2790
rect 357084 2446 357112 3062
rect 372620 2848 372672 2854
rect 372620 2790 372672 2796
rect 372632 2446 372660 2790
rect 387996 2446 388024 3062
rect 389008 2922 389036 4014
rect 402532 3058 402560 5102
rect 404556 4486 404584 5102
rect 405801 4922 406121 5425
rect 405801 4870 405807 4922
rect 405859 4870 405871 4922
rect 405923 4870 405935 4922
rect 405987 4870 405999 4922
rect 406051 4870 406063 4922
rect 406115 4870 406121 4922
rect 404544 4480 404596 4486
rect 404544 4422 404596 4428
rect 405801 4362 406121 4870
rect 406461 9784 406781 9796
rect 406461 9728 406473 9784
rect 406529 9728 406553 9784
rect 406609 9728 406633 9784
rect 406689 9728 406713 9784
rect 406769 9728 406781 9784
rect 406461 9704 406781 9728
rect 406461 9648 406473 9704
rect 406529 9648 406553 9704
rect 406609 9648 406633 9704
rect 406689 9648 406713 9704
rect 406769 9648 406781 9704
rect 406461 9624 406781 9648
rect 406461 9568 406473 9624
rect 406529 9568 406553 9624
rect 406609 9568 406633 9624
rect 406689 9568 406713 9624
rect 406769 9568 406781 9624
rect 406461 9544 406781 9568
rect 406461 9488 406473 9544
rect 406529 9488 406553 9544
rect 406609 9488 406633 9544
rect 406689 9488 406713 9544
rect 406769 9488 406781 9544
rect 406461 7740 406781 9488
rect 406461 7684 406473 7740
rect 406529 7684 406553 7740
rect 406609 7684 406633 7740
rect 406689 7684 406713 7740
rect 406769 7684 406781 7740
rect 406461 7660 406781 7684
rect 406461 7642 406473 7660
rect 406529 7642 406553 7660
rect 406609 7642 406633 7660
rect 406689 7642 406713 7660
rect 406769 7642 406781 7660
rect 406461 7590 406467 7642
rect 406529 7604 406531 7642
rect 406711 7604 406713 7642
rect 406519 7590 406531 7604
rect 406583 7590 406595 7604
rect 406647 7590 406659 7604
rect 406711 7590 406723 7604
rect 406775 7590 406781 7642
rect 406461 7580 406781 7590
rect 406461 7524 406473 7580
rect 406529 7524 406553 7580
rect 406609 7524 406633 7580
rect 406689 7524 406713 7580
rect 406769 7524 406781 7580
rect 406461 7500 406781 7524
rect 406461 7444 406473 7500
rect 406529 7444 406553 7500
rect 406609 7444 406633 7500
rect 406689 7444 406713 7500
rect 406769 7444 406781 7500
rect 406461 6554 406781 7444
rect 406461 6502 406467 6554
rect 406519 6502 406531 6554
rect 406583 6502 406595 6554
rect 406647 6502 406659 6554
rect 406711 6502 406723 6554
rect 406775 6502 406781 6554
rect 406461 6381 406781 6502
rect 406461 6325 406473 6381
rect 406529 6325 406553 6381
rect 406609 6325 406633 6381
rect 406689 6325 406713 6381
rect 406769 6325 406781 6381
rect 406461 6301 406781 6325
rect 406461 6245 406473 6301
rect 406529 6245 406553 6301
rect 406609 6245 406633 6301
rect 406689 6245 406713 6301
rect 406769 6245 406781 6301
rect 406461 6221 406781 6245
rect 406461 6165 406473 6221
rect 406529 6165 406553 6221
rect 406609 6165 406633 6221
rect 406689 6165 406713 6221
rect 406769 6165 406781 6221
rect 406461 6141 406781 6165
rect 406461 6085 406473 6141
rect 406529 6085 406553 6141
rect 406609 6085 406633 6141
rect 406689 6085 406713 6141
rect 406769 6085 406781 6141
rect 406461 5466 406781 6085
rect 406461 5414 406467 5466
rect 406519 5414 406531 5466
rect 406583 5414 406595 5466
rect 406647 5414 406659 5466
rect 406711 5414 406723 5466
rect 406775 5414 406781 5466
rect 406461 5022 406781 5414
rect 567744 9124 568064 9796
rect 567744 9068 567756 9124
rect 567812 9068 567836 9124
rect 567892 9068 567916 9124
rect 567972 9068 567996 9124
rect 568052 9068 568064 9124
rect 567744 9044 568064 9068
rect 567744 8988 567756 9044
rect 567812 8988 567836 9044
rect 567892 8988 567916 9044
rect 567972 8988 567996 9044
rect 568052 8988 568064 9044
rect 567744 8964 568064 8988
rect 567744 8908 567756 8964
rect 567812 8908 567836 8964
rect 567892 8908 567916 8964
rect 567972 8908 567996 8964
rect 568052 8908 568064 8964
rect 567744 8884 568064 8908
rect 567744 8828 567756 8884
rect 567812 8828 567836 8884
rect 567892 8828 567916 8884
rect 567972 8828 567996 8884
rect 568052 8828 568064 8884
rect 567744 7098 568064 8828
rect 567744 7046 567750 7098
rect 567802 7080 567814 7098
rect 567866 7080 567878 7098
rect 567930 7080 567942 7098
rect 567994 7080 568006 7098
rect 567812 7046 567814 7080
rect 567994 7046 567996 7080
rect 568058 7046 568064 7098
rect 567744 7024 567756 7046
rect 567812 7024 567836 7046
rect 567892 7024 567916 7046
rect 567972 7024 567996 7046
rect 568052 7024 568064 7046
rect 567744 7000 568064 7024
rect 567744 6944 567756 7000
rect 567812 6944 567836 7000
rect 567892 6944 567916 7000
rect 567972 6944 567996 7000
rect 568052 6944 568064 7000
rect 567744 6920 568064 6944
rect 567744 6864 567756 6920
rect 567812 6864 567836 6920
rect 567892 6864 567916 6920
rect 567972 6864 567996 6920
rect 568052 6864 568064 6920
rect 567744 6840 568064 6864
rect 567744 6784 567756 6840
rect 567812 6784 567836 6840
rect 567892 6784 567916 6840
rect 567972 6784 567996 6840
rect 568052 6784 568064 6840
rect 567744 6010 568064 6784
rect 567744 5958 567750 6010
rect 567802 5958 567814 6010
rect 567866 5958 567878 6010
rect 567930 5958 567942 6010
rect 567994 5958 568006 6010
rect 568058 5958 568064 6010
rect 567744 5721 568064 5958
rect 567744 5665 567756 5721
rect 567812 5665 567836 5721
rect 567892 5665 567916 5721
rect 567972 5665 567996 5721
rect 568052 5665 568064 5721
rect 567744 5641 568064 5665
rect 567744 5585 567756 5641
rect 567812 5585 567836 5641
rect 567892 5585 567916 5641
rect 567972 5585 567996 5641
rect 568052 5585 568064 5641
rect 567744 5561 568064 5585
rect 567744 5505 567756 5561
rect 567812 5505 567836 5561
rect 567892 5505 567916 5561
rect 567972 5505 567996 5561
rect 568052 5505 568064 5561
rect 567744 5481 568064 5505
rect 567744 5425 567756 5481
rect 567812 5425 567836 5481
rect 567892 5425 567916 5481
rect 567972 5425 567996 5481
rect 568052 5425 568064 5481
rect 432144 5228 432196 5234
rect 432144 5170 432196 5176
rect 406461 4966 406473 5022
rect 406529 4966 406553 5022
rect 406609 4966 406633 5022
rect 406689 4966 406713 5022
rect 406769 4966 406781 5022
rect 407304 5024 407356 5030
rect 407304 4966 407356 4972
rect 406461 4942 406781 4966
rect 406461 4886 406473 4942
rect 406529 4886 406553 4942
rect 406609 4886 406633 4942
rect 406689 4886 406713 4942
rect 406769 4886 406781 4942
rect 406461 4862 406781 4886
rect 406461 4806 406473 4862
rect 406529 4806 406553 4862
rect 406609 4806 406633 4862
rect 406689 4806 406713 4862
rect 406769 4806 406781 4862
rect 407316 4826 407344 4966
rect 406461 4782 406781 4806
rect 406461 4726 406473 4782
rect 406529 4726 406553 4782
rect 406609 4726 406633 4782
rect 406689 4726 406713 4782
rect 406769 4726 406781 4782
rect 407304 4820 407356 4826
rect 407304 4762 407356 4768
rect 432156 4758 432184 5170
rect 433248 5160 433300 5166
rect 433248 5102 433300 5108
rect 448796 5160 448848 5166
rect 448796 5102 448848 5108
rect 406200 4480 406252 4486
rect 406200 4422 406252 4428
rect 405801 4306 405813 4362
rect 405869 4306 405893 4362
rect 405949 4306 405973 4362
rect 406029 4306 406053 4362
rect 406109 4306 406121 4362
rect 405801 4282 406121 4306
rect 405801 4226 405813 4282
rect 405869 4226 405893 4282
rect 405949 4226 405973 4282
rect 406029 4226 406053 4282
rect 406109 4226 406121 4282
rect 405801 4202 406121 4226
rect 405801 4146 405813 4202
rect 405869 4146 405893 4202
rect 405949 4146 405973 4202
rect 406029 4146 406053 4202
rect 406109 4146 406121 4202
rect 402612 4140 402664 4146
rect 402612 4082 402664 4088
rect 405801 4122 406121 4146
rect 402624 3942 402652 4082
rect 404452 4072 404504 4078
rect 404452 4014 404504 4020
rect 405801 4066 405813 4122
rect 405869 4066 405893 4122
rect 405949 4066 405973 4122
rect 406029 4066 406053 4122
rect 406109 4066 406121 4122
rect 402612 3936 402664 3942
rect 402612 3878 402664 3884
rect 402624 3738 402652 3878
rect 404464 3738 404492 4014
rect 405801 3834 406121 4066
rect 405801 3782 405807 3834
rect 405859 3782 405871 3834
rect 405923 3782 405935 3834
rect 405987 3782 405999 3834
rect 406051 3782 406063 3834
rect 406115 3782 406121 3834
rect 402612 3732 402664 3738
rect 402612 3674 402664 3680
rect 404452 3732 404504 3738
rect 404452 3674 404504 3680
rect 403348 3528 403400 3534
rect 403348 3470 403400 3476
rect 402520 3052 402572 3058
rect 402520 2994 402572 3000
rect 403360 2990 403388 3470
rect 405801 3003 406121 3782
rect 406212 3466 406240 4422
rect 406461 4378 406781 4726
rect 432144 4752 432196 4758
rect 432144 4694 432196 4700
rect 406461 4326 406467 4378
rect 406519 4326 406531 4378
rect 406583 4326 406595 4378
rect 406647 4326 406659 4378
rect 406711 4326 406723 4378
rect 406775 4326 406781 4378
rect 406461 3663 406781 4326
rect 433260 3942 433288 5102
rect 447416 5024 447468 5030
rect 447416 4966 447468 4972
rect 447428 4690 447456 4966
rect 447416 4684 447468 4690
rect 447416 4626 447468 4632
rect 435364 4072 435416 4078
rect 435364 4014 435416 4020
rect 433248 3936 433300 3942
rect 433248 3878 433300 3884
rect 406461 3607 406473 3663
rect 406529 3607 406553 3663
rect 406609 3607 406633 3663
rect 406689 3607 406713 3663
rect 406769 3607 406781 3663
rect 406461 3583 406781 3607
rect 406461 3527 406473 3583
rect 406529 3527 406553 3583
rect 406609 3527 406633 3583
rect 406689 3527 406713 3583
rect 406769 3527 406781 3583
rect 406461 3503 406781 3527
rect 406200 3460 406252 3466
rect 406200 3402 406252 3408
rect 406461 3447 406473 3503
rect 406529 3447 406553 3503
rect 406609 3447 406633 3503
rect 406689 3447 406713 3503
rect 406769 3447 406781 3503
rect 406461 3423 406781 3447
rect 403348 2984 403400 2990
rect 403348 2926 403400 2932
rect 405801 2947 405813 3003
rect 405869 2947 405893 3003
rect 405949 2947 405973 3003
rect 406029 2947 406053 3003
rect 406109 2947 406121 3003
rect 388996 2916 389048 2922
rect 388996 2858 389048 2864
rect 342076 2440 342128 2446
rect 342076 2382 342128 2388
rect 357072 2440 357124 2446
rect 357072 2382 357124 2388
rect 372620 2440 372672 2446
rect 372620 2382 372672 2388
rect 387984 2440 388036 2446
rect 387984 2382 388036 2388
rect 279608 2372 279660 2378
rect 279608 2314 279660 2320
rect 307116 2372 307168 2378
rect 307116 2314 307168 2320
rect 326528 2372 326580 2378
rect 326528 2314 326580 2320
rect 249156 2304 249208 2310
rect 249156 2246 249208 2252
rect 264612 2304 264664 2310
rect 264612 2246 264664 2252
rect 244518 2150 244524 2202
rect 244576 2150 244588 2202
rect 244640 2150 244652 2202
rect 244704 2150 244716 2202
rect 244768 2150 244780 2202
rect 244832 2150 244838 2202
rect 244518 304 244838 2150
rect 249168 814 249196 2246
rect 264624 814 264652 2246
rect 279620 814 279648 2314
rect 293960 2304 294012 2310
rect 293960 2246 294012 2252
rect 309140 2304 309192 2310
rect 309140 2246 309192 2252
rect 293972 814 294000 2246
rect 249156 808 249208 814
rect 249156 750 249208 756
rect 264612 808 264664 814
rect 264612 750 264664 756
rect 279608 808 279660 814
rect 279608 750 279660 756
rect 293960 808 294012 814
rect 293960 750 294012 756
rect 244518 248 244530 304
rect 244586 248 244610 304
rect 244666 248 244690 304
rect 244746 248 244770 304
rect 244826 248 244838 304
rect 244518 224 244838 248
rect 244518 168 244530 224
rect 244586 168 244610 224
rect 244666 168 244690 224
rect 244746 168 244770 224
rect 244826 168 244838 224
rect 244518 144 244838 168
rect 244518 88 244530 144
rect 244586 88 244610 144
rect 244666 88 244690 144
rect 244746 88 244770 144
rect 244826 88 244838 144
rect 244518 64 244838 88
rect 309152 66 309180 2246
rect 326540 814 326568 2314
rect 339500 2304 339552 2310
rect 339500 2246 339552 2252
rect 357348 2304 357400 2310
rect 357348 2246 357400 2252
rect 339512 814 339540 2246
rect 357360 814 357388 2246
rect 372632 814 372660 2382
rect 403360 2378 403388 2926
rect 405801 2923 406121 2947
rect 405801 2867 405813 2923
rect 405869 2867 405893 2923
rect 405949 2867 405973 2923
rect 406029 2867 406053 2923
rect 406109 2867 406121 2923
rect 405801 2843 406121 2867
rect 405801 2787 405813 2843
rect 405869 2787 405893 2843
rect 405949 2787 405973 2843
rect 406029 2787 406053 2843
rect 406109 2787 406121 2843
rect 405801 2763 406121 2787
rect 405801 2746 405813 2763
rect 405869 2746 405893 2763
rect 405949 2746 405973 2763
rect 406029 2746 406053 2763
rect 406109 2746 406121 2763
rect 405801 2694 405807 2746
rect 405869 2707 405871 2746
rect 406051 2707 406053 2746
rect 405859 2694 405871 2707
rect 405923 2694 405935 2707
rect 405987 2694 405999 2707
rect 406051 2694 406063 2707
rect 406115 2694 406121 2746
rect 403348 2372 403400 2378
rect 403348 2314 403400 2320
rect 386420 2304 386472 2310
rect 386420 2246 386472 2252
rect 402704 2304 402756 2310
rect 402704 2246 402756 2252
rect 326528 808 326580 814
rect 326528 750 326580 756
rect 339500 808 339552 814
rect 339500 750 339552 756
rect 357348 808 357400 814
rect 357348 750 357400 756
rect 372620 808 372672 814
rect 372620 750 372672 756
rect 386432 66 386460 2246
rect 402716 814 402744 2246
rect 405801 964 406121 2694
rect 405801 908 405813 964
rect 405869 908 405893 964
rect 405949 908 405973 964
rect 406029 908 406053 964
rect 406109 908 406121 964
rect 405801 884 406121 908
rect 405801 828 405813 884
rect 405869 828 405893 884
rect 405949 828 405973 884
rect 406029 828 406053 884
rect 406109 828 406121 884
rect 402704 808 402756 814
rect 402704 750 402756 756
rect 405801 804 406121 828
rect 405801 748 405813 804
rect 405869 748 405893 804
rect 405949 748 405973 804
rect 406029 748 406053 804
rect 406109 748 406121 804
rect 405801 724 406121 748
rect 405801 668 405813 724
rect 405869 668 405893 724
rect 405949 668 405973 724
rect 406029 668 406053 724
rect 406109 668 406121 724
rect 244518 8 244530 64
rect 244586 8 244610 64
rect 244666 8 244690 64
rect 244746 8 244770 64
rect 244826 8 244838 64
rect 244518 -4 244838 8
rect 309140 60 309192 66
rect 309140 2 309192 8
rect 386420 60 386472 66
rect 386420 2 386472 8
rect 405801 -4 406121 668
rect 406461 3367 406473 3423
rect 406529 3367 406553 3423
rect 406609 3367 406633 3423
rect 406689 3367 406713 3423
rect 406769 3367 406781 3423
rect 406461 3290 406781 3367
rect 434352 3392 434404 3398
rect 434352 3334 434404 3340
rect 406461 3238 406467 3290
rect 406519 3238 406531 3290
rect 406583 3238 406595 3290
rect 406647 3238 406659 3290
rect 406711 3238 406723 3290
rect 406775 3238 406781 3290
rect 406461 2202 406781 3238
rect 434364 3126 434392 3334
rect 435376 3126 435404 4014
rect 448808 3398 448836 5102
rect 567744 4922 568064 5425
rect 567744 4870 567750 4922
rect 567802 4870 567814 4922
rect 567866 4870 567878 4922
rect 567930 4870 567942 4922
rect 567994 4870 568006 4922
rect 568058 4870 568064 4922
rect 499948 4820 500000 4826
rect 499948 4762 500000 4768
rect 499960 4214 499988 4762
rect 567744 4362 568064 4870
rect 567744 4306 567756 4362
rect 567812 4306 567836 4362
rect 567892 4306 567916 4362
rect 567972 4306 567996 4362
rect 568052 4306 568064 4362
rect 567744 4282 568064 4306
rect 567744 4226 567756 4282
rect 567812 4226 567836 4282
rect 567892 4226 567916 4282
rect 567972 4226 567996 4282
rect 568052 4226 568064 4282
rect 499948 4208 500000 4214
rect 499948 4150 500000 4156
rect 567744 4202 568064 4226
rect 567744 4146 567756 4202
rect 567812 4146 567836 4202
rect 567892 4146 567916 4202
rect 567972 4146 567996 4202
rect 568052 4146 568064 4202
rect 479892 4140 479944 4146
rect 479892 4082 479944 4088
rect 495440 4140 495492 4146
rect 495440 4082 495492 4088
rect 500500 4140 500552 4146
rect 500500 4082 500552 4088
rect 567744 4122 568064 4146
rect 450820 4072 450872 4078
rect 450820 4014 450872 4020
rect 448796 3392 448848 3398
rect 448796 3334 448848 3340
rect 450832 3194 450860 4014
rect 479904 3942 479932 4082
rect 495452 3942 495480 4082
rect 497188 4072 497240 4078
rect 497188 4014 497240 4020
rect 479892 3936 479944 3942
rect 479892 3878 479944 3884
rect 495440 3936 495492 3942
rect 495440 3878 495492 3884
rect 479904 3602 479932 3878
rect 479892 3596 479944 3602
rect 479892 3538 479944 3544
rect 450268 3188 450320 3194
rect 450268 3130 450320 3136
rect 450820 3188 450872 3194
rect 450820 3130 450872 3136
rect 434352 3120 434404 3126
rect 434352 3062 434404 3068
rect 435364 3120 435416 3126
rect 435364 3062 435416 3068
rect 415308 2848 415360 2854
rect 415308 2790 415360 2796
rect 415320 2650 415348 2790
rect 415308 2644 415360 2650
rect 415308 2586 415360 2592
rect 434364 2446 434392 3062
rect 450280 2446 450308 3130
rect 495452 3058 495480 3878
rect 497200 3738 497228 4014
rect 500512 3942 500540 4082
rect 567744 4066 567756 4122
rect 567812 4066 567836 4122
rect 567892 4066 567916 4122
rect 567972 4066 567996 4122
rect 568052 4066 568064 4122
rect 500500 3936 500552 3942
rect 500500 3878 500552 3884
rect 567744 3834 568064 4066
rect 567744 3782 567750 3834
rect 567802 3782 567814 3834
rect 567866 3782 567878 3834
rect 567930 3782 567942 3834
rect 567994 3782 568006 3834
rect 568058 3782 568064 3834
rect 496176 3732 496228 3738
rect 496176 3674 496228 3680
rect 497188 3732 497240 3738
rect 497188 3674 497240 3680
rect 496188 3058 496216 3674
rect 497280 3528 497332 3534
rect 497280 3470 497332 3476
rect 499856 3528 499908 3534
rect 499856 3470 499908 3476
rect 497292 3058 497320 3470
rect 499868 3398 499896 3470
rect 499856 3392 499908 3398
rect 499856 3334 499908 3340
rect 495440 3052 495492 3058
rect 495440 2994 495492 3000
rect 496176 3052 496228 3058
rect 496176 2994 496228 3000
rect 497280 3052 497332 3058
rect 497280 2994 497332 3000
rect 465264 2848 465316 2854
rect 465264 2790 465316 2796
rect 480812 2848 480864 2854
rect 480812 2790 480864 2796
rect 465276 2446 465304 2790
rect 480824 2446 480852 2790
rect 496188 2446 496216 2994
rect 418068 2440 418120 2446
rect 418068 2382 418120 2388
rect 434352 2440 434404 2446
rect 434352 2382 434404 2388
rect 450268 2440 450320 2446
rect 450268 2382 450320 2388
rect 465264 2440 465316 2446
rect 465264 2382 465316 2388
rect 480812 2440 480864 2446
rect 480812 2382 480864 2388
rect 496176 2440 496228 2446
rect 496176 2382 496228 2388
rect 406461 2150 406467 2202
rect 406519 2150 406531 2202
rect 406583 2150 406595 2202
rect 406647 2150 406659 2202
rect 406711 2150 406723 2202
rect 406775 2150 406781 2202
rect 406461 304 406781 2150
rect 418080 814 418108 2382
rect 432788 2304 432840 2310
rect 432788 2246 432840 2252
rect 450084 2304 450136 2310
rect 450084 2246 450136 2252
rect 432800 814 432828 2246
rect 450096 814 450124 2246
rect 418068 808 418120 814
rect 418068 750 418120 756
rect 432788 808 432840 814
rect 432788 750 432840 756
rect 450084 808 450136 814
rect 450084 750 450136 756
rect 406461 248 406473 304
rect 406529 248 406553 304
rect 406609 248 406633 304
rect 406689 248 406713 304
rect 406769 248 406781 304
rect 406461 224 406781 248
rect 406461 168 406473 224
rect 406529 168 406553 224
rect 406609 168 406633 224
rect 406689 168 406713 224
rect 406769 168 406781 224
rect 406461 144 406781 168
rect 406461 88 406473 144
rect 406529 88 406553 144
rect 406609 88 406633 144
rect 406689 88 406713 144
rect 406769 88 406781 144
rect 406461 64 406781 88
rect 465276 66 465304 2382
rect 499868 2378 499896 3334
rect 543004 3188 543056 3194
rect 543004 3130 543056 3136
rect 527548 3120 527600 3126
rect 527548 3062 527600 3068
rect 510528 3052 510580 3058
rect 510528 2994 510580 3000
rect 510540 2650 510568 2994
rect 510528 2644 510580 2650
rect 510528 2586 510580 2592
rect 527560 2446 527588 3062
rect 543016 2446 543044 3130
rect 567744 3003 568064 3782
rect 567744 2947 567756 3003
rect 567812 2947 567836 3003
rect 567892 2947 567916 3003
rect 567972 2947 567996 3003
rect 568052 2947 568064 3003
rect 567744 2923 568064 2947
rect 567744 2867 567756 2923
rect 567812 2867 567836 2923
rect 567892 2867 567916 2923
rect 567972 2867 567996 2923
rect 568052 2867 568064 2923
rect 558000 2848 558052 2854
rect 558000 2790 558052 2796
rect 567744 2843 568064 2867
rect 558012 2446 558040 2790
rect 567744 2787 567756 2843
rect 567812 2787 567836 2843
rect 567892 2787 567916 2843
rect 567972 2787 567996 2843
rect 568052 2787 568064 2843
rect 567744 2763 568064 2787
rect 567744 2746 567756 2763
rect 567812 2746 567836 2763
rect 567892 2746 567916 2763
rect 567972 2746 567996 2763
rect 568052 2746 568064 2763
rect 567744 2694 567750 2746
rect 567812 2707 567814 2746
rect 567994 2707 567996 2746
rect 567802 2694 567814 2707
rect 567866 2694 567878 2707
rect 567930 2694 567942 2707
rect 567994 2694 568006 2707
rect 568058 2694 568064 2746
rect 511908 2440 511960 2446
rect 511908 2382 511960 2388
rect 527548 2440 527600 2446
rect 527548 2382 527600 2388
rect 543004 2440 543056 2446
rect 543004 2382 543056 2388
rect 558000 2440 558052 2446
rect 558000 2382 558052 2388
rect 499856 2372 499908 2378
rect 499856 2314 499908 2320
rect 480996 2304 481048 2310
rect 480996 2246 481048 2252
rect 496452 2304 496504 2310
rect 496452 2246 496504 2252
rect 481008 814 481036 2246
rect 480996 808 481048 814
rect 480996 750 481048 756
rect 496464 66 496492 2246
rect 511920 814 511948 2382
rect 527364 2304 527416 2310
rect 527364 2246 527416 2252
rect 542820 2304 542872 2310
rect 542820 2246 542872 2252
rect 527376 814 527404 2246
rect 511908 808 511960 814
rect 511908 750 511960 756
rect 527364 808 527416 814
rect 527364 750 527416 756
rect 542832 66 542860 2246
rect 558012 814 558040 2382
rect 567744 964 568064 2694
rect 567744 908 567756 964
rect 567812 908 567836 964
rect 567892 908 567916 964
rect 567972 908 567996 964
rect 568052 908 568064 964
rect 567744 884 568064 908
rect 567744 828 567756 884
rect 567812 828 567836 884
rect 567892 828 567916 884
rect 567972 828 567996 884
rect 568052 828 568064 884
rect 558000 808 558052 814
rect 558000 750 558052 756
rect 567744 804 568064 828
rect 567744 748 567756 804
rect 567812 748 567836 804
rect 567892 748 567916 804
rect 567972 748 567996 804
rect 568052 748 568064 804
rect 567744 724 568064 748
rect 567744 668 567756 724
rect 567812 668 567836 724
rect 567892 668 567916 724
rect 567972 668 567996 724
rect 568052 668 568064 724
rect 406461 8 406473 64
rect 406529 8 406553 64
rect 406609 8 406633 64
rect 406689 8 406713 64
rect 406769 8 406781 64
rect 406461 -4 406781 8
rect 465264 60 465316 66
rect 465264 2 465316 8
rect 496452 60 496504 66
rect 496452 2 496504 8
rect 542820 60 542872 66
rect 542820 2 542872 8
rect 567744 -4 568064 668
rect 568404 9784 568724 9796
rect 568404 9728 568416 9784
rect 568472 9728 568496 9784
rect 568552 9728 568576 9784
rect 568632 9728 568656 9784
rect 568712 9728 568724 9784
rect 568404 9704 568724 9728
rect 568404 9648 568416 9704
rect 568472 9648 568496 9704
rect 568552 9648 568576 9704
rect 568632 9648 568656 9704
rect 568712 9648 568724 9704
rect 568404 9624 568724 9648
rect 568404 9568 568416 9624
rect 568472 9568 568496 9624
rect 568552 9568 568576 9624
rect 568632 9568 568656 9624
rect 568712 9568 568724 9624
rect 568404 9544 568724 9568
rect 568404 9488 568416 9544
rect 568472 9488 568496 9544
rect 568552 9488 568576 9544
rect 568632 9488 568656 9544
rect 568712 9488 568724 9544
rect 568404 7740 568724 9488
rect 650736 9784 651056 9796
rect 650736 9728 650748 9784
rect 650804 9728 650828 9784
rect 650884 9728 650908 9784
rect 650964 9728 650988 9784
rect 651044 9728 651056 9784
rect 650736 9704 651056 9728
rect 650736 9648 650748 9704
rect 650804 9648 650828 9704
rect 650884 9648 650908 9704
rect 650964 9648 650988 9704
rect 651044 9648 651056 9704
rect 650736 9624 651056 9648
rect 650736 9568 650748 9624
rect 650804 9568 650828 9624
rect 650884 9568 650908 9624
rect 650964 9568 650988 9624
rect 651044 9568 651056 9624
rect 650736 9544 651056 9568
rect 650736 9488 650748 9544
rect 650804 9488 650828 9544
rect 650884 9488 650908 9544
rect 650964 9488 650988 9544
rect 651044 9488 651056 9544
rect 568404 7684 568416 7740
rect 568472 7684 568496 7740
rect 568552 7684 568576 7740
rect 568632 7684 568656 7740
rect 568712 7684 568724 7740
rect 568404 7660 568724 7684
rect 568404 7642 568416 7660
rect 568472 7642 568496 7660
rect 568552 7642 568576 7660
rect 568632 7642 568656 7660
rect 568712 7642 568724 7660
rect 568404 7590 568410 7642
rect 568472 7604 568474 7642
rect 568654 7604 568656 7642
rect 568462 7590 568474 7604
rect 568526 7590 568538 7604
rect 568590 7590 568602 7604
rect 568654 7590 568666 7604
rect 568718 7590 568724 7642
rect 568404 7580 568724 7590
rect 568404 7524 568416 7580
rect 568472 7524 568496 7580
rect 568552 7524 568576 7580
rect 568632 7524 568656 7580
rect 568712 7524 568724 7580
rect 568404 7500 568724 7524
rect 568404 7444 568416 7500
rect 568472 7444 568496 7500
rect 568552 7444 568576 7500
rect 568632 7444 568656 7500
rect 568712 7444 568724 7500
rect 568404 6554 568724 7444
rect 568404 6502 568410 6554
rect 568462 6502 568474 6554
rect 568526 6502 568538 6554
rect 568590 6502 568602 6554
rect 568654 6502 568666 6554
rect 568718 6502 568724 6554
rect 568404 6381 568724 6502
rect 568404 6325 568416 6381
rect 568472 6325 568496 6381
rect 568552 6325 568576 6381
rect 568632 6325 568656 6381
rect 568712 6325 568724 6381
rect 568404 6301 568724 6325
rect 568404 6245 568416 6301
rect 568472 6245 568496 6301
rect 568552 6245 568576 6301
rect 568632 6245 568656 6301
rect 568712 6245 568724 6301
rect 568404 6221 568724 6245
rect 568404 6165 568416 6221
rect 568472 6165 568496 6221
rect 568552 6165 568576 6221
rect 568632 6165 568656 6221
rect 568712 6165 568724 6221
rect 568404 6141 568724 6165
rect 568404 6085 568416 6141
rect 568472 6085 568496 6141
rect 568552 6085 568576 6141
rect 568632 6085 568656 6141
rect 568712 6085 568724 6141
rect 568404 5466 568724 6085
rect 568404 5414 568410 5466
rect 568462 5414 568474 5466
rect 568526 5414 568538 5466
rect 568590 5414 568602 5466
rect 568654 5414 568666 5466
rect 568718 5414 568724 5466
rect 568404 5022 568724 5414
rect 568404 4966 568416 5022
rect 568472 4966 568496 5022
rect 568552 4966 568576 5022
rect 568632 4966 568656 5022
rect 568712 4966 568724 5022
rect 568404 4942 568724 4966
rect 568404 4886 568416 4942
rect 568472 4886 568496 4942
rect 568552 4886 568576 4942
rect 568632 4886 568656 4942
rect 568712 4886 568724 4942
rect 568404 4862 568724 4886
rect 568404 4806 568416 4862
rect 568472 4806 568496 4862
rect 568552 4806 568576 4862
rect 568632 4806 568656 4862
rect 568712 4806 568724 4862
rect 568404 4782 568724 4806
rect 568404 4726 568416 4782
rect 568472 4726 568496 4782
rect 568552 4726 568576 4782
rect 568632 4726 568656 4782
rect 568712 4726 568724 4782
rect 568404 4378 568724 4726
rect 568404 4326 568410 4378
rect 568462 4326 568474 4378
rect 568526 4326 568538 4378
rect 568590 4326 568602 4378
rect 568654 4326 568666 4378
rect 568718 4326 568724 4378
rect 568404 3663 568724 4326
rect 650076 9124 650396 9136
rect 650076 9068 650088 9124
rect 650144 9068 650168 9124
rect 650224 9068 650248 9124
rect 650304 9068 650328 9124
rect 650384 9068 650396 9124
rect 650076 9044 650396 9068
rect 650076 8988 650088 9044
rect 650144 8988 650168 9044
rect 650224 8988 650248 9044
rect 650304 8988 650328 9044
rect 650384 8988 650396 9044
rect 650076 8964 650396 8988
rect 650076 8908 650088 8964
rect 650144 8908 650168 8964
rect 650224 8908 650248 8964
rect 650304 8908 650328 8964
rect 650384 8908 650396 8964
rect 650076 8884 650396 8908
rect 650076 8828 650088 8884
rect 650144 8828 650168 8884
rect 650224 8828 650248 8884
rect 650304 8828 650328 8884
rect 650384 8828 650396 8884
rect 650076 7080 650396 8828
rect 650076 7024 650088 7080
rect 650144 7024 650168 7080
rect 650224 7024 650248 7080
rect 650304 7024 650328 7080
rect 650384 7024 650396 7080
rect 650076 7000 650396 7024
rect 650076 6944 650088 7000
rect 650144 6944 650168 7000
rect 650224 6944 650248 7000
rect 650304 6944 650328 7000
rect 650384 6944 650396 7000
rect 650076 6920 650396 6944
rect 650076 6864 650088 6920
rect 650144 6864 650168 6920
rect 650224 6864 650248 6920
rect 650304 6864 650328 6920
rect 650384 6864 650396 6920
rect 650076 6840 650396 6864
rect 650076 6784 650088 6840
rect 650144 6784 650168 6840
rect 650224 6784 650248 6840
rect 650304 6784 650328 6840
rect 650384 6784 650396 6840
rect 650076 5721 650396 6784
rect 650076 5665 650088 5721
rect 650144 5665 650168 5721
rect 650224 5665 650248 5721
rect 650304 5665 650328 5721
rect 650384 5665 650396 5721
rect 650076 5641 650396 5665
rect 650076 5585 650088 5641
rect 650144 5585 650168 5641
rect 650224 5585 650248 5641
rect 650304 5585 650328 5641
rect 650384 5585 650396 5641
rect 650076 5561 650396 5585
rect 650076 5505 650088 5561
rect 650144 5505 650168 5561
rect 650224 5505 650248 5561
rect 650304 5505 650328 5561
rect 650384 5505 650396 5561
rect 650076 5481 650396 5505
rect 650076 5425 650088 5481
rect 650144 5425 650168 5481
rect 650224 5425 650248 5481
rect 650304 5425 650328 5481
rect 650384 5425 650396 5481
rect 650076 4362 650396 5425
rect 650076 4306 650088 4362
rect 650144 4306 650168 4362
rect 650224 4306 650248 4362
rect 650304 4306 650328 4362
rect 650384 4306 650396 4362
rect 650076 4282 650396 4306
rect 650076 4226 650088 4282
rect 650144 4226 650168 4282
rect 650224 4226 650248 4282
rect 650304 4226 650328 4282
rect 650384 4226 650396 4282
rect 650076 4202 650396 4226
rect 650076 4146 650088 4202
rect 650144 4146 650168 4202
rect 650224 4146 650248 4202
rect 650304 4146 650328 4202
rect 650384 4146 650396 4202
rect 650076 4122 650396 4146
rect 619824 4072 619876 4078
rect 619824 4014 619876 4020
rect 650076 4066 650088 4122
rect 650144 4066 650168 4122
rect 650224 4066 650248 4122
rect 650304 4066 650328 4122
rect 650384 4066 650396 4122
rect 573456 4004 573508 4010
rect 573456 3946 573508 3952
rect 568404 3607 568416 3663
rect 568472 3607 568496 3663
rect 568552 3607 568576 3663
rect 568632 3607 568656 3663
rect 568712 3607 568724 3663
rect 568404 3583 568724 3607
rect 568404 3527 568416 3583
rect 568472 3527 568496 3583
rect 568552 3527 568576 3583
rect 568632 3527 568656 3583
rect 568712 3527 568724 3583
rect 568404 3503 568724 3527
rect 568404 3447 568416 3503
rect 568472 3447 568496 3503
rect 568552 3447 568576 3503
rect 568632 3447 568656 3503
rect 568712 3447 568724 3503
rect 568404 3423 568724 3447
rect 568404 3367 568416 3423
rect 568472 3367 568496 3423
rect 568552 3367 568576 3423
rect 568632 3367 568656 3423
rect 568712 3367 568724 3423
rect 568404 3290 568724 3367
rect 568404 3238 568410 3290
rect 568462 3238 568474 3290
rect 568526 3238 568538 3290
rect 568590 3238 568602 3290
rect 568654 3238 568666 3290
rect 568718 3238 568724 3290
rect 568404 2202 568724 3238
rect 573468 3194 573496 3946
rect 594064 3936 594116 3942
rect 594064 3878 594116 3884
rect 588912 3732 588964 3738
rect 588912 3674 588964 3680
rect 588924 3194 588952 3674
rect 573456 3188 573508 3194
rect 573456 3130 573508 3136
rect 588912 3188 588964 3194
rect 588912 3130 588964 3136
rect 573468 2446 573496 3130
rect 588924 2446 588952 3130
rect 594076 3126 594104 3878
rect 619836 3194 619864 4014
rect 635280 3460 635332 3466
rect 635280 3402 635332 3408
rect 635292 3194 635320 3402
rect 619824 3188 619876 3194
rect 619824 3130 619876 3136
rect 635280 3188 635332 3194
rect 635280 3130 635332 3136
rect 594064 3120 594116 3126
rect 594064 3062 594116 3068
rect 602896 3052 602948 3058
rect 602896 2994 602948 3000
rect 602908 2650 602936 2994
rect 602896 2644 602948 2650
rect 602896 2586 602948 2592
rect 619836 2446 619864 3130
rect 635292 2446 635320 3130
rect 650076 3003 650396 4066
rect 650076 2947 650088 3003
rect 650144 2947 650168 3003
rect 650224 2947 650248 3003
rect 650304 2947 650328 3003
rect 650384 2947 650396 3003
rect 650076 2923 650396 2947
rect 650076 2867 650088 2923
rect 650144 2867 650168 2923
rect 650224 2867 650248 2923
rect 650304 2867 650328 2923
rect 650384 2867 650396 2923
rect 650076 2843 650396 2867
rect 650076 2787 650088 2843
rect 650144 2787 650168 2843
rect 650224 2787 650248 2843
rect 650304 2787 650328 2843
rect 650384 2787 650396 2843
rect 650076 2763 650396 2787
rect 650076 2707 650088 2763
rect 650144 2707 650168 2763
rect 650224 2707 650248 2763
rect 650304 2707 650328 2763
rect 650384 2707 650396 2763
rect 573456 2440 573508 2446
rect 573456 2382 573508 2388
rect 588912 2440 588964 2446
rect 588912 2382 588964 2388
rect 604368 2440 604420 2446
rect 604368 2382 604420 2388
rect 619824 2440 619876 2446
rect 619824 2382 619876 2388
rect 635280 2440 635332 2446
rect 635280 2382 635332 2388
rect 573732 2304 573784 2310
rect 573732 2246 573784 2252
rect 589188 2304 589240 2310
rect 589188 2246 589240 2252
rect 568404 2150 568410 2202
rect 568462 2150 568474 2202
rect 568526 2150 568538 2202
rect 568590 2150 568602 2202
rect 568654 2150 568666 2202
rect 568718 2150 568724 2202
rect 568404 304 568724 2150
rect 568404 248 568416 304
rect 568472 248 568496 304
rect 568552 248 568576 304
rect 568632 248 568656 304
rect 568712 248 568724 304
rect 568404 224 568724 248
rect 568404 168 568416 224
rect 568472 168 568496 224
rect 568552 168 568576 224
rect 568632 168 568656 224
rect 568712 168 568724 224
rect 568404 144 568724 168
rect 568404 88 568416 144
rect 568472 88 568496 144
rect 568552 88 568576 144
rect 568632 88 568656 144
rect 568712 88 568724 144
rect 568404 64 568724 88
rect 573744 66 573772 2246
rect 589200 814 589228 2246
rect 604380 814 604408 2382
rect 618260 2304 618312 2310
rect 618260 2246 618312 2252
rect 633440 2304 633492 2310
rect 633440 2246 633492 2252
rect 589188 808 589240 814
rect 589188 750 589240 756
rect 604368 808 604420 814
rect 604368 750 604420 756
rect 618272 66 618300 2246
rect 633452 814 633480 2246
rect 650076 964 650396 2707
rect 650076 908 650088 964
rect 650144 908 650168 964
rect 650224 908 650248 964
rect 650304 908 650328 964
rect 650384 908 650396 964
rect 650076 884 650396 908
rect 650076 828 650088 884
rect 650144 828 650168 884
rect 650224 828 650248 884
rect 650304 828 650328 884
rect 650384 828 650396 884
rect 633440 808 633492 814
rect 633440 750 633492 756
rect 650076 804 650396 828
rect 650076 748 650088 804
rect 650144 748 650168 804
rect 650224 748 650248 804
rect 650304 748 650328 804
rect 650384 748 650396 804
rect 650076 724 650396 748
rect 650076 668 650088 724
rect 650144 668 650168 724
rect 650224 668 650248 724
rect 650304 668 650328 724
rect 650384 668 650396 724
rect 650076 656 650396 668
rect 650736 7740 651056 9488
rect 650736 7684 650748 7740
rect 650804 7684 650828 7740
rect 650884 7684 650908 7740
rect 650964 7684 650988 7740
rect 651044 7684 651056 7740
rect 650736 7660 651056 7684
rect 650736 7604 650748 7660
rect 650804 7604 650828 7660
rect 650884 7604 650908 7660
rect 650964 7604 650988 7660
rect 651044 7604 651056 7660
rect 650736 7580 651056 7604
rect 650736 7524 650748 7580
rect 650804 7524 650828 7580
rect 650884 7524 650908 7580
rect 650964 7524 650988 7580
rect 651044 7524 651056 7580
rect 650736 7500 651056 7524
rect 650736 7444 650748 7500
rect 650804 7444 650828 7500
rect 650884 7444 650908 7500
rect 650964 7444 650988 7500
rect 651044 7444 651056 7500
rect 650736 6381 651056 7444
rect 650736 6325 650748 6381
rect 650804 6325 650828 6381
rect 650884 6325 650908 6381
rect 650964 6325 650988 6381
rect 651044 6325 651056 6381
rect 650736 6301 651056 6325
rect 650736 6245 650748 6301
rect 650804 6245 650828 6301
rect 650884 6245 650908 6301
rect 650964 6245 650988 6301
rect 651044 6245 651056 6301
rect 650736 6221 651056 6245
rect 650736 6165 650748 6221
rect 650804 6165 650828 6221
rect 650884 6165 650908 6221
rect 650964 6165 650988 6221
rect 651044 6165 651056 6221
rect 650736 6141 651056 6165
rect 650736 6085 650748 6141
rect 650804 6085 650828 6141
rect 650884 6085 650908 6141
rect 650964 6085 650988 6141
rect 651044 6085 651056 6141
rect 650736 5022 651056 6085
rect 650736 4966 650748 5022
rect 650804 4966 650828 5022
rect 650884 4966 650908 5022
rect 650964 4966 650988 5022
rect 651044 4966 651056 5022
rect 650736 4942 651056 4966
rect 650736 4886 650748 4942
rect 650804 4886 650828 4942
rect 650884 4886 650908 4942
rect 650964 4886 650988 4942
rect 651044 4886 651056 4942
rect 650736 4862 651056 4886
rect 650736 4806 650748 4862
rect 650804 4806 650828 4862
rect 650884 4806 650908 4862
rect 650964 4806 650988 4862
rect 651044 4806 651056 4862
rect 650736 4782 651056 4806
rect 650736 4726 650748 4782
rect 650804 4726 650828 4782
rect 650884 4726 650908 4782
rect 650964 4726 650988 4782
rect 651044 4726 651056 4782
rect 650736 3663 651056 4726
rect 650736 3607 650748 3663
rect 650804 3607 650828 3663
rect 650884 3607 650908 3663
rect 650964 3607 650988 3663
rect 651044 3607 651056 3663
rect 650736 3583 651056 3607
rect 650736 3527 650748 3583
rect 650804 3527 650828 3583
rect 650884 3527 650908 3583
rect 650964 3527 650988 3583
rect 651044 3527 651056 3583
rect 650736 3503 651056 3527
rect 650736 3447 650748 3503
rect 650804 3447 650828 3503
rect 650884 3447 650908 3503
rect 650964 3447 650988 3503
rect 651044 3447 651056 3503
rect 650736 3423 651056 3447
rect 650736 3367 650748 3423
rect 650804 3367 650828 3423
rect 650884 3367 650908 3423
rect 650964 3367 650988 3423
rect 651044 3367 651056 3423
rect 650736 304 651056 3367
rect 650736 248 650748 304
rect 650804 248 650828 304
rect 650884 248 650908 304
rect 650964 248 650988 304
rect 651044 248 651056 304
rect 650736 224 651056 248
rect 650736 168 650748 224
rect 650804 168 650828 224
rect 650884 168 650908 224
rect 650964 168 650988 224
rect 651044 168 651056 224
rect 650736 144 651056 168
rect 650736 88 650748 144
rect 650804 88 650828 144
rect 650884 88 650908 144
rect 650964 88 650988 144
rect 651044 88 651056 144
rect 568404 8 568416 64
rect 568472 8 568496 64
rect 568552 8 568576 64
rect 568632 8 568656 64
rect 568712 8 568724 64
rect 568404 -4 568724 8
rect 573732 60 573784 66
rect 573732 2 573784 8
rect 618260 60 618312 66
rect 618260 2 618312 8
rect 650736 64 651056 88
rect 650736 8 650748 64
rect 650804 8 650828 64
rect 650884 8 650908 64
rect 650964 8 650988 64
rect 651044 8 651056 64
rect 650736 -4 651056 8
<< via2 >>
rect -1064 9728 -1008 9784
rect -984 9728 -928 9784
rect -904 9728 -848 9784
rect -824 9728 -768 9784
rect -1064 9648 -1008 9704
rect -984 9648 -928 9704
rect -904 9648 -848 9704
rect -824 9648 -768 9704
rect -1064 9568 -1008 9624
rect -984 9568 -928 9624
rect -904 9568 -848 9624
rect -824 9568 -768 9624
rect -1064 9488 -1008 9544
rect -984 9488 -928 9544
rect -904 9488 -848 9544
rect -824 9488 -768 9544
rect -1064 7684 -1008 7740
rect -984 7684 -928 7740
rect -904 7684 -848 7740
rect -824 7684 -768 7740
rect -1064 7604 -1008 7660
rect -984 7604 -928 7660
rect -904 7604 -848 7660
rect -824 7604 -768 7660
rect -1064 7524 -1008 7580
rect -984 7524 -928 7580
rect -904 7524 -848 7580
rect -824 7524 -768 7580
rect -1064 7444 -1008 7500
rect -984 7444 -928 7500
rect -904 7444 -848 7500
rect -824 7444 -768 7500
rect -1064 6325 -1008 6381
rect -984 6325 -928 6381
rect -904 6325 -848 6381
rect -824 6325 -768 6381
rect -1064 6245 -1008 6301
rect -984 6245 -928 6301
rect -904 6245 -848 6301
rect -824 6245 -768 6301
rect -1064 6165 -1008 6221
rect -984 6165 -928 6221
rect -904 6165 -848 6221
rect -824 6165 -768 6221
rect -1064 6085 -1008 6141
rect -984 6085 -928 6141
rect -904 6085 -848 6141
rect -824 6085 -768 6141
rect -1064 4966 -1008 5022
rect -984 4966 -928 5022
rect -904 4966 -848 5022
rect -824 4966 -768 5022
rect -1064 4886 -1008 4942
rect -984 4886 -928 4942
rect -904 4886 -848 4942
rect -824 4886 -768 4942
rect -1064 4806 -1008 4862
rect -984 4806 -928 4862
rect -904 4806 -848 4862
rect -824 4806 -768 4862
rect -1064 4726 -1008 4782
rect -984 4726 -928 4782
rect -904 4726 -848 4782
rect -824 4726 -768 4782
rect -1064 3607 -1008 3663
rect -984 3607 -928 3663
rect -904 3607 -848 3663
rect -824 3607 -768 3663
rect -1064 3527 -1008 3583
rect -984 3527 -928 3583
rect -904 3527 -848 3583
rect -824 3527 -768 3583
rect -1064 3447 -1008 3503
rect -984 3447 -928 3503
rect -904 3447 -848 3503
rect -824 3447 -768 3503
rect -1064 3367 -1008 3423
rect -984 3367 -928 3423
rect -904 3367 -848 3423
rect -824 3367 -768 3423
rect -404 9068 -348 9124
rect -324 9068 -268 9124
rect -244 9068 -188 9124
rect -164 9068 -108 9124
rect -404 8988 -348 9044
rect -324 8988 -268 9044
rect -244 8988 -188 9044
rect -164 8988 -108 9044
rect -404 8908 -348 8964
rect -324 8908 -268 8964
rect -244 8908 -188 8964
rect -164 8908 -108 8964
rect -404 8828 -348 8884
rect -324 8828 -268 8884
rect -244 8828 -188 8884
rect -164 8828 -108 8884
rect -404 7024 -348 7080
rect -324 7024 -268 7080
rect -244 7024 -188 7080
rect -164 7024 -108 7080
rect -404 6944 -348 7000
rect -324 6944 -268 7000
rect -244 6944 -188 7000
rect -164 6944 -108 7000
rect -404 6864 -348 6920
rect -324 6864 -268 6920
rect -244 6864 -188 6920
rect -164 6864 -108 6920
rect -404 6784 -348 6840
rect -324 6784 -268 6840
rect -244 6784 -188 6840
rect -164 6784 -108 6840
rect -404 5665 -348 5721
rect -324 5665 -268 5721
rect -244 5665 -188 5721
rect -164 5665 -108 5721
rect -404 5585 -348 5641
rect -324 5585 -268 5641
rect -244 5585 -188 5641
rect -164 5585 -108 5641
rect -404 5505 -348 5561
rect -324 5505 -268 5561
rect -244 5505 -188 5561
rect -164 5505 -108 5561
rect -404 5425 -348 5481
rect -324 5425 -268 5481
rect -244 5425 -188 5481
rect -164 5425 -108 5481
rect -404 4306 -348 4362
rect -324 4306 -268 4362
rect -244 4306 -188 4362
rect -164 4306 -108 4362
rect -404 4226 -348 4282
rect -324 4226 -268 4282
rect -244 4226 -188 4282
rect -164 4226 -108 4282
rect -404 4146 -348 4202
rect -324 4146 -268 4202
rect -244 4146 -188 4202
rect -164 4146 -108 4202
rect -404 4066 -348 4122
rect -324 4066 -268 4122
rect -244 4066 -188 4122
rect -164 4066 -108 4122
rect -404 2947 -348 3003
rect -324 2947 -268 3003
rect -244 2947 -188 3003
rect -164 2947 -108 3003
rect -404 2867 -348 2923
rect -324 2867 -268 2923
rect -244 2867 -188 2923
rect -164 2867 -108 2923
rect -404 2787 -348 2843
rect -324 2787 -268 2843
rect -244 2787 -188 2843
rect -164 2787 -108 2843
rect -404 2707 -348 2763
rect -324 2707 -268 2763
rect -244 2707 -188 2763
rect -164 2707 -108 2763
rect -404 908 -348 964
rect -324 908 -268 964
rect -244 908 -188 964
rect -164 908 -108 964
rect -404 828 -348 884
rect -324 828 -268 884
rect -244 828 -188 884
rect -164 828 -108 884
rect 28354 8064 28410 8120
rect 29182 7928 29238 7984
rect 81927 9068 81983 9124
rect 82007 9068 82063 9124
rect 82087 9068 82143 9124
rect 82167 9068 82223 9124
rect 81927 8988 81983 9044
rect 82007 8988 82063 9044
rect 82087 8988 82143 9044
rect 82167 8988 82223 9044
rect 81927 8908 81983 8964
rect 82007 8908 82063 8964
rect 82087 8908 82143 8964
rect 82167 8908 82223 8964
rect 81927 8828 81983 8884
rect 82007 8828 82063 8884
rect 82087 8828 82143 8884
rect 82167 8828 82223 8884
rect 30838 6568 30894 6624
rect 79322 5888 79378 5944
rect 81927 7046 81973 7080
rect 81973 7046 81983 7080
rect 82007 7046 82037 7080
rect 82037 7046 82049 7080
rect 82049 7046 82063 7080
rect 82087 7046 82101 7080
rect 82101 7046 82113 7080
rect 82113 7046 82143 7080
rect 82167 7046 82177 7080
rect 82177 7046 82223 7080
rect 81927 7024 81983 7046
rect 82007 7024 82063 7046
rect 82087 7024 82143 7046
rect 82167 7024 82223 7046
rect 81927 6944 81983 7000
rect 82007 6944 82063 7000
rect 82087 6944 82143 7000
rect 82167 6944 82223 7000
rect 81927 6864 81983 6920
rect 82007 6864 82063 6920
rect 82087 6864 82143 6920
rect 82167 6864 82223 6920
rect 81927 6784 81983 6840
rect 82007 6784 82063 6840
rect 82087 6784 82143 6840
rect 82167 6784 82223 6840
rect 82587 9728 82643 9784
rect 82667 9728 82723 9784
rect 82747 9728 82803 9784
rect 82827 9728 82883 9784
rect 82587 9648 82643 9704
rect 82667 9648 82723 9704
rect 82747 9648 82803 9704
rect 82827 9648 82883 9704
rect 82587 9568 82643 9624
rect 82667 9568 82723 9624
rect 82747 9568 82803 9624
rect 82827 9568 82883 9624
rect 82587 9488 82643 9544
rect 82667 9488 82723 9544
rect 82747 9488 82803 9544
rect 82827 9488 82883 9544
rect 82587 7684 82643 7740
rect 82667 7684 82723 7740
rect 82747 7684 82803 7740
rect 82827 7684 82883 7740
rect 82587 7642 82643 7660
rect 82667 7642 82723 7660
rect 82747 7642 82803 7660
rect 82827 7642 82883 7660
rect 82587 7604 82633 7642
rect 82633 7604 82643 7642
rect 82667 7604 82697 7642
rect 82697 7604 82709 7642
rect 82709 7604 82723 7642
rect 82747 7604 82761 7642
rect 82761 7604 82773 7642
rect 82773 7604 82803 7642
rect 82827 7604 82837 7642
rect 82837 7604 82883 7642
rect 82587 7524 82643 7580
rect 82667 7524 82723 7580
rect 82747 7524 82803 7580
rect 82827 7524 82883 7580
rect 82587 7444 82643 7500
rect 82667 7444 82723 7500
rect 82747 7444 82803 7500
rect 82827 7444 82883 7500
rect 81927 5665 81983 5721
rect 82007 5665 82063 5721
rect 82087 5665 82143 5721
rect 82167 5665 82223 5721
rect 81927 5585 81983 5641
rect 82007 5585 82063 5641
rect 82087 5585 82143 5641
rect 82167 5585 82223 5641
rect 81927 5505 81983 5561
rect 82007 5505 82063 5561
rect 82087 5505 82143 5561
rect 82167 5505 82223 5561
rect 81927 5425 81983 5481
rect 82007 5425 82063 5481
rect 82087 5425 82143 5481
rect 82167 5425 82223 5481
rect 81927 4306 81983 4362
rect 82007 4306 82063 4362
rect 82087 4306 82143 4362
rect 82167 4306 82223 4362
rect 81927 4226 81983 4282
rect 82007 4226 82063 4282
rect 82087 4226 82143 4282
rect 82167 4226 82223 4282
rect 81927 4146 81983 4202
rect 82007 4146 82063 4202
rect 82087 4146 82143 4202
rect 82167 4146 82223 4202
rect 81927 4066 81983 4122
rect 82007 4066 82063 4122
rect 82087 4066 82143 4122
rect 82167 4066 82223 4122
rect 81927 2947 81983 3003
rect 82007 2947 82063 3003
rect 82087 2947 82143 3003
rect 82167 2947 82223 3003
rect 82587 6325 82643 6381
rect 82667 6325 82723 6381
rect 82747 6325 82803 6381
rect 82827 6325 82883 6381
rect 82587 6245 82643 6301
rect 82667 6245 82723 6301
rect 82747 6245 82803 6301
rect 82827 6245 82883 6301
rect 82587 6165 82643 6221
rect 82667 6165 82723 6221
rect 82747 6165 82803 6221
rect 82827 6165 82883 6221
rect 82587 6085 82643 6141
rect 82667 6085 82723 6141
rect 82747 6085 82803 6141
rect 82827 6085 82883 6141
rect 82587 4966 82643 5022
rect 82667 4966 82723 5022
rect 82747 4966 82803 5022
rect 82827 4966 82883 5022
rect 82587 4886 82643 4942
rect 82667 4886 82723 4942
rect 82747 4886 82803 4942
rect 82827 4886 82883 4942
rect 82587 4806 82643 4862
rect 82667 4806 82723 4862
rect 82747 4806 82803 4862
rect 82827 4806 82883 4862
rect 82587 4726 82643 4782
rect 82667 4726 82723 4782
rect 82747 4726 82803 4782
rect 82827 4726 82883 4782
rect 82587 3607 82643 3663
rect 82667 3607 82723 3663
rect 82747 3607 82803 3663
rect 82827 3607 82883 3663
rect 82587 3527 82643 3583
rect 82667 3527 82723 3583
rect 82747 3527 82803 3583
rect 82827 3527 82883 3583
rect 82587 3447 82643 3503
rect 82667 3447 82723 3503
rect 82747 3447 82803 3503
rect 82827 3447 82883 3503
rect 82587 3367 82643 3423
rect 82667 3367 82723 3423
rect 82747 3367 82803 3423
rect 82827 3367 82883 3423
rect 81927 2867 81983 2923
rect 82007 2867 82063 2923
rect 82087 2867 82143 2923
rect 82167 2867 82223 2923
rect 81927 2787 81983 2843
rect 82007 2787 82063 2843
rect 82087 2787 82143 2843
rect 82167 2787 82223 2843
rect 81927 2746 81983 2763
rect 82007 2746 82063 2763
rect 82087 2746 82143 2763
rect 82167 2746 82223 2763
rect 81927 2707 81973 2746
rect 81973 2707 81983 2746
rect 82007 2707 82037 2746
rect 82037 2707 82049 2746
rect 82049 2707 82063 2746
rect 82087 2707 82101 2746
rect 82101 2707 82113 2746
rect 82113 2707 82143 2746
rect 82167 2707 82177 2746
rect 82177 2707 82223 2746
rect 81927 908 81983 964
rect 82007 908 82063 964
rect 82087 908 82143 964
rect 82167 908 82223 964
rect 81927 828 81983 884
rect 82007 828 82063 884
rect 82087 828 82143 884
rect 82167 828 82223 884
rect -404 748 -348 804
rect -324 748 -268 804
rect -244 748 -188 804
rect -164 748 -108 804
rect -404 668 -348 724
rect -324 668 -268 724
rect -244 668 -188 724
rect -164 668 -108 724
rect 81927 748 81983 804
rect 82007 748 82063 804
rect 82087 748 82143 804
rect 82167 748 82223 804
rect 81927 668 81983 724
rect 82007 668 82063 724
rect 82087 668 82143 724
rect 82167 668 82223 724
rect -1064 248 -1008 304
rect -984 248 -928 304
rect -904 248 -848 304
rect -824 248 -768 304
rect -1064 168 -1008 224
rect -984 168 -928 224
rect -904 168 -848 224
rect -824 168 -768 224
rect -1064 88 -1008 144
rect -984 88 -928 144
rect -904 88 -848 144
rect -824 88 -768 144
rect -1064 8 -1008 64
rect -984 8 -928 64
rect -904 8 -848 64
rect -824 8 -768 64
rect 243870 9068 243926 9124
rect 243950 9068 244006 9124
rect 244030 9068 244086 9124
rect 244110 9068 244166 9124
rect 243870 8988 243926 9044
rect 243950 8988 244006 9044
rect 244030 8988 244086 9044
rect 244110 8988 244166 9044
rect 243870 8908 243926 8964
rect 243950 8908 244006 8964
rect 244030 8908 244086 8964
rect 244110 8908 244166 8964
rect 243870 8828 243926 8884
rect 243950 8828 244006 8884
rect 244030 8828 244086 8884
rect 244110 8828 244166 8884
rect 121458 8064 121514 8120
rect 122838 7928 122894 7984
rect 124678 6568 124734 6624
rect 125506 6568 125562 6624
rect 154302 6568 154358 6624
rect 154486 6568 154542 6624
rect 126978 5888 127034 5944
rect 154302 5888 154358 5944
rect 166998 5888 167054 5944
rect 167182 5888 167238 5944
rect 244530 9728 244586 9784
rect 244610 9728 244666 9784
rect 244690 9728 244746 9784
rect 244770 9728 244826 9784
rect 244530 9648 244586 9704
rect 244610 9648 244666 9704
rect 244690 9648 244746 9704
rect 244770 9648 244826 9704
rect 244530 9568 244586 9624
rect 244610 9568 244666 9624
rect 244690 9568 244746 9624
rect 244770 9568 244826 9624
rect 244530 9488 244586 9544
rect 244610 9488 244666 9544
rect 244690 9488 244746 9544
rect 244770 9488 244826 9544
rect 244530 7684 244586 7740
rect 244610 7684 244666 7740
rect 244690 7684 244746 7740
rect 244770 7684 244826 7740
rect 244530 7642 244586 7660
rect 244610 7642 244666 7660
rect 244690 7642 244746 7660
rect 244770 7642 244826 7660
rect 244530 7604 244576 7642
rect 244576 7604 244586 7642
rect 244610 7604 244640 7642
rect 244640 7604 244652 7642
rect 244652 7604 244666 7642
rect 244690 7604 244704 7642
rect 244704 7604 244716 7642
rect 244716 7604 244746 7642
rect 244770 7604 244780 7642
rect 244780 7604 244826 7642
rect 244530 7524 244586 7580
rect 244610 7524 244666 7580
rect 244690 7524 244746 7580
rect 244770 7524 244826 7580
rect 244530 7444 244586 7500
rect 244610 7444 244666 7500
rect 244690 7444 244746 7500
rect 244770 7444 244826 7500
rect 243870 7046 243916 7080
rect 243916 7046 243926 7080
rect 243950 7046 243980 7080
rect 243980 7046 243992 7080
rect 243992 7046 244006 7080
rect 244030 7046 244044 7080
rect 244044 7046 244056 7080
rect 244056 7046 244086 7080
rect 244110 7046 244120 7080
rect 244120 7046 244166 7080
rect 243870 7024 243926 7046
rect 243950 7024 244006 7046
rect 244030 7024 244086 7046
rect 244110 7024 244166 7046
rect 243870 6944 243926 7000
rect 243950 6944 244006 7000
rect 244030 6944 244086 7000
rect 244110 6944 244166 7000
rect 243870 6864 243926 6920
rect 243950 6864 244006 6920
rect 244030 6864 244086 6920
rect 244110 6864 244166 6920
rect 243870 6784 243926 6840
rect 243950 6784 244006 6840
rect 244030 6784 244086 6840
rect 244110 6784 244166 6840
rect 243870 5665 243926 5721
rect 243950 5665 244006 5721
rect 244030 5665 244086 5721
rect 244110 5665 244166 5721
rect 243870 5585 243926 5641
rect 243950 5585 244006 5641
rect 244030 5585 244086 5641
rect 244110 5585 244166 5641
rect 243870 5505 243926 5561
rect 243950 5505 244006 5561
rect 244030 5505 244086 5561
rect 244110 5505 244166 5561
rect 243870 5425 243926 5481
rect 243950 5425 244006 5481
rect 244030 5425 244086 5481
rect 244110 5425 244166 5481
rect 243870 4306 243926 4362
rect 243950 4306 244006 4362
rect 244030 4306 244086 4362
rect 244110 4306 244166 4362
rect 243870 4226 243926 4282
rect 243950 4226 244006 4282
rect 244030 4226 244086 4282
rect 244110 4226 244166 4282
rect 243870 4146 243926 4202
rect 243950 4146 244006 4202
rect 244030 4146 244086 4202
rect 244110 4146 244166 4202
rect 243870 4066 243926 4122
rect 243950 4066 244006 4122
rect 244030 4066 244086 4122
rect 244110 4066 244166 4122
rect 243870 2947 243926 3003
rect 243950 2947 244006 3003
rect 244030 2947 244086 3003
rect 244110 2947 244166 3003
rect 243870 2867 243926 2923
rect 243950 2867 244006 2923
rect 244030 2867 244086 2923
rect 244110 2867 244166 2923
rect 243870 2787 243926 2843
rect 243950 2787 244006 2843
rect 244030 2787 244086 2843
rect 244110 2787 244166 2843
rect 243870 2746 243926 2763
rect 243950 2746 244006 2763
rect 244030 2746 244086 2763
rect 244110 2746 244166 2763
rect 243870 2707 243916 2746
rect 243916 2707 243926 2746
rect 243950 2707 243980 2746
rect 243980 2707 243992 2746
rect 243992 2707 244006 2746
rect 244030 2707 244044 2746
rect 244044 2707 244056 2746
rect 244056 2707 244086 2746
rect 244110 2707 244120 2746
rect 244120 2707 244166 2746
rect 243870 908 243926 964
rect 243950 908 244006 964
rect 244030 908 244086 964
rect 244110 908 244166 964
rect 243870 828 243926 884
rect 243950 828 244006 884
rect 244030 828 244086 884
rect 244110 828 244166 884
rect 82587 248 82643 304
rect 82667 248 82723 304
rect 82747 248 82803 304
rect 82827 248 82883 304
rect 82587 168 82643 224
rect 82667 168 82723 224
rect 82747 168 82803 224
rect 82827 168 82883 224
rect 82587 88 82643 144
rect 82667 88 82723 144
rect 82747 88 82803 144
rect 82827 88 82883 144
rect 82587 8 82643 64
rect 82667 8 82723 64
rect 82747 8 82803 64
rect 82827 8 82883 64
rect 243870 748 243926 804
rect 243950 748 244006 804
rect 244030 748 244086 804
rect 244110 748 244166 804
rect 243870 668 243926 724
rect 243950 668 244006 724
rect 244030 668 244086 724
rect 244110 668 244166 724
rect 405813 9068 405869 9124
rect 405893 9068 405949 9124
rect 405973 9068 406029 9124
rect 406053 9068 406109 9124
rect 405813 8988 405869 9044
rect 405893 8988 405949 9044
rect 405973 8988 406029 9044
rect 406053 8988 406109 9044
rect 405813 8908 405869 8964
rect 405893 8908 405949 8964
rect 405973 8908 406029 8964
rect 406053 8908 406109 8964
rect 405813 8828 405869 8884
rect 405893 8828 405949 8884
rect 405973 8828 406029 8884
rect 406053 8828 406109 8884
rect 244530 6325 244586 6381
rect 244610 6325 244666 6381
rect 244690 6325 244746 6381
rect 244770 6325 244826 6381
rect 244530 6245 244586 6301
rect 244610 6245 244666 6301
rect 244690 6245 244746 6301
rect 244770 6245 244826 6301
rect 244530 6165 244586 6221
rect 244610 6165 244666 6221
rect 244690 6165 244746 6221
rect 244770 6165 244826 6221
rect 244530 6085 244586 6141
rect 244610 6085 244666 6141
rect 244690 6085 244746 6141
rect 244770 6085 244826 6141
rect 246118 6604 246120 6624
rect 246120 6604 246172 6624
rect 246172 6604 246174 6624
rect 246118 6568 246174 6604
rect 246762 6568 246818 6624
rect 405813 7046 405859 7080
rect 405859 7046 405869 7080
rect 405893 7046 405923 7080
rect 405923 7046 405935 7080
rect 405935 7046 405949 7080
rect 405973 7046 405987 7080
rect 405987 7046 405999 7080
rect 405999 7046 406029 7080
rect 406053 7046 406063 7080
rect 406063 7046 406109 7080
rect 405813 7024 405869 7046
rect 405893 7024 405949 7046
rect 405973 7024 406029 7046
rect 406053 7024 406109 7046
rect 405813 6944 405869 7000
rect 405893 6944 405949 7000
rect 405973 6944 406029 7000
rect 406053 6944 406109 7000
rect 405813 6864 405869 6920
rect 405893 6864 405949 6920
rect 405973 6864 406029 6920
rect 406053 6864 406109 6920
rect 247590 5888 247646 5944
rect 244530 4966 244586 5022
rect 244610 4966 244666 5022
rect 244690 4966 244746 5022
rect 244770 4966 244826 5022
rect 244530 4886 244586 4942
rect 244610 4886 244666 4942
rect 244690 4886 244746 4942
rect 244770 4886 244826 4942
rect 244530 4806 244586 4862
rect 244610 4806 244666 4862
rect 244690 4806 244746 4862
rect 244770 4806 244826 4862
rect 244530 4726 244586 4782
rect 244610 4726 244666 4782
rect 244690 4726 244746 4782
rect 244770 4726 244826 4782
rect 405813 6784 405869 6840
rect 405893 6784 405949 6840
rect 405973 6784 406029 6840
rect 406053 6784 406109 6840
rect 244530 3607 244586 3663
rect 244610 3607 244666 3663
rect 244690 3607 244746 3663
rect 244770 3607 244826 3663
rect 244530 3527 244586 3583
rect 244610 3527 244666 3583
rect 244690 3527 244746 3583
rect 244770 3527 244826 3583
rect 244530 3447 244586 3503
rect 244610 3447 244666 3503
rect 244690 3447 244746 3503
rect 244770 3447 244826 3503
rect 244530 3367 244586 3423
rect 244610 3367 244666 3423
rect 244690 3367 244746 3423
rect 244770 3367 244826 3423
rect 405813 5665 405869 5721
rect 405893 5665 405949 5721
rect 405973 5665 406029 5721
rect 406053 5665 406109 5721
rect 405813 5585 405869 5641
rect 405893 5585 405949 5641
rect 405973 5585 406029 5641
rect 406053 5585 406109 5641
rect 405813 5505 405869 5561
rect 405893 5505 405949 5561
rect 405973 5505 406029 5561
rect 406053 5505 406109 5561
rect 405813 5425 405869 5481
rect 405893 5425 405949 5481
rect 405973 5425 406029 5481
rect 406053 5425 406109 5481
rect 406473 9728 406529 9784
rect 406553 9728 406609 9784
rect 406633 9728 406689 9784
rect 406713 9728 406769 9784
rect 406473 9648 406529 9704
rect 406553 9648 406609 9704
rect 406633 9648 406689 9704
rect 406713 9648 406769 9704
rect 406473 9568 406529 9624
rect 406553 9568 406609 9624
rect 406633 9568 406689 9624
rect 406713 9568 406769 9624
rect 406473 9488 406529 9544
rect 406553 9488 406609 9544
rect 406633 9488 406689 9544
rect 406713 9488 406769 9544
rect 406473 7684 406529 7740
rect 406553 7684 406609 7740
rect 406633 7684 406689 7740
rect 406713 7684 406769 7740
rect 406473 7642 406529 7660
rect 406553 7642 406609 7660
rect 406633 7642 406689 7660
rect 406713 7642 406769 7660
rect 406473 7604 406519 7642
rect 406519 7604 406529 7642
rect 406553 7604 406583 7642
rect 406583 7604 406595 7642
rect 406595 7604 406609 7642
rect 406633 7604 406647 7642
rect 406647 7604 406659 7642
rect 406659 7604 406689 7642
rect 406713 7604 406723 7642
rect 406723 7604 406769 7642
rect 406473 7524 406529 7580
rect 406553 7524 406609 7580
rect 406633 7524 406689 7580
rect 406713 7524 406769 7580
rect 406473 7444 406529 7500
rect 406553 7444 406609 7500
rect 406633 7444 406689 7500
rect 406713 7444 406769 7500
rect 406473 6325 406529 6381
rect 406553 6325 406609 6381
rect 406633 6325 406689 6381
rect 406713 6325 406769 6381
rect 406473 6245 406529 6301
rect 406553 6245 406609 6301
rect 406633 6245 406689 6301
rect 406713 6245 406769 6301
rect 406473 6165 406529 6221
rect 406553 6165 406609 6221
rect 406633 6165 406689 6221
rect 406713 6165 406769 6221
rect 406473 6085 406529 6141
rect 406553 6085 406609 6141
rect 406633 6085 406689 6141
rect 406713 6085 406769 6141
rect 567756 9068 567812 9124
rect 567836 9068 567892 9124
rect 567916 9068 567972 9124
rect 567996 9068 568052 9124
rect 567756 8988 567812 9044
rect 567836 8988 567892 9044
rect 567916 8988 567972 9044
rect 567996 8988 568052 9044
rect 567756 8908 567812 8964
rect 567836 8908 567892 8964
rect 567916 8908 567972 8964
rect 567996 8908 568052 8964
rect 567756 8828 567812 8884
rect 567836 8828 567892 8884
rect 567916 8828 567972 8884
rect 567996 8828 568052 8884
rect 567756 7046 567802 7080
rect 567802 7046 567812 7080
rect 567836 7046 567866 7080
rect 567866 7046 567878 7080
rect 567878 7046 567892 7080
rect 567916 7046 567930 7080
rect 567930 7046 567942 7080
rect 567942 7046 567972 7080
rect 567996 7046 568006 7080
rect 568006 7046 568052 7080
rect 567756 7024 567812 7046
rect 567836 7024 567892 7046
rect 567916 7024 567972 7046
rect 567996 7024 568052 7046
rect 567756 6944 567812 7000
rect 567836 6944 567892 7000
rect 567916 6944 567972 7000
rect 567996 6944 568052 7000
rect 567756 6864 567812 6920
rect 567836 6864 567892 6920
rect 567916 6864 567972 6920
rect 567996 6864 568052 6920
rect 567756 6784 567812 6840
rect 567836 6784 567892 6840
rect 567916 6784 567972 6840
rect 567996 6784 568052 6840
rect 567756 5665 567812 5721
rect 567836 5665 567892 5721
rect 567916 5665 567972 5721
rect 567996 5665 568052 5721
rect 567756 5585 567812 5641
rect 567836 5585 567892 5641
rect 567916 5585 567972 5641
rect 567996 5585 568052 5641
rect 567756 5505 567812 5561
rect 567836 5505 567892 5561
rect 567916 5505 567972 5561
rect 567996 5505 568052 5561
rect 567756 5425 567812 5481
rect 567836 5425 567892 5481
rect 567916 5425 567972 5481
rect 567996 5425 568052 5481
rect 406473 4966 406529 5022
rect 406553 4966 406609 5022
rect 406633 4966 406689 5022
rect 406713 4966 406769 5022
rect 406473 4886 406529 4942
rect 406553 4886 406609 4942
rect 406633 4886 406689 4942
rect 406713 4886 406769 4942
rect 406473 4806 406529 4862
rect 406553 4806 406609 4862
rect 406633 4806 406689 4862
rect 406713 4806 406769 4862
rect 406473 4726 406529 4782
rect 406553 4726 406609 4782
rect 406633 4726 406689 4782
rect 406713 4726 406769 4782
rect 405813 4306 405869 4362
rect 405893 4306 405949 4362
rect 405973 4306 406029 4362
rect 406053 4306 406109 4362
rect 405813 4226 405869 4282
rect 405893 4226 405949 4282
rect 405973 4226 406029 4282
rect 406053 4226 406109 4282
rect 405813 4146 405869 4202
rect 405893 4146 405949 4202
rect 405973 4146 406029 4202
rect 406053 4146 406109 4202
rect 405813 4066 405869 4122
rect 405893 4066 405949 4122
rect 405973 4066 406029 4122
rect 406053 4066 406109 4122
rect 406473 3607 406529 3663
rect 406553 3607 406609 3663
rect 406633 3607 406689 3663
rect 406713 3607 406769 3663
rect 406473 3527 406529 3583
rect 406553 3527 406609 3583
rect 406633 3527 406689 3583
rect 406713 3527 406769 3583
rect 406473 3447 406529 3503
rect 406553 3447 406609 3503
rect 406633 3447 406689 3503
rect 406713 3447 406769 3503
rect 405813 2947 405869 3003
rect 405893 2947 405949 3003
rect 405973 2947 406029 3003
rect 406053 2947 406109 3003
rect 244530 248 244586 304
rect 244610 248 244666 304
rect 244690 248 244746 304
rect 244770 248 244826 304
rect 244530 168 244586 224
rect 244610 168 244666 224
rect 244690 168 244746 224
rect 244770 168 244826 224
rect 244530 88 244586 144
rect 244610 88 244666 144
rect 244690 88 244746 144
rect 244770 88 244826 144
rect 405813 2867 405869 2923
rect 405893 2867 405949 2923
rect 405973 2867 406029 2923
rect 406053 2867 406109 2923
rect 405813 2787 405869 2843
rect 405893 2787 405949 2843
rect 405973 2787 406029 2843
rect 406053 2787 406109 2843
rect 405813 2746 405869 2763
rect 405893 2746 405949 2763
rect 405973 2746 406029 2763
rect 406053 2746 406109 2763
rect 405813 2707 405859 2746
rect 405859 2707 405869 2746
rect 405893 2707 405923 2746
rect 405923 2707 405935 2746
rect 405935 2707 405949 2746
rect 405973 2707 405987 2746
rect 405987 2707 405999 2746
rect 405999 2707 406029 2746
rect 406053 2707 406063 2746
rect 406063 2707 406109 2746
rect 405813 908 405869 964
rect 405893 908 405949 964
rect 405973 908 406029 964
rect 406053 908 406109 964
rect 405813 828 405869 884
rect 405893 828 405949 884
rect 405973 828 406029 884
rect 406053 828 406109 884
rect 405813 748 405869 804
rect 405893 748 405949 804
rect 405973 748 406029 804
rect 406053 748 406109 804
rect 405813 668 405869 724
rect 405893 668 405949 724
rect 405973 668 406029 724
rect 406053 668 406109 724
rect 244530 8 244586 64
rect 244610 8 244666 64
rect 244690 8 244746 64
rect 244770 8 244826 64
rect 406473 3367 406529 3423
rect 406553 3367 406609 3423
rect 406633 3367 406689 3423
rect 406713 3367 406769 3423
rect 567756 4306 567812 4362
rect 567836 4306 567892 4362
rect 567916 4306 567972 4362
rect 567996 4306 568052 4362
rect 567756 4226 567812 4282
rect 567836 4226 567892 4282
rect 567916 4226 567972 4282
rect 567996 4226 568052 4282
rect 567756 4146 567812 4202
rect 567836 4146 567892 4202
rect 567916 4146 567972 4202
rect 567996 4146 568052 4202
rect 567756 4066 567812 4122
rect 567836 4066 567892 4122
rect 567916 4066 567972 4122
rect 567996 4066 568052 4122
rect 406473 248 406529 304
rect 406553 248 406609 304
rect 406633 248 406689 304
rect 406713 248 406769 304
rect 406473 168 406529 224
rect 406553 168 406609 224
rect 406633 168 406689 224
rect 406713 168 406769 224
rect 406473 88 406529 144
rect 406553 88 406609 144
rect 406633 88 406689 144
rect 406713 88 406769 144
rect 567756 2947 567812 3003
rect 567836 2947 567892 3003
rect 567916 2947 567972 3003
rect 567996 2947 568052 3003
rect 567756 2867 567812 2923
rect 567836 2867 567892 2923
rect 567916 2867 567972 2923
rect 567996 2867 568052 2923
rect 567756 2787 567812 2843
rect 567836 2787 567892 2843
rect 567916 2787 567972 2843
rect 567996 2787 568052 2843
rect 567756 2746 567812 2763
rect 567836 2746 567892 2763
rect 567916 2746 567972 2763
rect 567996 2746 568052 2763
rect 567756 2707 567802 2746
rect 567802 2707 567812 2746
rect 567836 2707 567866 2746
rect 567866 2707 567878 2746
rect 567878 2707 567892 2746
rect 567916 2707 567930 2746
rect 567930 2707 567942 2746
rect 567942 2707 567972 2746
rect 567996 2707 568006 2746
rect 568006 2707 568052 2746
rect 567756 908 567812 964
rect 567836 908 567892 964
rect 567916 908 567972 964
rect 567996 908 568052 964
rect 567756 828 567812 884
rect 567836 828 567892 884
rect 567916 828 567972 884
rect 567996 828 568052 884
rect 567756 748 567812 804
rect 567836 748 567892 804
rect 567916 748 567972 804
rect 567996 748 568052 804
rect 567756 668 567812 724
rect 567836 668 567892 724
rect 567916 668 567972 724
rect 567996 668 568052 724
rect 406473 8 406529 64
rect 406553 8 406609 64
rect 406633 8 406689 64
rect 406713 8 406769 64
rect 568416 9728 568472 9784
rect 568496 9728 568552 9784
rect 568576 9728 568632 9784
rect 568656 9728 568712 9784
rect 568416 9648 568472 9704
rect 568496 9648 568552 9704
rect 568576 9648 568632 9704
rect 568656 9648 568712 9704
rect 568416 9568 568472 9624
rect 568496 9568 568552 9624
rect 568576 9568 568632 9624
rect 568656 9568 568712 9624
rect 568416 9488 568472 9544
rect 568496 9488 568552 9544
rect 568576 9488 568632 9544
rect 568656 9488 568712 9544
rect 650748 9728 650804 9784
rect 650828 9728 650884 9784
rect 650908 9728 650964 9784
rect 650988 9728 651044 9784
rect 650748 9648 650804 9704
rect 650828 9648 650884 9704
rect 650908 9648 650964 9704
rect 650988 9648 651044 9704
rect 650748 9568 650804 9624
rect 650828 9568 650884 9624
rect 650908 9568 650964 9624
rect 650988 9568 651044 9624
rect 650748 9488 650804 9544
rect 650828 9488 650884 9544
rect 650908 9488 650964 9544
rect 650988 9488 651044 9544
rect 568416 7684 568472 7740
rect 568496 7684 568552 7740
rect 568576 7684 568632 7740
rect 568656 7684 568712 7740
rect 568416 7642 568472 7660
rect 568496 7642 568552 7660
rect 568576 7642 568632 7660
rect 568656 7642 568712 7660
rect 568416 7604 568462 7642
rect 568462 7604 568472 7642
rect 568496 7604 568526 7642
rect 568526 7604 568538 7642
rect 568538 7604 568552 7642
rect 568576 7604 568590 7642
rect 568590 7604 568602 7642
rect 568602 7604 568632 7642
rect 568656 7604 568666 7642
rect 568666 7604 568712 7642
rect 568416 7524 568472 7580
rect 568496 7524 568552 7580
rect 568576 7524 568632 7580
rect 568656 7524 568712 7580
rect 568416 7444 568472 7500
rect 568496 7444 568552 7500
rect 568576 7444 568632 7500
rect 568656 7444 568712 7500
rect 568416 6325 568472 6381
rect 568496 6325 568552 6381
rect 568576 6325 568632 6381
rect 568656 6325 568712 6381
rect 568416 6245 568472 6301
rect 568496 6245 568552 6301
rect 568576 6245 568632 6301
rect 568656 6245 568712 6301
rect 568416 6165 568472 6221
rect 568496 6165 568552 6221
rect 568576 6165 568632 6221
rect 568656 6165 568712 6221
rect 568416 6085 568472 6141
rect 568496 6085 568552 6141
rect 568576 6085 568632 6141
rect 568656 6085 568712 6141
rect 568416 4966 568472 5022
rect 568496 4966 568552 5022
rect 568576 4966 568632 5022
rect 568656 4966 568712 5022
rect 568416 4886 568472 4942
rect 568496 4886 568552 4942
rect 568576 4886 568632 4942
rect 568656 4886 568712 4942
rect 568416 4806 568472 4862
rect 568496 4806 568552 4862
rect 568576 4806 568632 4862
rect 568656 4806 568712 4862
rect 568416 4726 568472 4782
rect 568496 4726 568552 4782
rect 568576 4726 568632 4782
rect 568656 4726 568712 4782
rect 650088 9068 650144 9124
rect 650168 9068 650224 9124
rect 650248 9068 650304 9124
rect 650328 9068 650384 9124
rect 650088 8988 650144 9044
rect 650168 8988 650224 9044
rect 650248 8988 650304 9044
rect 650328 8988 650384 9044
rect 650088 8908 650144 8964
rect 650168 8908 650224 8964
rect 650248 8908 650304 8964
rect 650328 8908 650384 8964
rect 650088 8828 650144 8884
rect 650168 8828 650224 8884
rect 650248 8828 650304 8884
rect 650328 8828 650384 8884
rect 650088 7024 650144 7080
rect 650168 7024 650224 7080
rect 650248 7024 650304 7080
rect 650328 7024 650384 7080
rect 650088 6944 650144 7000
rect 650168 6944 650224 7000
rect 650248 6944 650304 7000
rect 650328 6944 650384 7000
rect 650088 6864 650144 6920
rect 650168 6864 650224 6920
rect 650248 6864 650304 6920
rect 650328 6864 650384 6920
rect 650088 6784 650144 6840
rect 650168 6784 650224 6840
rect 650248 6784 650304 6840
rect 650328 6784 650384 6840
rect 650088 5665 650144 5721
rect 650168 5665 650224 5721
rect 650248 5665 650304 5721
rect 650328 5665 650384 5721
rect 650088 5585 650144 5641
rect 650168 5585 650224 5641
rect 650248 5585 650304 5641
rect 650328 5585 650384 5641
rect 650088 5505 650144 5561
rect 650168 5505 650224 5561
rect 650248 5505 650304 5561
rect 650328 5505 650384 5561
rect 650088 5425 650144 5481
rect 650168 5425 650224 5481
rect 650248 5425 650304 5481
rect 650328 5425 650384 5481
rect 650088 4306 650144 4362
rect 650168 4306 650224 4362
rect 650248 4306 650304 4362
rect 650328 4306 650384 4362
rect 650088 4226 650144 4282
rect 650168 4226 650224 4282
rect 650248 4226 650304 4282
rect 650328 4226 650384 4282
rect 650088 4146 650144 4202
rect 650168 4146 650224 4202
rect 650248 4146 650304 4202
rect 650328 4146 650384 4202
rect 650088 4066 650144 4122
rect 650168 4066 650224 4122
rect 650248 4066 650304 4122
rect 650328 4066 650384 4122
rect 568416 3607 568472 3663
rect 568496 3607 568552 3663
rect 568576 3607 568632 3663
rect 568656 3607 568712 3663
rect 568416 3527 568472 3583
rect 568496 3527 568552 3583
rect 568576 3527 568632 3583
rect 568656 3527 568712 3583
rect 568416 3447 568472 3503
rect 568496 3447 568552 3503
rect 568576 3447 568632 3503
rect 568656 3447 568712 3503
rect 568416 3367 568472 3423
rect 568496 3367 568552 3423
rect 568576 3367 568632 3423
rect 568656 3367 568712 3423
rect 650088 2947 650144 3003
rect 650168 2947 650224 3003
rect 650248 2947 650304 3003
rect 650328 2947 650384 3003
rect 650088 2867 650144 2923
rect 650168 2867 650224 2923
rect 650248 2867 650304 2923
rect 650328 2867 650384 2923
rect 650088 2787 650144 2843
rect 650168 2787 650224 2843
rect 650248 2787 650304 2843
rect 650328 2787 650384 2843
rect 650088 2707 650144 2763
rect 650168 2707 650224 2763
rect 650248 2707 650304 2763
rect 650328 2707 650384 2763
rect 568416 248 568472 304
rect 568496 248 568552 304
rect 568576 248 568632 304
rect 568656 248 568712 304
rect 568416 168 568472 224
rect 568496 168 568552 224
rect 568576 168 568632 224
rect 568656 168 568712 224
rect 568416 88 568472 144
rect 568496 88 568552 144
rect 568576 88 568632 144
rect 568656 88 568712 144
rect 650088 908 650144 964
rect 650168 908 650224 964
rect 650248 908 650304 964
rect 650328 908 650384 964
rect 650088 828 650144 884
rect 650168 828 650224 884
rect 650248 828 650304 884
rect 650328 828 650384 884
rect 650088 748 650144 804
rect 650168 748 650224 804
rect 650248 748 650304 804
rect 650328 748 650384 804
rect 650088 668 650144 724
rect 650168 668 650224 724
rect 650248 668 650304 724
rect 650328 668 650384 724
rect 650748 7684 650804 7740
rect 650828 7684 650884 7740
rect 650908 7684 650964 7740
rect 650988 7684 651044 7740
rect 650748 7604 650804 7660
rect 650828 7604 650884 7660
rect 650908 7604 650964 7660
rect 650988 7604 651044 7660
rect 650748 7524 650804 7580
rect 650828 7524 650884 7580
rect 650908 7524 650964 7580
rect 650988 7524 651044 7580
rect 650748 7444 650804 7500
rect 650828 7444 650884 7500
rect 650908 7444 650964 7500
rect 650988 7444 651044 7500
rect 650748 6325 650804 6381
rect 650828 6325 650884 6381
rect 650908 6325 650964 6381
rect 650988 6325 651044 6381
rect 650748 6245 650804 6301
rect 650828 6245 650884 6301
rect 650908 6245 650964 6301
rect 650988 6245 651044 6301
rect 650748 6165 650804 6221
rect 650828 6165 650884 6221
rect 650908 6165 650964 6221
rect 650988 6165 651044 6221
rect 650748 6085 650804 6141
rect 650828 6085 650884 6141
rect 650908 6085 650964 6141
rect 650988 6085 651044 6141
rect 650748 4966 650804 5022
rect 650828 4966 650884 5022
rect 650908 4966 650964 5022
rect 650988 4966 651044 5022
rect 650748 4886 650804 4942
rect 650828 4886 650884 4942
rect 650908 4886 650964 4942
rect 650988 4886 651044 4942
rect 650748 4806 650804 4862
rect 650828 4806 650884 4862
rect 650908 4806 650964 4862
rect 650988 4806 651044 4862
rect 650748 4726 650804 4782
rect 650828 4726 650884 4782
rect 650908 4726 650964 4782
rect 650988 4726 651044 4782
rect 650748 3607 650804 3663
rect 650828 3607 650884 3663
rect 650908 3607 650964 3663
rect 650988 3607 651044 3663
rect 650748 3527 650804 3583
rect 650828 3527 650884 3583
rect 650908 3527 650964 3583
rect 650988 3527 651044 3583
rect 650748 3447 650804 3503
rect 650828 3447 650884 3503
rect 650908 3447 650964 3503
rect 650988 3447 651044 3503
rect 650748 3367 650804 3423
rect 650828 3367 650884 3423
rect 650908 3367 650964 3423
rect 650988 3367 651044 3423
rect 650748 248 650804 304
rect 650828 248 650884 304
rect 650908 248 650964 304
rect 650988 248 651044 304
rect 650748 168 650804 224
rect 650828 168 650884 224
rect 650908 168 650964 224
rect 650988 168 651044 224
rect 650748 88 650804 144
rect 650828 88 650884 144
rect 650908 88 650964 144
rect 650988 88 651044 144
rect 568416 8 568472 64
rect 568496 8 568552 64
rect 568576 8 568632 64
rect 568656 8 568712 64
rect 650748 8 650804 64
rect 650828 8 650884 64
rect 650908 8 650964 64
rect 650988 8 651044 64
<< metal3 >>
rect -1076 9784 651056 9796
rect -1076 9728 -1064 9784
rect -1008 9728 -984 9784
rect -928 9728 -904 9784
rect -848 9728 -824 9784
rect -768 9728 82587 9784
rect 82643 9728 82667 9784
rect 82723 9728 82747 9784
rect 82803 9728 82827 9784
rect 82883 9728 244530 9784
rect 244586 9728 244610 9784
rect 244666 9728 244690 9784
rect 244746 9728 244770 9784
rect 244826 9728 406473 9784
rect 406529 9728 406553 9784
rect 406609 9728 406633 9784
rect 406689 9728 406713 9784
rect 406769 9728 568416 9784
rect 568472 9728 568496 9784
rect 568552 9728 568576 9784
rect 568632 9728 568656 9784
rect 568712 9728 650748 9784
rect 650804 9728 650828 9784
rect 650884 9728 650908 9784
rect 650964 9728 650988 9784
rect 651044 9728 651056 9784
rect -1076 9704 651056 9728
rect -1076 9648 -1064 9704
rect -1008 9648 -984 9704
rect -928 9648 -904 9704
rect -848 9648 -824 9704
rect -768 9648 82587 9704
rect 82643 9648 82667 9704
rect 82723 9648 82747 9704
rect 82803 9648 82827 9704
rect 82883 9648 244530 9704
rect 244586 9648 244610 9704
rect 244666 9648 244690 9704
rect 244746 9648 244770 9704
rect 244826 9648 406473 9704
rect 406529 9648 406553 9704
rect 406609 9648 406633 9704
rect 406689 9648 406713 9704
rect 406769 9648 568416 9704
rect 568472 9648 568496 9704
rect 568552 9648 568576 9704
rect 568632 9648 568656 9704
rect 568712 9648 650748 9704
rect 650804 9648 650828 9704
rect 650884 9648 650908 9704
rect 650964 9648 650988 9704
rect 651044 9648 651056 9704
rect -1076 9624 651056 9648
rect -1076 9568 -1064 9624
rect -1008 9568 -984 9624
rect -928 9568 -904 9624
rect -848 9568 -824 9624
rect -768 9568 82587 9624
rect 82643 9568 82667 9624
rect 82723 9568 82747 9624
rect 82803 9568 82827 9624
rect 82883 9568 244530 9624
rect 244586 9568 244610 9624
rect 244666 9568 244690 9624
rect 244746 9568 244770 9624
rect 244826 9568 406473 9624
rect 406529 9568 406553 9624
rect 406609 9568 406633 9624
rect 406689 9568 406713 9624
rect 406769 9568 568416 9624
rect 568472 9568 568496 9624
rect 568552 9568 568576 9624
rect 568632 9568 568656 9624
rect 568712 9568 650748 9624
rect 650804 9568 650828 9624
rect 650884 9568 650908 9624
rect 650964 9568 650988 9624
rect 651044 9568 651056 9624
rect -1076 9544 651056 9568
rect -1076 9488 -1064 9544
rect -1008 9488 -984 9544
rect -928 9488 -904 9544
rect -848 9488 -824 9544
rect -768 9488 82587 9544
rect 82643 9488 82667 9544
rect 82723 9488 82747 9544
rect 82803 9488 82827 9544
rect 82883 9488 244530 9544
rect 244586 9488 244610 9544
rect 244666 9488 244690 9544
rect 244746 9488 244770 9544
rect 244826 9488 406473 9544
rect 406529 9488 406553 9544
rect 406609 9488 406633 9544
rect 406689 9488 406713 9544
rect 406769 9488 568416 9544
rect 568472 9488 568496 9544
rect 568552 9488 568576 9544
rect 568632 9488 568656 9544
rect 568712 9488 650748 9544
rect 650804 9488 650828 9544
rect 650884 9488 650908 9544
rect 650964 9488 650988 9544
rect 651044 9488 651056 9544
rect -1076 9476 651056 9488
rect -416 9124 650396 9136
rect -416 9068 -404 9124
rect -348 9068 -324 9124
rect -268 9068 -244 9124
rect -188 9068 -164 9124
rect -108 9068 81927 9124
rect 81983 9068 82007 9124
rect 82063 9068 82087 9124
rect 82143 9068 82167 9124
rect 82223 9068 243870 9124
rect 243926 9068 243950 9124
rect 244006 9068 244030 9124
rect 244086 9068 244110 9124
rect 244166 9068 405813 9124
rect 405869 9068 405893 9124
rect 405949 9068 405973 9124
rect 406029 9068 406053 9124
rect 406109 9068 567756 9124
rect 567812 9068 567836 9124
rect 567892 9068 567916 9124
rect 567972 9068 567996 9124
rect 568052 9068 650088 9124
rect 650144 9068 650168 9124
rect 650224 9068 650248 9124
rect 650304 9068 650328 9124
rect 650384 9068 650396 9124
rect -416 9044 650396 9068
rect -416 8988 -404 9044
rect -348 8988 -324 9044
rect -268 8988 -244 9044
rect -188 8988 -164 9044
rect -108 8988 81927 9044
rect 81983 8988 82007 9044
rect 82063 8988 82087 9044
rect 82143 8988 82167 9044
rect 82223 8988 243870 9044
rect 243926 8988 243950 9044
rect 244006 8988 244030 9044
rect 244086 8988 244110 9044
rect 244166 8988 405813 9044
rect 405869 8988 405893 9044
rect 405949 8988 405973 9044
rect 406029 8988 406053 9044
rect 406109 8988 567756 9044
rect 567812 8988 567836 9044
rect 567892 8988 567916 9044
rect 567972 8988 567996 9044
rect 568052 8988 650088 9044
rect 650144 8988 650168 9044
rect 650224 8988 650248 9044
rect 650304 8988 650328 9044
rect 650384 8988 650396 9044
rect -416 8964 650396 8988
rect -416 8908 -404 8964
rect -348 8908 -324 8964
rect -268 8908 -244 8964
rect -188 8908 -164 8964
rect -108 8908 81927 8964
rect 81983 8908 82007 8964
rect 82063 8908 82087 8964
rect 82143 8908 82167 8964
rect 82223 8908 243870 8964
rect 243926 8908 243950 8964
rect 244006 8908 244030 8964
rect 244086 8908 244110 8964
rect 244166 8908 405813 8964
rect 405869 8908 405893 8964
rect 405949 8908 405973 8964
rect 406029 8908 406053 8964
rect 406109 8908 567756 8964
rect 567812 8908 567836 8964
rect 567892 8908 567916 8964
rect 567972 8908 567996 8964
rect 568052 8908 650088 8964
rect 650144 8908 650168 8964
rect 650224 8908 650248 8964
rect 650304 8908 650328 8964
rect 650384 8908 650396 8964
rect -416 8884 650396 8908
rect -416 8828 -404 8884
rect -348 8828 -324 8884
rect -268 8828 -244 8884
rect -188 8828 -164 8884
rect -108 8828 81927 8884
rect 81983 8828 82007 8884
rect 82063 8828 82087 8884
rect 82143 8828 82167 8884
rect 82223 8828 243870 8884
rect 243926 8828 243950 8884
rect 244006 8828 244030 8884
rect 244086 8828 244110 8884
rect 244166 8828 405813 8884
rect 405869 8828 405893 8884
rect 405949 8828 405973 8884
rect 406029 8828 406053 8884
rect 406109 8828 567756 8884
rect 567812 8828 567836 8884
rect 567892 8828 567916 8884
rect 567972 8828 567996 8884
rect 568052 8828 650088 8884
rect 650144 8828 650168 8884
rect 650224 8828 650248 8884
rect 650304 8828 650328 8884
rect 650384 8828 650396 8884
rect -416 8816 650396 8828
rect 28349 8122 28415 8125
rect 121453 8122 121519 8125
rect 28349 8120 121519 8122
rect 28349 8064 28354 8120
rect 28410 8064 121458 8120
rect 121514 8064 121519 8120
rect 28349 8062 121519 8064
rect 28349 8059 28415 8062
rect 121453 8059 121519 8062
rect 29177 7986 29243 7989
rect 122833 7986 122899 7989
rect 29177 7984 122899 7986
rect 29177 7928 29182 7984
rect 29238 7928 122838 7984
rect 122894 7928 122899 7984
rect 29177 7926 122899 7928
rect 29177 7923 29243 7926
rect 122833 7923 122899 7926
rect -1076 7740 651056 7752
rect -1076 7684 -1064 7740
rect -1008 7684 -984 7740
rect -928 7684 -904 7740
rect -848 7684 -824 7740
rect -768 7684 82587 7740
rect 82643 7684 82667 7740
rect 82723 7684 82747 7740
rect 82803 7684 82827 7740
rect 82883 7684 244530 7740
rect 244586 7684 244610 7740
rect 244666 7684 244690 7740
rect 244746 7684 244770 7740
rect 244826 7684 406473 7740
rect 406529 7684 406553 7740
rect 406609 7684 406633 7740
rect 406689 7684 406713 7740
rect 406769 7684 568416 7740
rect 568472 7684 568496 7740
rect 568552 7684 568576 7740
rect 568632 7684 568656 7740
rect 568712 7684 650748 7740
rect 650804 7684 650828 7740
rect 650884 7684 650908 7740
rect 650964 7684 650988 7740
rect 651044 7684 651056 7740
rect -1076 7660 651056 7684
rect -1076 7604 -1064 7660
rect -1008 7604 -984 7660
rect -928 7604 -904 7660
rect -848 7604 -824 7660
rect -768 7604 82587 7660
rect 82643 7604 82667 7660
rect 82723 7604 82747 7660
rect 82803 7604 82827 7660
rect 82883 7604 244530 7660
rect 244586 7604 244610 7660
rect 244666 7604 244690 7660
rect 244746 7604 244770 7660
rect 244826 7604 406473 7660
rect 406529 7604 406553 7660
rect 406609 7604 406633 7660
rect 406689 7604 406713 7660
rect 406769 7604 568416 7660
rect 568472 7604 568496 7660
rect 568552 7604 568576 7660
rect 568632 7604 568656 7660
rect 568712 7604 650748 7660
rect 650804 7604 650828 7660
rect 650884 7604 650908 7660
rect 650964 7604 650988 7660
rect 651044 7604 651056 7660
rect -1076 7580 651056 7604
rect -1076 7524 -1064 7580
rect -1008 7524 -984 7580
rect -928 7524 -904 7580
rect -848 7524 -824 7580
rect -768 7524 82587 7580
rect 82643 7524 82667 7580
rect 82723 7524 82747 7580
rect 82803 7524 82827 7580
rect 82883 7524 244530 7580
rect 244586 7524 244610 7580
rect 244666 7524 244690 7580
rect 244746 7524 244770 7580
rect 244826 7524 406473 7580
rect 406529 7524 406553 7580
rect 406609 7524 406633 7580
rect 406689 7524 406713 7580
rect 406769 7524 568416 7580
rect 568472 7524 568496 7580
rect 568552 7524 568576 7580
rect 568632 7524 568656 7580
rect 568712 7524 650748 7580
rect 650804 7524 650828 7580
rect 650884 7524 650908 7580
rect 650964 7524 650988 7580
rect 651044 7524 651056 7580
rect -1076 7500 651056 7524
rect -1076 7444 -1064 7500
rect -1008 7444 -984 7500
rect -928 7444 -904 7500
rect -848 7444 -824 7500
rect -768 7444 82587 7500
rect 82643 7444 82667 7500
rect 82723 7444 82747 7500
rect 82803 7444 82827 7500
rect 82883 7444 244530 7500
rect 244586 7444 244610 7500
rect 244666 7444 244690 7500
rect 244746 7444 244770 7500
rect 244826 7444 406473 7500
rect 406529 7444 406553 7500
rect 406609 7444 406633 7500
rect 406689 7444 406713 7500
rect 406769 7444 568416 7500
rect 568472 7444 568496 7500
rect 568552 7444 568576 7500
rect 568632 7444 568656 7500
rect 568712 7444 650748 7500
rect 650804 7444 650828 7500
rect 650884 7444 650908 7500
rect 650964 7444 650988 7500
rect 651044 7444 651056 7500
rect -1076 7432 651056 7444
rect -1076 7080 651056 7092
rect -1076 7024 -404 7080
rect -348 7024 -324 7080
rect -268 7024 -244 7080
rect -188 7024 -164 7080
rect -108 7024 81927 7080
rect 81983 7024 82007 7080
rect 82063 7024 82087 7080
rect 82143 7024 82167 7080
rect 82223 7024 243870 7080
rect 243926 7024 243950 7080
rect 244006 7024 244030 7080
rect 244086 7024 244110 7080
rect 244166 7024 405813 7080
rect 405869 7024 405893 7080
rect 405949 7024 405973 7080
rect 406029 7024 406053 7080
rect 406109 7024 567756 7080
rect 567812 7024 567836 7080
rect 567892 7024 567916 7080
rect 567972 7024 567996 7080
rect 568052 7024 650088 7080
rect 650144 7024 650168 7080
rect 650224 7024 650248 7080
rect 650304 7024 650328 7080
rect 650384 7024 651056 7080
rect -1076 7000 651056 7024
rect -1076 6944 -404 7000
rect -348 6944 -324 7000
rect -268 6944 -244 7000
rect -188 6944 -164 7000
rect -108 6944 81927 7000
rect 81983 6944 82007 7000
rect 82063 6944 82087 7000
rect 82143 6944 82167 7000
rect 82223 6944 243870 7000
rect 243926 6944 243950 7000
rect 244006 6944 244030 7000
rect 244086 6944 244110 7000
rect 244166 6944 405813 7000
rect 405869 6944 405893 7000
rect 405949 6944 405973 7000
rect 406029 6944 406053 7000
rect 406109 6944 567756 7000
rect 567812 6944 567836 7000
rect 567892 6944 567916 7000
rect 567972 6944 567996 7000
rect 568052 6944 650088 7000
rect 650144 6944 650168 7000
rect 650224 6944 650248 7000
rect 650304 6944 650328 7000
rect 650384 6944 651056 7000
rect -1076 6920 651056 6944
rect -1076 6864 -404 6920
rect -348 6864 -324 6920
rect -268 6864 -244 6920
rect -188 6864 -164 6920
rect -108 6864 81927 6920
rect 81983 6864 82007 6920
rect 82063 6864 82087 6920
rect 82143 6864 82167 6920
rect 82223 6864 243870 6920
rect 243926 6864 243950 6920
rect 244006 6864 244030 6920
rect 244086 6864 244110 6920
rect 244166 6864 405813 6920
rect 405869 6864 405893 6920
rect 405949 6864 405973 6920
rect 406029 6864 406053 6920
rect 406109 6864 567756 6920
rect 567812 6864 567836 6920
rect 567892 6864 567916 6920
rect 567972 6864 567996 6920
rect 568052 6864 650088 6920
rect 650144 6864 650168 6920
rect 650224 6864 650248 6920
rect 650304 6864 650328 6920
rect 650384 6864 651056 6920
rect -1076 6840 651056 6864
rect -1076 6784 -404 6840
rect -348 6784 -324 6840
rect -268 6784 -244 6840
rect -188 6784 -164 6840
rect -108 6784 81927 6840
rect 81983 6784 82007 6840
rect 82063 6784 82087 6840
rect 82143 6784 82167 6840
rect 82223 6784 243870 6840
rect 243926 6784 243950 6840
rect 244006 6784 244030 6840
rect 244086 6784 244110 6840
rect 244166 6784 405813 6840
rect 405869 6784 405893 6840
rect 405949 6784 405973 6840
rect 406029 6784 406053 6840
rect 406109 6784 567756 6840
rect 567812 6784 567836 6840
rect 567892 6784 567916 6840
rect 567972 6784 567996 6840
rect 568052 6784 650088 6840
rect 650144 6784 650168 6840
rect 650224 6784 650248 6840
rect 650304 6784 650328 6840
rect 650384 6784 651056 6840
rect -1076 6772 651056 6784
rect 30833 6626 30899 6629
rect 124673 6626 124739 6629
rect 30833 6624 124739 6626
rect 30833 6568 30838 6624
rect 30894 6568 124678 6624
rect 124734 6568 124739 6624
rect 30833 6566 124739 6568
rect 30833 6563 30899 6566
rect 124673 6563 124739 6566
rect 125501 6626 125567 6629
rect 154297 6626 154363 6629
rect 125501 6624 154363 6626
rect 125501 6568 125506 6624
rect 125562 6568 154302 6624
rect 154358 6568 154363 6624
rect 125501 6566 154363 6568
rect 125501 6563 125567 6566
rect 154297 6563 154363 6566
rect 154481 6626 154547 6629
rect 246113 6626 246179 6629
rect 246757 6626 246823 6629
rect 154481 6624 246823 6626
rect 154481 6568 154486 6624
rect 154542 6568 246118 6624
rect 246174 6568 246762 6624
rect 246818 6568 246823 6624
rect 154481 6566 246823 6568
rect 154481 6563 154547 6566
rect 246113 6563 246179 6566
rect 246757 6563 246823 6566
rect -1076 6381 651056 6393
rect -1076 6325 -1064 6381
rect -1008 6325 -984 6381
rect -928 6325 -904 6381
rect -848 6325 -824 6381
rect -768 6325 82587 6381
rect 82643 6325 82667 6381
rect 82723 6325 82747 6381
rect 82803 6325 82827 6381
rect 82883 6325 244530 6381
rect 244586 6325 244610 6381
rect 244666 6325 244690 6381
rect 244746 6325 244770 6381
rect 244826 6325 406473 6381
rect 406529 6325 406553 6381
rect 406609 6325 406633 6381
rect 406689 6325 406713 6381
rect 406769 6325 568416 6381
rect 568472 6325 568496 6381
rect 568552 6325 568576 6381
rect 568632 6325 568656 6381
rect 568712 6325 650748 6381
rect 650804 6325 650828 6381
rect 650884 6325 650908 6381
rect 650964 6325 650988 6381
rect 651044 6325 651056 6381
rect -1076 6301 651056 6325
rect -1076 6245 -1064 6301
rect -1008 6245 -984 6301
rect -928 6245 -904 6301
rect -848 6245 -824 6301
rect -768 6245 82587 6301
rect 82643 6245 82667 6301
rect 82723 6245 82747 6301
rect 82803 6245 82827 6301
rect 82883 6245 244530 6301
rect 244586 6245 244610 6301
rect 244666 6245 244690 6301
rect 244746 6245 244770 6301
rect 244826 6245 406473 6301
rect 406529 6245 406553 6301
rect 406609 6245 406633 6301
rect 406689 6245 406713 6301
rect 406769 6245 568416 6301
rect 568472 6245 568496 6301
rect 568552 6245 568576 6301
rect 568632 6245 568656 6301
rect 568712 6245 650748 6301
rect 650804 6245 650828 6301
rect 650884 6245 650908 6301
rect 650964 6245 650988 6301
rect 651044 6245 651056 6301
rect -1076 6221 651056 6245
rect -1076 6165 -1064 6221
rect -1008 6165 -984 6221
rect -928 6165 -904 6221
rect -848 6165 -824 6221
rect -768 6165 82587 6221
rect 82643 6165 82667 6221
rect 82723 6165 82747 6221
rect 82803 6165 82827 6221
rect 82883 6165 244530 6221
rect 244586 6165 244610 6221
rect 244666 6165 244690 6221
rect 244746 6165 244770 6221
rect 244826 6165 406473 6221
rect 406529 6165 406553 6221
rect 406609 6165 406633 6221
rect 406689 6165 406713 6221
rect 406769 6165 568416 6221
rect 568472 6165 568496 6221
rect 568552 6165 568576 6221
rect 568632 6165 568656 6221
rect 568712 6165 650748 6221
rect 650804 6165 650828 6221
rect 650884 6165 650908 6221
rect 650964 6165 650988 6221
rect 651044 6165 651056 6221
rect -1076 6141 651056 6165
rect -1076 6085 -1064 6141
rect -1008 6085 -984 6141
rect -928 6085 -904 6141
rect -848 6085 -824 6141
rect -768 6085 82587 6141
rect 82643 6085 82667 6141
rect 82723 6085 82747 6141
rect 82803 6085 82827 6141
rect 82883 6085 244530 6141
rect 244586 6085 244610 6141
rect 244666 6085 244690 6141
rect 244746 6085 244770 6141
rect 244826 6085 406473 6141
rect 406529 6085 406553 6141
rect 406609 6085 406633 6141
rect 406689 6085 406713 6141
rect 406769 6085 568416 6141
rect 568472 6085 568496 6141
rect 568552 6085 568576 6141
rect 568632 6085 568656 6141
rect 568712 6085 650748 6141
rect 650804 6085 650828 6141
rect 650884 6085 650908 6141
rect 650964 6085 650988 6141
rect 651044 6085 651056 6141
rect -1076 6073 651056 6085
rect 79317 5946 79383 5949
rect 126973 5946 127039 5949
rect 79317 5944 127039 5946
rect 79317 5888 79322 5944
rect 79378 5888 126978 5944
rect 127034 5888 127039 5944
rect 79317 5886 127039 5888
rect 79317 5883 79383 5886
rect 126973 5883 127039 5886
rect 154297 5946 154363 5949
rect 166993 5946 167059 5949
rect 154297 5944 167059 5946
rect 154297 5888 154302 5944
rect 154358 5888 166998 5944
rect 167054 5888 167059 5944
rect 154297 5886 167059 5888
rect 154297 5883 154363 5886
rect 166993 5883 167059 5886
rect 167177 5946 167243 5949
rect 247585 5946 247651 5949
rect 167177 5944 247651 5946
rect 167177 5888 167182 5944
rect 167238 5888 247590 5944
rect 247646 5888 247651 5944
rect 167177 5886 247651 5888
rect 167177 5883 167243 5886
rect 247585 5883 247651 5886
rect -1076 5721 651056 5733
rect -1076 5665 -404 5721
rect -348 5665 -324 5721
rect -268 5665 -244 5721
rect -188 5665 -164 5721
rect -108 5665 81927 5721
rect 81983 5665 82007 5721
rect 82063 5665 82087 5721
rect 82143 5665 82167 5721
rect 82223 5665 243870 5721
rect 243926 5665 243950 5721
rect 244006 5665 244030 5721
rect 244086 5665 244110 5721
rect 244166 5665 405813 5721
rect 405869 5665 405893 5721
rect 405949 5665 405973 5721
rect 406029 5665 406053 5721
rect 406109 5665 567756 5721
rect 567812 5665 567836 5721
rect 567892 5665 567916 5721
rect 567972 5665 567996 5721
rect 568052 5665 650088 5721
rect 650144 5665 650168 5721
rect 650224 5665 650248 5721
rect 650304 5665 650328 5721
rect 650384 5665 651056 5721
rect -1076 5641 651056 5665
rect -1076 5585 -404 5641
rect -348 5585 -324 5641
rect -268 5585 -244 5641
rect -188 5585 -164 5641
rect -108 5585 81927 5641
rect 81983 5585 82007 5641
rect 82063 5585 82087 5641
rect 82143 5585 82167 5641
rect 82223 5585 243870 5641
rect 243926 5585 243950 5641
rect 244006 5585 244030 5641
rect 244086 5585 244110 5641
rect 244166 5585 405813 5641
rect 405869 5585 405893 5641
rect 405949 5585 405973 5641
rect 406029 5585 406053 5641
rect 406109 5585 567756 5641
rect 567812 5585 567836 5641
rect 567892 5585 567916 5641
rect 567972 5585 567996 5641
rect 568052 5585 650088 5641
rect 650144 5585 650168 5641
rect 650224 5585 650248 5641
rect 650304 5585 650328 5641
rect 650384 5585 651056 5641
rect -1076 5561 651056 5585
rect -1076 5505 -404 5561
rect -348 5505 -324 5561
rect -268 5505 -244 5561
rect -188 5505 -164 5561
rect -108 5505 81927 5561
rect 81983 5505 82007 5561
rect 82063 5505 82087 5561
rect 82143 5505 82167 5561
rect 82223 5505 243870 5561
rect 243926 5505 243950 5561
rect 244006 5505 244030 5561
rect 244086 5505 244110 5561
rect 244166 5505 405813 5561
rect 405869 5505 405893 5561
rect 405949 5505 405973 5561
rect 406029 5505 406053 5561
rect 406109 5505 567756 5561
rect 567812 5505 567836 5561
rect 567892 5505 567916 5561
rect 567972 5505 567996 5561
rect 568052 5505 650088 5561
rect 650144 5505 650168 5561
rect 650224 5505 650248 5561
rect 650304 5505 650328 5561
rect 650384 5505 651056 5561
rect -1076 5481 651056 5505
rect -1076 5425 -404 5481
rect -348 5425 -324 5481
rect -268 5425 -244 5481
rect -188 5425 -164 5481
rect -108 5425 81927 5481
rect 81983 5425 82007 5481
rect 82063 5425 82087 5481
rect 82143 5425 82167 5481
rect 82223 5425 243870 5481
rect 243926 5425 243950 5481
rect 244006 5425 244030 5481
rect 244086 5425 244110 5481
rect 244166 5425 405813 5481
rect 405869 5425 405893 5481
rect 405949 5425 405973 5481
rect 406029 5425 406053 5481
rect 406109 5425 567756 5481
rect 567812 5425 567836 5481
rect 567892 5425 567916 5481
rect 567972 5425 567996 5481
rect 568052 5425 650088 5481
rect 650144 5425 650168 5481
rect 650224 5425 650248 5481
rect 650304 5425 650328 5481
rect 650384 5425 651056 5481
rect -1076 5413 651056 5425
rect -1076 5022 651056 5034
rect -1076 4966 -1064 5022
rect -1008 4966 -984 5022
rect -928 4966 -904 5022
rect -848 4966 -824 5022
rect -768 4966 82587 5022
rect 82643 4966 82667 5022
rect 82723 4966 82747 5022
rect 82803 4966 82827 5022
rect 82883 4966 244530 5022
rect 244586 4966 244610 5022
rect 244666 4966 244690 5022
rect 244746 4966 244770 5022
rect 244826 4966 406473 5022
rect 406529 4966 406553 5022
rect 406609 4966 406633 5022
rect 406689 4966 406713 5022
rect 406769 4966 568416 5022
rect 568472 4966 568496 5022
rect 568552 4966 568576 5022
rect 568632 4966 568656 5022
rect 568712 4966 650748 5022
rect 650804 4966 650828 5022
rect 650884 4966 650908 5022
rect 650964 4966 650988 5022
rect 651044 4966 651056 5022
rect -1076 4942 651056 4966
rect -1076 4886 -1064 4942
rect -1008 4886 -984 4942
rect -928 4886 -904 4942
rect -848 4886 -824 4942
rect -768 4886 82587 4942
rect 82643 4886 82667 4942
rect 82723 4886 82747 4942
rect 82803 4886 82827 4942
rect 82883 4886 244530 4942
rect 244586 4886 244610 4942
rect 244666 4886 244690 4942
rect 244746 4886 244770 4942
rect 244826 4886 406473 4942
rect 406529 4886 406553 4942
rect 406609 4886 406633 4942
rect 406689 4886 406713 4942
rect 406769 4886 568416 4942
rect 568472 4886 568496 4942
rect 568552 4886 568576 4942
rect 568632 4886 568656 4942
rect 568712 4886 650748 4942
rect 650804 4886 650828 4942
rect 650884 4886 650908 4942
rect 650964 4886 650988 4942
rect 651044 4886 651056 4942
rect -1076 4862 651056 4886
rect -1076 4806 -1064 4862
rect -1008 4806 -984 4862
rect -928 4806 -904 4862
rect -848 4806 -824 4862
rect -768 4806 82587 4862
rect 82643 4806 82667 4862
rect 82723 4806 82747 4862
rect 82803 4806 82827 4862
rect 82883 4806 244530 4862
rect 244586 4806 244610 4862
rect 244666 4806 244690 4862
rect 244746 4806 244770 4862
rect 244826 4806 406473 4862
rect 406529 4806 406553 4862
rect 406609 4806 406633 4862
rect 406689 4806 406713 4862
rect 406769 4806 568416 4862
rect 568472 4806 568496 4862
rect 568552 4806 568576 4862
rect 568632 4806 568656 4862
rect 568712 4806 650748 4862
rect 650804 4806 650828 4862
rect 650884 4806 650908 4862
rect 650964 4806 650988 4862
rect 651044 4806 651056 4862
rect -1076 4782 651056 4806
rect -1076 4726 -1064 4782
rect -1008 4726 -984 4782
rect -928 4726 -904 4782
rect -848 4726 -824 4782
rect -768 4726 82587 4782
rect 82643 4726 82667 4782
rect 82723 4726 82747 4782
rect 82803 4726 82827 4782
rect 82883 4726 244530 4782
rect 244586 4726 244610 4782
rect 244666 4726 244690 4782
rect 244746 4726 244770 4782
rect 244826 4726 406473 4782
rect 406529 4726 406553 4782
rect 406609 4726 406633 4782
rect 406689 4726 406713 4782
rect 406769 4726 568416 4782
rect 568472 4726 568496 4782
rect 568552 4726 568576 4782
rect 568632 4726 568656 4782
rect 568712 4726 650748 4782
rect 650804 4726 650828 4782
rect 650884 4726 650908 4782
rect 650964 4726 650988 4782
rect 651044 4726 651056 4782
rect -1076 4714 651056 4726
rect -1076 4362 651056 4374
rect -1076 4306 -404 4362
rect -348 4306 -324 4362
rect -268 4306 -244 4362
rect -188 4306 -164 4362
rect -108 4306 81927 4362
rect 81983 4306 82007 4362
rect 82063 4306 82087 4362
rect 82143 4306 82167 4362
rect 82223 4306 243870 4362
rect 243926 4306 243950 4362
rect 244006 4306 244030 4362
rect 244086 4306 244110 4362
rect 244166 4306 405813 4362
rect 405869 4306 405893 4362
rect 405949 4306 405973 4362
rect 406029 4306 406053 4362
rect 406109 4306 567756 4362
rect 567812 4306 567836 4362
rect 567892 4306 567916 4362
rect 567972 4306 567996 4362
rect 568052 4306 650088 4362
rect 650144 4306 650168 4362
rect 650224 4306 650248 4362
rect 650304 4306 650328 4362
rect 650384 4306 651056 4362
rect -1076 4282 651056 4306
rect -1076 4226 -404 4282
rect -348 4226 -324 4282
rect -268 4226 -244 4282
rect -188 4226 -164 4282
rect -108 4226 81927 4282
rect 81983 4226 82007 4282
rect 82063 4226 82087 4282
rect 82143 4226 82167 4282
rect 82223 4226 243870 4282
rect 243926 4226 243950 4282
rect 244006 4226 244030 4282
rect 244086 4226 244110 4282
rect 244166 4226 405813 4282
rect 405869 4226 405893 4282
rect 405949 4226 405973 4282
rect 406029 4226 406053 4282
rect 406109 4226 567756 4282
rect 567812 4226 567836 4282
rect 567892 4226 567916 4282
rect 567972 4226 567996 4282
rect 568052 4226 650088 4282
rect 650144 4226 650168 4282
rect 650224 4226 650248 4282
rect 650304 4226 650328 4282
rect 650384 4226 651056 4282
rect -1076 4202 651056 4226
rect -1076 4146 -404 4202
rect -348 4146 -324 4202
rect -268 4146 -244 4202
rect -188 4146 -164 4202
rect -108 4146 81927 4202
rect 81983 4146 82007 4202
rect 82063 4146 82087 4202
rect 82143 4146 82167 4202
rect 82223 4146 243870 4202
rect 243926 4146 243950 4202
rect 244006 4146 244030 4202
rect 244086 4146 244110 4202
rect 244166 4146 405813 4202
rect 405869 4146 405893 4202
rect 405949 4146 405973 4202
rect 406029 4146 406053 4202
rect 406109 4146 567756 4202
rect 567812 4146 567836 4202
rect 567892 4146 567916 4202
rect 567972 4146 567996 4202
rect 568052 4146 650088 4202
rect 650144 4146 650168 4202
rect 650224 4146 650248 4202
rect 650304 4146 650328 4202
rect 650384 4146 651056 4202
rect -1076 4122 651056 4146
rect -1076 4066 -404 4122
rect -348 4066 -324 4122
rect -268 4066 -244 4122
rect -188 4066 -164 4122
rect -108 4066 81927 4122
rect 81983 4066 82007 4122
rect 82063 4066 82087 4122
rect 82143 4066 82167 4122
rect 82223 4066 243870 4122
rect 243926 4066 243950 4122
rect 244006 4066 244030 4122
rect 244086 4066 244110 4122
rect 244166 4066 405813 4122
rect 405869 4066 405893 4122
rect 405949 4066 405973 4122
rect 406029 4066 406053 4122
rect 406109 4066 567756 4122
rect 567812 4066 567836 4122
rect 567892 4066 567916 4122
rect 567972 4066 567996 4122
rect 568052 4066 650088 4122
rect 650144 4066 650168 4122
rect 650224 4066 650248 4122
rect 650304 4066 650328 4122
rect 650384 4066 651056 4122
rect -1076 4054 651056 4066
rect -1076 3663 651056 3675
rect -1076 3607 -1064 3663
rect -1008 3607 -984 3663
rect -928 3607 -904 3663
rect -848 3607 -824 3663
rect -768 3607 82587 3663
rect 82643 3607 82667 3663
rect 82723 3607 82747 3663
rect 82803 3607 82827 3663
rect 82883 3607 244530 3663
rect 244586 3607 244610 3663
rect 244666 3607 244690 3663
rect 244746 3607 244770 3663
rect 244826 3607 406473 3663
rect 406529 3607 406553 3663
rect 406609 3607 406633 3663
rect 406689 3607 406713 3663
rect 406769 3607 568416 3663
rect 568472 3607 568496 3663
rect 568552 3607 568576 3663
rect 568632 3607 568656 3663
rect 568712 3607 650748 3663
rect 650804 3607 650828 3663
rect 650884 3607 650908 3663
rect 650964 3607 650988 3663
rect 651044 3607 651056 3663
rect -1076 3583 651056 3607
rect -1076 3527 -1064 3583
rect -1008 3527 -984 3583
rect -928 3527 -904 3583
rect -848 3527 -824 3583
rect -768 3527 82587 3583
rect 82643 3527 82667 3583
rect 82723 3527 82747 3583
rect 82803 3527 82827 3583
rect 82883 3527 244530 3583
rect 244586 3527 244610 3583
rect 244666 3527 244690 3583
rect 244746 3527 244770 3583
rect 244826 3527 406473 3583
rect 406529 3527 406553 3583
rect 406609 3527 406633 3583
rect 406689 3527 406713 3583
rect 406769 3527 568416 3583
rect 568472 3527 568496 3583
rect 568552 3527 568576 3583
rect 568632 3527 568656 3583
rect 568712 3527 650748 3583
rect 650804 3527 650828 3583
rect 650884 3527 650908 3583
rect 650964 3527 650988 3583
rect 651044 3527 651056 3583
rect -1076 3503 651056 3527
rect -1076 3447 -1064 3503
rect -1008 3447 -984 3503
rect -928 3447 -904 3503
rect -848 3447 -824 3503
rect -768 3447 82587 3503
rect 82643 3447 82667 3503
rect 82723 3447 82747 3503
rect 82803 3447 82827 3503
rect 82883 3447 244530 3503
rect 244586 3447 244610 3503
rect 244666 3447 244690 3503
rect 244746 3447 244770 3503
rect 244826 3447 406473 3503
rect 406529 3447 406553 3503
rect 406609 3447 406633 3503
rect 406689 3447 406713 3503
rect 406769 3447 568416 3503
rect 568472 3447 568496 3503
rect 568552 3447 568576 3503
rect 568632 3447 568656 3503
rect 568712 3447 650748 3503
rect 650804 3447 650828 3503
rect 650884 3447 650908 3503
rect 650964 3447 650988 3503
rect 651044 3447 651056 3503
rect -1076 3423 651056 3447
rect -1076 3367 -1064 3423
rect -1008 3367 -984 3423
rect -928 3367 -904 3423
rect -848 3367 -824 3423
rect -768 3367 82587 3423
rect 82643 3367 82667 3423
rect 82723 3367 82747 3423
rect 82803 3367 82827 3423
rect 82883 3367 244530 3423
rect 244586 3367 244610 3423
rect 244666 3367 244690 3423
rect 244746 3367 244770 3423
rect 244826 3367 406473 3423
rect 406529 3367 406553 3423
rect 406609 3367 406633 3423
rect 406689 3367 406713 3423
rect 406769 3367 568416 3423
rect 568472 3367 568496 3423
rect 568552 3367 568576 3423
rect 568632 3367 568656 3423
rect 568712 3367 650748 3423
rect 650804 3367 650828 3423
rect 650884 3367 650908 3423
rect 650964 3367 650988 3423
rect 651044 3367 651056 3423
rect -1076 3355 651056 3367
rect -1076 3003 651056 3015
rect -1076 2947 -404 3003
rect -348 2947 -324 3003
rect -268 2947 -244 3003
rect -188 2947 -164 3003
rect -108 2947 81927 3003
rect 81983 2947 82007 3003
rect 82063 2947 82087 3003
rect 82143 2947 82167 3003
rect 82223 2947 243870 3003
rect 243926 2947 243950 3003
rect 244006 2947 244030 3003
rect 244086 2947 244110 3003
rect 244166 2947 405813 3003
rect 405869 2947 405893 3003
rect 405949 2947 405973 3003
rect 406029 2947 406053 3003
rect 406109 2947 567756 3003
rect 567812 2947 567836 3003
rect 567892 2947 567916 3003
rect 567972 2947 567996 3003
rect 568052 2947 650088 3003
rect 650144 2947 650168 3003
rect 650224 2947 650248 3003
rect 650304 2947 650328 3003
rect 650384 2947 651056 3003
rect -1076 2923 651056 2947
rect -1076 2867 -404 2923
rect -348 2867 -324 2923
rect -268 2867 -244 2923
rect -188 2867 -164 2923
rect -108 2867 81927 2923
rect 81983 2867 82007 2923
rect 82063 2867 82087 2923
rect 82143 2867 82167 2923
rect 82223 2867 243870 2923
rect 243926 2867 243950 2923
rect 244006 2867 244030 2923
rect 244086 2867 244110 2923
rect 244166 2867 405813 2923
rect 405869 2867 405893 2923
rect 405949 2867 405973 2923
rect 406029 2867 406053 2923
rect 406109 2867 567756 2923
rect 567812 2867 567836 2923
rect 567892 2867 567916 2923
rect 567972 2867 567996 2923
rect 568052 2867 650088 2923
rect 650144 2867 650168 2923
rect 650224 2867 650248 2923
rect 650304 2867 650328 2923
rect 650384 2867 651056 2923
rect -1076 2843 651056 2867
rect -1076 2787 -404 2843
rect -348 2787 -324 2843
rect -268 2787 -244 2843
rect -188 2787 -164 2843
rect -108 2787 81927 2843
rect 81983 2787 82007 2843
rect 82063 2787 82087 2843
rect 82143 2787 82167 2843
rect 82223 2787 243870 2843
rect 243926 2787 243950 2843
rect 244006 2787 244030 2843
rect 244086 2787 244110 2843
rect 244166 2787 405813 2843
rect 405869 2787 405893 2843
rect 405949 2787 405973 2843
rect 406029 2787 406053 2843
rect 406109 2787 567756 2843
rect 567812 2787 567836 2843
rect 567892 2787 567916 2843
rect 567972 2787 567996 2843
rect 568052 2787 650088 2843
rect 650144 2787 650168 2843
rect 650224 2787 650248 2843
rect 650304 2787 650328 2843
rect 650384 2787 651056 2843
rect -1076 2763 651056 2787
rect -1076 2707 -404 2763
rect -348 2707 -324 2763
rect -268 2707 -244 2763
rect -188 2707 -164 2763
rect -108 2707 81927 2763
rect 81983 2707 82007 2763
rect 82063 2707 82087 2763
rect 82143 2707 82167 2763
rect 82223 2707 243870 2763
rect 243926 2707 243950 2763
rect 244006 2707 244030 2763
rect 244086 2707 244110 2763
rect 244166 2707 405813 2763
rect 405869 2707 405893 2763
rect 405949 2707 405973 2763
rect 406029 2707 406053 2763
rect 406109 2707 567756 2763
rect 567812 2707 567836 2763
rect 567892 2707 567916 2763
rect 567972 2707 567996 2763
rect 568052 2707 650088 2763
rect 650144 2707 650168 2763
rect 650224 2707 650248 2763
rect 650304 2707 650328 2763
rect 650384 2707 651056 2763
rect -1076 2695 651056 2707
rect -416 964 650396 976
rect -416 908 -404 964
rect -348 908 -324 964
rect -268 908 -244 964
rect -188 908 -164 964
rect -108 908 81927 964
rect 81983 908 82007 964
rect 82063 908 82087 964
rect 82143 908 82167 964
rect 82223 908 243870 964
rect 243926 908 243950 964
rect 244006 908 244030 964
rect 244086 908 244110 964
rect 244166 908 405813 964
rect 405869 908 405893 964
rect 405949 908 405973 964
rect 406029 908 406053 964
rect 406109 908 567756 964
rect 567812 908 567836 964
rect 567892 908 567916 964
rect 567972 908 567996 964
rect 568052 908 650088 964
rect 650144 908 650168 964
rect 650224 908 650248 964
rect 650304 908 650328 964
rect 650384 908 650396 964
rect -416 884 650396 908
rect -416 828 -404 884
rect -348 828 -324 884
rect -268 828 -244 884
rect -188 828 -164 884
rect -108 828 81927 884
rect 81983 828 82007 884
rect 82063 828 82087 884
rect 82143 828 82167 884
rect 82223 828 243870 884
rect 243926 828 243950 884
rect 244006 828 244030 884
rect 244086 828 244110 884
rect 244166 828 405813 884
rect 405869 828 405893 884
rect 405949 828 405973 884
rect 406029 828 406053 884
rect 406109 828 567756 884
rect 567812 828 567836 884
rect 567892 828 567916 884
rect 567972 828 567996 884
rect 568052 828 650088 884
rect 650144 828 650168 884
rect 650224 828 650248 884
rect 650304 828 650328 884
rect 650384 828 650396 884
rect -416 804 650396 828
rect -416 748 -404 804
rect -348 748 -324 804
rect -268 748 -244 804
rect -188 748 -164 804
rect -108 748 81927 804
rect 81983 748 82007 804
rect 82063 748 82087 804
rect 82143 748 82167 804
rect 82223 748 243870 804
rect 243926 748 243950 804
rect 244006 748 244030 804
rect 244086 748 244110 804
rect 244166 748 405813 804
rect 405869 748 405893 804
rect 405949 748 405973 804
rect 406029 748 406053 804
rect 406109 748 567756 804
rect 567812 748 567836 804
rect 567892 748 567916 804
rect 567972 748 567996 804
rect 568052 748 650088 804
rect 650144 748 650168 804
rect 650224 748 650248 804
rect 650304 748 650328 804
rect 650384 748 650396 804
rect -416 724 650396 748
rect -416 668 -404 724
rect -348 668 -324 724
rect -268 668 -244 724
rect -188 668 -164 724
rect -108 668 81927 724
rect 81983 668 82007 724
rect 82063 668 82087 724
rect 82143 668 82167 724
rect 82223 668 243870 724
rect 243926 668 243950 724
rect 244006 668 244030 724
rect 244086 668 244110 724
rect 244166 668 405813 724
rect 405869 668 405893 724
rect 405949 668 405973 724
rect 406029 668 406053 724
rect 406109 668 567756 724
rect 567812 668 567836 724
rect 567892 668 567916 724
rect 567972 668 567996 724
rect 568052 668 650088 724
rect 650144 668 650168 724
rect 650224 668 650248 724
rect 650304 668 650328 724
rect 650384 668 650396 724
rect -416 656 650396 668
rect -1076 304 651056 316
rect -1076 248 -1064 304
rect -1008 248 -984 304
rect -928 248 -904 304
rect -848 248 -824 304
rect -768 248 82587 304
rect 82643 248 82667 304
rect 82723 248 82747 304
rect 82803 248 82827 304
rect 82883 248 244530 304
rect 244586 248 244610 304
rect 244666 248 244690 304
rect 244746 248 244770 304
rect 244826 248 406473 304
rect 406529 248 406553 304
rect 406609 248 406633 304
rect 406689 248 406713 304
rect 406769 248 568416 304
rect 568472 248 568496 304
rect 568552 248 568576 304
rect 568632 248 568656 304
rect 568712 248 650748 304
rect 650804 248 650828 304
rect 650884 248 650908 304
rect 650964 248 650988 304
rect 651044 248 651056 304
rect -1076 224 651056 248
rect -1076 168 -1064 224
rect -1008 168 -984 224
rect -928 168 -904 224
rect -848 168 -824 224
rect -768 168 82587 224
rect 82643 168 82667 224
rect 82723 168 82747 224
rect 82803 168 82827 224
rect 82883 168 244530 224
rect 244586 168 244610 224
rect 244666 168 244690 224
rect 244746 168 244770 224
rect 244826 168 406473 224
rect 406529 168 406553 224
rect 406609 168 406633 224
rect 406689 168 406713 224
rect 406769 168 568416 224
rect 568472 168 568496 224
rect 568552 168 568576 224
rect 568632 168 568656 224
rect 568712 168 650748 224
rect 650804 168 650828 224
rect 650884 168 650908 224
rect 650964 168 650988 224
rect 651044 168 651056 224
rect -1076 144 651056 168
rect -1076 88 -1064 144
rect -1008 88 -984 144
rect -928 88 -904 144
rect -848 88 -824 144
rect -768 88 82587 144
rect 82643 88 82667 144
rect 82723 88 82747 144
rect 82803 88 82827 144
rect 82883 88 244530 144
rect 244586 88 244610 144
rect 244666 88 244690 144
rect 244746 88 244770 144
rect 244826 88 406473 144
rect 406529 88 406553 144
rect 406609 88 406633 144
rect 406689 88 406713 144
rect 406769 88 568416 144
rect 568472 88 568496 144
rect 568552 88 568576 144
rect 568632 88 568656 144
rect 568712 88 650748 144
rect 650804 88 650828 144
rect 650884 88 650908 144
rect 650964 88 650988 144
rect 651044 88 651056 144
rect -1076 64 651056 88
rect -1076 8 -1064 64
rect -1008 8 -984 64
rect -928 8 -904 64
rect -848 8 -824 64
rect -768 8 82587 64
rect 82643 8 82667 64
rect 82723 8 82747 64
rect 82803 8 82827 64
rect 82883 8 244530 64
rect 244586 8 244610 64
rect 244666 8 244690 64
rect 244746 8 244770 64
rect 244826 8 406473 64
rect 406529 8 406553 64
rect 406609 8 406633 64
rect 406689 8 406713 64
rect 406769 8 568416 64
rect 568472 8 568496 64
rect 568552 8 568576 64
rect 568632 8 568656 64
rect 568712 8 650748 64
rect 650804 8 650828 64
rect 650884 8 650908 64
rect 650964 8 650988 64
rect 651044 8 651056 64
rect -1076 -4 651056 8
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[0\].u_buf_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 1748 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[1\].u_buf_A
timestamp 1676037725
transform 1 0 17940 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[2\].u_buf_A
timestamp 1676037725
transform 1 0 32476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[3\].u_buf_A
timestamp 1676037725
transform -1 0 48116 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[4\].u_buf_A
timestamp 1676037725
transform 1 0 63388 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[5\].u_buf_A
timestamp 1676037725
transform 1 0 78844 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[6\].u_buf_A
timestamp 1676037725
transform -1 0 94484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[7\].u_buf_A
timestamp 1676037725
transform 1 0 109756 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[8\].u_buf_A
timestamp 1676037725
transform 1 0 125212 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[9\].u_buf_A
timestamp 1676037725
transform -1 0 140852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[10\].u_buf_A
timestamp 1676037725
transform 1 0 156124 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[11\].u_buf_A
timestamp 1676037725
transform 1 0 171580 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[12\].u_buf_A
timestamp 1676037725
transform -1 0 187036 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[13\].u_buf_A
timestamp 1676037725
transform 1 0 202492 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[14\].u_buf_A
timestamp 1676037725
transform 1 0 217948 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[15\].u_buf_A
timestamp 1676037725
transform -1 0 233588 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[16\].u_buf_A
timestamp 1676037725
transform 1 0 248860 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[17\].u_buf_A
timestamp 1676037725
transform 1 0 264316 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[18\].u_buf_A
timestamp 1676037725
transform -1 0 279772 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[19\].u_buf_A
timestamp 1676037725
transform 1 0 295228 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[20\].u_buf_A
timestamp 1676037725
transform 1 0 310684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[21\].u_buf_A
timestamp 1676037725
transform -1 0 326324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[22\].u_buf_A
timestamp 1676037725
transform 1 0 341596 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[23\].u_buf_A
timestamp 1676037725
transform 1 0 357052 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[24\].u_buf_A
timestamp 1676037725
transform -1 0 372692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[25\].u_buf_A
timestamp 1676037725
transform 1 0 387964 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[26\].u_buf_A
timestamp 1676037725
transform 1 0 402592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[27\].u_buf_A
timestamp 1676037725
transform -1 0 419980 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[28\].u_buf_A
timestamp 1676037725
transform 1 0 434332 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[29\].u_buf_A
timestamp 1676037725
transform 1 0 449788 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[30\].u_buf_A
timestamp 1676037725
transform -1 0 465428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[31\].u_buf_A
timestamp 1676037725
transform 1 0 480700 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[32\].u_buf_A
timestamp 1676037725
transform 1 0 496156 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[33\].u_buf_A
timestamp 1676037725
transform -1 0 512716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[34\].u_buf_A
timestamp 1676037725
transform 1 0 527068 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[35\].u_buf_A
timestamp 1676037725
transform 1 0 542524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[36\].u_buf_A
timestamp 1676037725
transform -1 0 558164 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[37\].u_buf_A
timestamp 1676037725
transform 1 0 573436 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[38\].u_buf_A
timestamp 1676037725
transform 1 0 588892 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[39\].u_buf_A
timestamp 1676037725
transform -1 0 605452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[40\].u_buf_A
timestamp 1676037725
transform 1 0 619804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[41\].u_buf_A
timestamp 1676037725
transform 1 0 635260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire1_A
timestamp 1676037725
transform -1 0 113252 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire2_A
timestamp 1676037725
transform 1 0 125764 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire3_A
timestamp 1676037725
transform 1 0 220340 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire4_A
timestamp 1676037725
transform 1 0 313628 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire5_A
timestamp 1676037725
transform 1 0 407192 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire6_A
timestamp 1676037725
transform 1 0 501124 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire8_A
timestamp 1676037725
transform -1 0 124384 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire9_A
timestamp 1676037725
transform -1 0 219328 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire10_A
timestamp 1676037725
transform 1 0 311788 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire11_A
timestamp 1676037725
transform -1 0 405996 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire12_A
timestamp 1676037725
transform -1 0 499928 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire13_A
timestamp 1676037725
transform -1 0 123004 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire14_A
timestamp 1676037725
transform 1 0 217764 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire15_A
timestamp 1676037725
transform 1 0 310960 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire16_A
timestamp 1676037725
transform -1 0 404892 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire18_A
timestamp 1676037725
transform -1 0 122084 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire19_A
timestamp 1676037725
transform 1 0 216384 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire20_A
timestamp 1676037725
transform 1 0 309856 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire21_A
timestamp 1676037725
transform 1 0 403236 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire22_A
timestamp 1676037725
transform -1 0 121532 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire23_A
timestamp 1676037725
transform 1 0 215188 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire24_A
timestamp 1676037725
transform 1 0 308752 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire25_A
timestamp 1676037725
transform 1 0 401488 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire26_A
timestamp 1676037725
transform -1 0 120520 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire27_A
timestamp 1676037725
transform 1 0 213624 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire28_A
timestamp 1676037725
transform 1 0 307004 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire29_A
timestamp 1676037725
transform 1 0 119232 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire30_A
timestamp 1676037725
transform -1 0 212796 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire31_A
timestamp 1676037725
transform 1 0 305348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire32_A
timestamp 1676037725
transform 1 0 117944 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire33_A
timestamp 1676037725
transform -1 0 211416 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire34_A
timestamp 1676037725
transform -1 0 117484 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire35_A
timestamp 1676037725
transform -1 0 209024 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire36_A
timestamp 1676037725
transform -1 0 115736 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire37_A
timestamp 1676037725
transform -1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire38_A
timestamp 1676037725
transform 1 0 541328 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire39_A
timestamp 1676037725
transform -1 0 447580 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire40_A
timestamp 1676037725
transform -1 0 353740 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire41_A
timestamp 1676037725
transform -1 0 259900 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire42_A
timestamp 1676037725
transform -1 0 166336 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire43_A
timestamp 1676037725
transform -1 0 72128 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire44_A
timestamp 1676037725
transform -1 0 526424 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire45_A
timestamp 1676037725
transform -1 0 432216 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire46_A
timestamp 1676037725
transform -1 0 338376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire47_A
timestamp 1676037725
transform -1 0 244444 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire48_A
timestamp 1676037725
transform -1 0 151064 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire49_A
timestamp 1676037725
transform -1 0 56672 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire50_A
timestamp 1676037725
transform -1 0 495512 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire51_A
timestamp 1676037725
transform -1 0 401304 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire52_A
timestamp 1676037725
transform -1 0 307648 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire53_A
timestamp 1676037725
transform -1 0 213532 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire54_A
timestamp 1676037725
transform -1 0 119140 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire55_A
timestamp 1676037725
transform -1 0 480056 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire56_A
timestamp 1676037725
transform -1 0 385848 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire57_A
timestamp 1676037725
transform -1 0 292284 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire58_A
timestamp 1676037725
transform -1 0 198076 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire59_A
timestamp 1676037725
transform -1 0 104788 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire60_A
timestamp 1676037725
transform -1 0 449144 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire61_A
timestamp 1676037725
transform -1 0 354936 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire62_A
timestamp 1676037725
transform -1 0 261924 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire63_A
timestamp 1676037725
transform -1 0 168360 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire64_A
timestamp 1676037725
transform -1 0 74244 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire65_A
timestamp 1676037725
transform -1 0 433688 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire66_A
timestamp 1676037725
transform -1 0 339480 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire67_A
timestamp 1676037725
transform 1 0 246100 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire68_A
timestamp 1676037725
transform -1 0 152904 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire69_A
timestamp 1676037725
transform -1 0 58972 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire70_A
timestamp 1676037725
transform -1 0 402776 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire71_A
timestamp 1676037725
transform -1 0 309488 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire72_A
timestamp 1676037725
transform -1 0 215556 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire73_A
timestamp 1676037725
transform -1 0 122636 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire74_A
timestamp 1676037725
transform -1 0 387320 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire75_A
timestamp 1676037725
transform 1 0 293664 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire76_A
timestamp 1676037725
transform -1 0 200284 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire77_A
timestamp 1676037725
transform -1 0 107180 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire78_A
timestamp 1676037725
transform -1 0 356408 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire79_A
timestamp 1676037725
transform 1 0 262936 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire80_A
timestamp 1676037725
transform -1 0 170016 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire81_A
timestamp 1676037725
transform -1 0 76268 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire82_A
timestamp 1676037725
transform -1 0 341504 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire83_A
timestamp 1676037725
transform 1 0 247572 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire84_A
timestamp 1676037725
transform -1 0 154652 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire85_A
timestamp 1676037725
transform -1 0 61088 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire86_A
timestamp 1676037725
transform -1 0 310960 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire87_A
timestamp 1676037725
transform -1 0 217304 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire88_A
timestamp 1676037725
transform -1 0 123832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire89_A
timestamp 1676037725
transform 1 0 294768 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire90_A
timestamp 1676037725
transform -1 0 201848 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire91_A
timestamp 1676037725
transform 1 0 108468 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire92_A
timestamp 1676037725
transform 1 0 264040 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire93_A
timestamp 1676037725
transform 1 0 171028 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire94_A
timestamp 1676037725
transform -1 0 78200 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire95_A
timestamp 1676037725
transform 1 0 248676 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire96_A
timestamp 1676037725
transform 1 0 155756 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire97_A
timestamp 1676037725
transform -1 0 63480 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire98_A
timestamp 1676037725
transform -1 0 218132 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire99_A
timestamp 1676037725
transform -1 0 125488 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire100_A
timestamp 1676037725
transform -1 0 32844 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire101_A
timestamp 1676037725
transform -1 0 202860 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire102_A
timestamp 1676037725
transform -1 0 110308 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire103_A
timestamp 1676037725
transform 1 0 172040 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire104_A
timestamp 1676037725
transform -1 0 79948 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire105_A
timestamp 1676037725
transform 1 0 156676 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire106_A
timestamp 1676037725
transform -1 0 64768 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire107_A
timestamp 1676037725
transform -1 0 126500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire108_A
timestamp 1676037725
transform -1 0 35236 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire109_A
timestamp 1676037725
transform -1 0 111320 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire110_A
timestamp 1676037725
transform -1 0 81420 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire111_A
timestamp 1676037725
transform -1 0 66056 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23
timestamp 1676037725
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1676037725
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1676037725
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1676037725
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1676037725
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_169 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_179
timestamp 1676037725
transform 1 0 17572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_185 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18124 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1676037725
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1676037725
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1676037725
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1676037725
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1676037725
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1676037725
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1676037725
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1676037725
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1676037725
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_347
timestamp 1676037725
transform 1 0 33028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_359
timestamp 1676037725
transform 1 0 34132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1676037725
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1676037725
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1676037725
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1676037725
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1676037725
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1676037725
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1676037725
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1676037725
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1676037725
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1676037725
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_515
timestamp 1676037725
transform 1 0 48484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_527
timestamp 1676037725
transform 1 0 49588 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_531
timestamp 1676037725
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1676037725
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_545
timestamp 1676037725
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1676037725
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_561
timestamp 1676037725
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_573
timestamp 1676037725
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1676037725
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_589
timestamp 1676037725
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_601
timestamp 1676037725
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1676037725
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_617
timestamp 1676037725
transform 1 0 57868 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_629
timestamp 1676037725
transform 1 0 58972 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_641
timestamp 1676037725
transform 1 0 60076 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_645
timestamp 1676037725
transform 1 0 60444 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_657
timestamp 1676037725
transform 1 0 61548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_669
timestamp 1676037725
transform 1 0 62652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_673
timestamp 1676037725
transform 1 0 63020 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_683
timestamp 1676037725
transform 1 0 63940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_695
timestamp 1676037725
transform 1 0 65044 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_699
timestamp 1676037725
transform 1 0 65412 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_701
timestamp 1676037725
transform 1 0 65596 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_713
timestamp 1676037725
transform 1 0 66700 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_725
timestamp 1676037725
transform 1 0 67804 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_729
timestamp 1676037725
transform 1 0 68172 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_741
timestamp 1676037725
transform 1 0 69276 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_753
timestamp 1676037725
transform 1 0 70380 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_757
timestamp 1676037725
transform 1 0 70748 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_769
timestamp 1676037725
transform 1 0 71852 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_781
timestamp 1676037725
transform 1 0 72956 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_785
timestamp 1676037725
transform 1 0 73324 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_797
timestamp 1676037725
transform 1 0 74428 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_809
timestamp 1676037725
transform 1 0 75532 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_813
timestamp 1676037725
transform 1 0 75900 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_825
timestamp 1676037725
transform 1 0 77004 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_837
timestamp 1676037725
transform 1 0 78108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_841
timestamp 1676037725
transform 1 0 78476 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_851
timestamp 1676037725
transform 1 0 79396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_863
timestamp 1676037725
transform 1 0 80500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_867
timestamp 1676037725
transform 1 0 80868 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_869
timestamp 1676037725
transform 1 0 81052 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_881
timestamp 1676037725
transform 1 0 82156 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_893
timestamp 1676037725
transform 1 0 83260 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_897
timestamp 1676037725
transform 1 0 83628 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_909
timestamp 1676037725
transform 1 0 84732 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_921
timestamp 1676037725
transform 1 0 85836 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_925
timestamp 1676037725
transform 1 0 86204 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_937
timestamp 1676037725
transform 1 0 87308 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_949
timestamp 1676037725
transform 1 0 88412 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_953
timestamp 1676037725
transform 1 0 88780 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_965
timestamp 1676037725
transform 1 0 89884 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_977
timestamp 1676037725
transform 1 0 90988 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_981
timestamp 1676037725
transform 1 0 91356 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_993
timestamp 1676037725
transform 1 0 92460 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1005
timestamp 1676037725
transform 1 0 93564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1009
timestamp 1676037725
transform 1 0 93932 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1019
timestamp 1676037725
transform 1 0 94852 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1031
timestamp 1676037725
transform 1 0 95956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1035
timestamp 1676037725
transform 1 0 96324 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1037
timestamp 1676037725
transform 1 0 96508 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1049
timestamp 1676037725
transform 1 0 97612 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1061
timestamp 1676037725
transform 1 0 98716 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1065
timestamp 1676037725
transform 1 0 99084 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1077
timestamp 1676037725
transform 1 0 100188 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1089
timestamp 1676037725
transform 1 0 101292 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1093
timestamp 1676037725
transform 1 0 101660 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1105
timestamp 1676037725
transform 1 0 102764 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1117
timestamp 1676037725
transform 1 0 103868 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1121
timestamp 1676037725
transform 1 0 104236 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1133
timestamp 1676037725
transform 1 0 105340 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1145
timestamp 1676037725
transform 1 0 106444 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1149
timestamp 1676037725
transform 1 0 106812 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1161
timestamp 1676037725
transform 1 0 107916 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1173
timestamp 1676037725
transform 1 0 109020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1177
timestamp 1676037725
transform 1 0 109388 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1187
timestamp 1676037725
transform 1 0 110308 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1199
timestamp 1676037725
transform 1 0 111412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1203
timestamp 1676037725
transform 1 0 111780 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1205
timestamp 1676037725
transform 1 0 111964 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1217
timestamp 1676037725
transform 1 0 113068 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1229
timestamp 1676037725
transform 1 0 114172 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1233
timestamp 1676037725
transform 1 0 114540 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1245
timestamp 1676037725
transform 1 0 115644 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1257
timestamp 1676037725
transform 1 0 116748 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1261
timestamp 1676037725
transform 1 0 117116 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1273
timestamp 1676037725
transform 1 0 118220 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1285
timestamp 1676037725
transform 1 0 119324 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1289
timestamp 1676037725
transform 1 0 119692 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1301
timestamp 1676037725
transform 1 0 120796 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1313
timestamp 1676037725
transform 1 0 121900 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1317
timestamp 1676037725
transform 1 0 122268 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1329
timestamp 1676037725
transform 1 0 123372 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1341
timestamp 1676037725
transform 1 0 124476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1345
timestamp 1676037725
transform 1 0 124844 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1355
timestamp 1676037725
transform 1 0 125764 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1367
timestamp 1676037725
transform 1 0 126868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1371
timestamp 1676037725
transform 1 0 127236 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1373
timestamp 1676037725
transform 1 0 127420 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1385
timestamp 1676037725
transform 1 0 128524 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1397
timestamp 1676037725
transform 1 0 129628 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1401
timestamp 1676037725
transform 1 0 129996 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1413
timestamp 1676037725
transform 1 0 131100 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1425
timestamp 1676037725
transform 1 0 132204 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1429
timestamp 1676037725
transform 1 0 132572 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1441
timestamp 1676037725
transform 1 0 133676 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1453
timestamp 1676037725
transform 1 0 134780 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1457
timestamp 1676037725
transform 1 0 135148 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1469
timestamp 1676037725
transform 1 0 136252 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1481
timestamp 1676037725
transform 1 0 137356 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1485
timestamp 1676037725
transform 1 0 137724 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1497
timestamp 1676037725
transform 1 0 138828 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1509
timestamp 1676037725
transform 1 0 139932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1513
timestamp 1676037725
transform 1 0 140300 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1523
timestamp 1676037725
transform 1 0 141220 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1535
timestamp 1676037725
transform 1 0 142324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1539
timestamp 1676037725
transform 1 0 142692 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1541
timestamp 1676037725
transform 1 0 142876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1553
timestamp 1676037725
transform 1 0 143980 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1565
timestamp 1676037725
transform 1 0 145084 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1569
timestamp 1676037725
transform 1 0 145452 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1581
timestamp 1676037725
transform 1 0 146556 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1593
timestamp 1676037725
transform 1 0 147660 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1597
timestamp 1676037725
transform 1 0 148028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1609
timestamp 1676037725
transform 1 0 149132 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1621
timestamp 1676037725
transform 1 0 150236 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1625
timestamp 1676037725
transform 1 0 150604 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1637
timestamp 1676037725
transform 1 0 151708 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1649
timestamp 1676037725
transform 1 0 152812 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1653
timestamp 1676037725
transform 1 0 153180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1665
timestamp 1676037725
transform 1 0 154284 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1677
timestamp 1676037725
transform 1 0 155388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1681
timestamp 1676037725
transform 1 0 155756 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1691
timestamp 1676037725
transform 1 0 156676 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1703
timestamp 1676037725
transform 1 0 157780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1707
timestamp 1676037725
transform 1 0 158148 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1709
timestamp 1676037725
transform 1 0 158332 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1721
timestamp 1676037725
transform 1 0 159436 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1733
timestamp 1676037725
transform 1 0 160540 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1737
timestamp 1676037725
transform 1 0 160908 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1749
timestamp 1676037725
transform 1 0 162012 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1761
timestamp 1676037725
transform 1 0 163116 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1765
timestamp 1676037725
transform 1 0 163484 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1777
timestamp 1676037725
transform 1 0 164588 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1789
timestamp 1676037725
transform 1 0 165692 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1793
timestamp 1676037725
transform 1 0 166060 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1805
timestamp 1676037725
transform 1 0 167164 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1817
timestamp 1676037725
transform 1 0 168268 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1821
timestamp 1676037725
transform 1 0 168636 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1833
timestamp 1676037725
transform 1 0 169740 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1845
timestamp 1676037725
transform 1 0 170844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1849
timestamp 1676037725
transform 1 0 171212 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1859
timestamp 1676037725
transform 1 0 172132 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1871
timestamp 1676037725
transform 1 0 173236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1875
timestamp 1676037725
transform 1 0 173604 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1877
timestamp 1676037725
transform 1 0 173788 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1889
timestamp 1676037725
transform 1 0 174892 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1901
timestamp 1676037725
transform 1 0 175996 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1905
timestamp 1676037725
transform 1 0 176364 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1917
timestamp 1676037725
transform 1 0 177468 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1929
timestamp 1676037725
transform 1 0 178572 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1933
timestamp 1676037725
transform 1 0 178940 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1945
timestamp 1676037725
transform 1 0 180044 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1957
timestamp 1676037725
transform 1 0 181148 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1961
timestamp 1676037725
transform 1 0 181516 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1973
timestamp 1676037725
transform 1 0 182620 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1985
timestamp 1676037725
transform 1 0 183724 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1989
timestamp 1676037725
transform 1 0 184092 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2001
timestamp 1676037725
transform 1 0 185196 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2013
timestamp 1676037725
transform 1 0 186300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2017
timestamp 1676037725
transform 1 0 186668 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2027
timestamp 1676037725
transform 1 0 187588 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2039
timestamp 1676037725
transform 1 0 188692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2043
timestamp 1676037725
transform 1 0 189060 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2045
timestamp 1676037725
transform 1 0 189244 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2057
timestamp 1676037725
transform 1 0 190348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2069
timestamp 1676037725
transform 1 0 191452 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2073
timestamp 1676037725
transform 1 0 191820 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2085
timestamp 1676037725
transform 1 0 192924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2097
timestamp 1676037725
transform 1 0 194028 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2101
timestamp 1676037725
transform 1 0 194396 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2113
timestamp 1676037725
transform 1 0 195500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2125
timestamp 1676037725
transform 1 0 196604 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2129
timestamp 1676037725
transform 1 0 196972 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2141
timestamp 1676037725
transform 1 0 198076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2153
timestamp 1676037725
transform 1 0 199180 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2157
timestamp 1676037725
transform 1 0 199548 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2169
timestamp 1676037725
transform 1 0 200652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2181
timestamp 1676037725
transform 1 0 201756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2185
timestamp 1676037725
transform 1 0 202124 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2195
timestamp 1676037725
transform 1 0 203044 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2207
timestamp 1676037725
transform 1 0 204148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2211
timestamp 1676037725
transform 1 0 204516 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2213
timestamp 1676037725
transform 1 0 204700 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2225
timestamp 1676037725
transform 1 0 205804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2237
timestamp 1676037725
transform 1 0 206908 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2241
timestamp 1676037725
transform 1 0 207276 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2253
timestamp 1676037725
transform 1 0 208380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2265
timestamp 1676037725
transform 1 0 209484 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2269
timestamp 1676037725
transform 1 0 209852 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2281
timestamp 1676037725
transform 1 0 210956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2293
timestamp 1676037725
transform 1 0 212060 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2297
timestamp 1676037725
transform 1 0 212428 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2309
timestamp 1676037725
transform 1 0 213532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2321
timestamp 1676037725
transform 1 0 214636 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2325
timestamp 1676037725
transform 1 0 215004 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2337
timestamp 1676037725
transform 1 0 216108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2349
timestamp 1676037725
transform 1 0 217212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2353
timestamp 1676037725
transform 1 0 217580 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2363
timestamp 1676037725
transform 1 0 218500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2375
timestamp 1676037725
transform 1 0 219604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2379
timestamp 1676037725
transform 1 0 219972 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2381
timestamp 1676037725
transform 1 0 220156 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2393
timestamp 1676037725
transform 1 0 221260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2405
timestamp 1676037725
transform 1 0 222364 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2409
timestamp 1676037725
transform 1 0 222732 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2421
timestamp 1676037725
transform 1 0 223836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2433
timestamp 1676037725
transform 1 0 224940 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2437
timestamp 1676037725
transform 1 0 225308 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2449
timestamp 1676037725
transform 1 0 226412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2461
timestamp 1676037725
transform 1 0 227516 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2465
timestamp 1676037725
transform 1 0 227884 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2477
timestamp 1676037725
transform 1 0 228988 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2489
timestamp 1676037725
transform 1 0 230092 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2493
timestamp 1676037725
transform 1 0 230460 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2505
timestamp 1676037725
transform 1 0 231564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2517
timestamp 1676037725
transform 1 0 232668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2521
timestamp 1676037725
transform 1 0 233036 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2531
timestamp 1676037725
transform 1 0 233956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2543
timestamp 1676037725
transform 1 0 235060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2547
timestamp 1676037725
transform 1 0 235428 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2549
timestamp 1676037725
transform 1 0 235612 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2561
timestamp 1676037725
transform 1 0 236716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2573
timestamp 1676037725
transform 1 0 237820 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2577
timestamp 1676037725
transform 1 0 238188 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2589
timestamp 1676037725
transform 1 0 239292 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2601
timestamp 1676037725
transform 1 0 240396 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2605
timestamp 1676037725
transform 1 0 240764 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2617
timestamp 1676037725
transform 1 0 241868 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2629
timestamp 1676037725
transform 1 0 242972 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2633
timestamp 1676037725
transform 1 0 243340 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2645
timestamp 1676037725
transform 1 0 244444 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2657
timestamp 1676037725
transform 1 0 245548 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2661
timestamp 1676037725
transform 1 0 245916 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2673
timestamp 1676037725
transform 1 0 247020 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2685
timestamp 1676037725
transform 1 0 248124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2689
timestamp 1676037725
transform 1 0 248492 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2699
timestamp 1676037725
transform 1 0 249412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2711
timestamp 1676037725
transform 1 0 250516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2715
timestamp 1676037725
transform 1 0 250884 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2717
timestamp 1676037725
transform 1 0 251068 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2729
timestamp 1676037725
transform 1 0 252172 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2741
timestamp 1676037725
transform 1 0 253276 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2745
timestamp 1676037725
transform 1 0 253644 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2757
timestamp 1676037725
transform 1 0 254748 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2769
timestamp 1676037725
transform 1 0 255852 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2773
timestamp 1676037725
transform 1 0 256220 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2785
timestamp 1676037725
transform 1 0 257324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2797
timestamp 1676037725
transform 1 0 258428 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2801
timestamp 1676037725
transform 1 0 258796 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2813
timestamp 1676037725
transform 1 0 259900 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2825
timestamp 1676037725
transform 1 0 261004 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2829
timestamp 1676037725
transform 1 0 261372 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2841
timestamp 1676037725
transform 1 0 262476 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2853
timestamp 1676037725
transform 1 0 263580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2857
timestamp 1676037725
transform 1 0 263948 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2867
timestamp 1676037725
transform 1 0 264868 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2879
timestamp 1676037725
transform 1 0 265972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2883
timestamp 1676037725
transform 1 0 266340 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2885
timestamp 1676037725
transform 1 0 266524 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2897
timestamp 1676037725
transform 1 0 267628 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2909
timestamp 1676037725
transform 1 0 268732 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2913
timestamp 1676037725
transform 1 0 269100 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2925
timestamp 1676037725
transform 1 0 270204 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2937
timestamp 1676037725
transform 1 0 271308 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2941
timestamp 1676037725
transform 1 0 271676 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2953
timestamp 1676037725
transform 1 0 272780 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2965
timestamp 1676037725
transform 1 0 273884 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2969
timestamp 1676037725
transform 1 0 274252 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2981
timestamp 1676037725
transform 1 0 275356 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2993
timestamp 1676037725
transform 1 0 276460 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2997
timestamp 1676037725
transform 1 0 276828 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3009
timestamp 1676037725
transform 1 0 277932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3021
timestamp 1676037725
transform 1 0 279036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3025
timestamp 1676037725
transform 1 0 279404 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3035
timestamp 1676037725
transform 1 0 280324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3047
timestamp 1676037725
transform 1 0 281428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3051
timestamp 1676037725
transform 1 0 281796 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3053
timestamp 1676037725
transform 1 0 281980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3065
timestamp 1676037725
transform 1 0 283084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3077
timestamp 1676037725
transform 1 0 284188 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3081
timestamp 1676037725
transform 1 0 284556 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3093
timestamp 1676037725
transform 1 0 285660 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3105
timestamp 1676037725
transform 1 0 286764 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3109
timestamp 1676037725
transform 1 0 287132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3121
timestamp 1676037725
transform 1 0 288236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3133
timestamp 1676037725
transform 1 0 289340 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3137
timestamp 1676037725
transform 1 0 289708 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3149
timestamp 1676037725
transform 1 0 290812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3161
timestamp 1676037725
transform 1 0 291916 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3165
timestamp 1676037725
transform 1 0 292284 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3177
timestamp 1676037725
transform 1 0 293388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3189
timestamp 1676037725
transform 1 0 294492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3193
timestamp 1676037725
transform 1 0 294860 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3203
timestamp 1676037725
transform 1 0 295780 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3215
timestamp 1676037725
transform 1 0 296884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3219
timestamp 1676037725
transform 1 0 297252 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3221
timestamp 1676037725
transform 1 0 297436 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3233
timestamp 1676037725
transform 1 0 298540 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3245
timestamp 1676037725
transform 1 0 299644 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3249
timestamp 1676037725
transform 1 0 300012 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3261
timestamp 1676037725
transform 1 0 301116 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3273
timestamp 1676037725
transform 1 0 302220 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3277
timestamp 1676037725
transform 1 0 302588 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3289
timestamp 1676037725
transform 1 0 303692 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3301
timestamp 1676037725
transform 1 0 304796 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3305
timestamp 1676037725
transform 1 0 305164 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3317
timestamp 1676037725
transform 1 0 306268 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3329
timestamp 1676037725
transform 1 0 307372 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3333
timestamp 1676037725
transform 1 0 307740 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3345
timestamp 1676037725
transform 1 0 308844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3357
timestamp 1676037725
transform 1 0 309948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3361
timestamp 1676037725
transform 1 0 310316 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3371
timestamp 1676037725
transform 1 0 311236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3383
timestamp 1676037725
transform 1 0 312340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3387
timestamp 1676037725
transform 1 0 312708 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3389
timestamp 1676037725
transform 1 0 312892 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3401
timestamp 1676037725
transform 1 0 313996 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3413
timestamp 1676037725
transform 1 0 315100 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3417
timestamp 1676037725
transform 1 0 315468 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3429
timestamp 1676037725
transform 1 0 316572 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3441
timestamp 1676037725
transform 1 0 317676 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3445
timestamp 1676037725
transform 1 0 318044 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3457
timestamp 1676037725
transform 1 0 319148 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3469
timestamp 1676037725
transform 1 0 320252 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3473
timestamp 1676037725
transform 1 0 320620 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3485
timestamp 1676037725
transform 1 0 321724 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3497
timestamp 1676037725
transform 1 0 322828 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3501
timestamp 1676037725
transform 1 0 323196 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3513
timestamp 1676037725
transform 1 0 324300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3525
timestamp 1676037725
transform 1 0 325404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3529
timestamp 1676037725
transform 1 0 325772 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3539
timestamp 1676037725
transform 1 0 326692 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3551
timestamp 1676037725
transform 1 0 327796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3555
timestamp 1676037725
transform 1 0 328164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3557
timestamp 1676037725
transform 1 0 328348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3569
timestamp 1676037725
transform 1 0 329452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3581
timestamp 1676037725
transform 1 0 330556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3585
timestamp 1676037725
transform 1 0 330924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3597
timestamp 1676037725
transform 1 0 332028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3609
timestamp 1676037725
transform 1 0 333132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3613
timestamp 1676037725
transform 1 0 333500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3625
timestamp 1676037725
transform 1 0 334604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3637
timestamp 1676037725
transform 1 0 335708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3641
timestamp 1676037725
transform 1 0 336076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3653
timestamp 1676037725
transform 1 0 337180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3665
timestamp 1676037725
transform 1 0 338284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3669
timestamp 1676037725
transform 1 0 338652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3681
timestamp 1676037725
transform 1 0 339756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3693
timestamp 1676037725
transform 1 0 340860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3697
timestamp 1676037725
transform 1 0 341228 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3707
timestamp 1676037725
transform 1 0 342148 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3719
timestamp 1676037725
transform 1 0 343252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3723
timestamp 1676037725
transform 1 0 343620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3725
timestamp 1676037725
transform 1 0 343804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3737
timestamp 1676037725
transform 1 0 344908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3749
timestamp 1676037725
transform 1 0 346012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3753
timestamp 1676037725
transform 1 0 346380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3765
timestamp 1676037725
transform 1 0 347484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3777
timestamp 1676037725
transform 1 0 348588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3781
timestamp 1676037725
transform 1 0 348956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3793
timestamp 1676037725
transform 1 0 350060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3805
timestamp 1676037725
transform 1 0 351164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3809
timestamp 1676037725
transform 1 0 351532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3821
timestamp 1676037725
transform 1 0 352636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3833
timestamp 1676037725
transform 1 0 353740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3837
timestamp 1676037725
transform 1 0 354108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3849
timestamp 1676037725
transform 1 0 355212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3861
timestamp 1676037725
transform 1 0 356316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3865
timestamp 1676037725
transform 1 0 356684 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3875
timestamp 1676037725
transform 1 0 357604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3887
timestamp 1676037725
transform 1 0 358708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3891
timestamp 1676037725
transform 1 0 359076 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3893
timestamp 1676037725
transform 1 0 359260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3905
timestamp 1676037725
transform 1 0 360364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3917
timestamp 1676037725
transform 1 0 361468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3921
timestamp 1676037725
transform 1 0 361836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3933
timestamp 1676037725
transform 1 0 362940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3945
timestamp 1676037725
transform 1 0 364044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3949
timestamp 1676037725
transform 1 0 364412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3961
timestamp 1676037725
transform 1 0 365516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3973
timestamp 1676037725
transform 1 0 366620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3977
timestamp 1676037725
transform 1 0 366988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3989
timestamp 1676037725
transform 1 0 368092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4001
timestamp 1676037725
transform 1 0 369196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4005
timestamp 1676037725
transform 1 0 369564 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4017
timestamp 1676037725
transform 1 0 370668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4029
timestamp 1676037725
transform 1 0 371772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4033
timestamp 1676037725
transform 1 0 372140 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4043
timestamp 1676037725
transform 1 0 373060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4055
timestamp 1676037725
transform 1 0 374164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4059
timestamp 1676037725
transform 1 0 374532 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4061
timestamp 1676037725
transform 1 0 374716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4073
timestamp 1676037725
transform 1 0 375820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4085
timestamp 1676037725
transform 1 0 376924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4089
timestamp 1676037725
transform 1 0 377292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4101
timestamp 1676037725
transform 1 0 378396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4113
timestamp 1676037725
transform 1 0 379500 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4117
timestamp 1676037725
transform 1 0 379868 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4129
timestamp 1676037725
transform 1 0 380972 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4141
timestamp 1676037725
transform 1 0 382076 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4145
timestamp 1676037725
transform 1 0 382444 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4157
timestamp 1676037725
transform 1 0 383548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4169
timestamp 1676037725
transform 1 0 384652 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4173
timestamp 1676037725
transform 1 0 385020 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4185
timestamp 1676037725
transform 1 0 386124 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4197
timestamp 1676037725
transform 1 0 387228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4201
timestamp 1676037725
transform 1 0 387596 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4211
timestamp 1676037725
transform 1 0 388516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4223
timestamp 1676037725
transform 1 0 389620 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4227
timestamp 1676037725
transform 1 0 389988 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4229
timestamp 1676037725
transform 1 0 390172 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4241
timestamp 1676037725
transform 1 0 391276 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4253
timestamp 1676037725
transform 1 0 392380 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4257
timestamp 1676037725
transform 1 0 392748 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4269
timestamp 1676037725
transform 1 0 393852 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4281
timestamp 1676037725
transform 1 0 394956 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4285
timestamp 1676037725
transform 1 0 395324 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4297
timestamp 1676037725
transform 1 0 396428 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4309
timestamp 1676037725
transform 1 0 397532 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4313
timestamp 1676037725
transform 1 0 397900 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4325
timestamp 1676037725
transform 1 0 399004 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4337
timestamp 1676037725
transform 1 0 400108 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4341
timestamp 1676037725
transform 1 0 400476 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4353
timestamp 1676037725
transform 1 0 401580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4361
timestamp 1676037725
transform 1 0 402316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4366 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 402776 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4369
timestamp 1676037725
transform 1 0 403052 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4379
timestamp 1676037725
transform 1 0 403972 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4391
timestamp 1676037725
transform 1 0 405076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4395
timestamp 1676037725
transform 1 0 405444 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4397
timestamp 1676037725
transform 1 0 405628 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4409
timestamp 1676037725
transform 1 0 406732 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4421
timestamp 1676037725
transform 1 0 407836 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4425
timestamp 1676037725
transform 1 0 408204 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4437
timestamp 1676037725
transform 1 0 409308 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4449
timestamp 1676037725
transform 1 0 410412 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4453
timestamp 1676037725
transform 1 0 410780 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4465
timestamp 1676037725
transform 1 0 411884 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4477
timestamp 1676037725
transform 1 0 412988 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4481
timestamp 1676037725
transform 1 0 413356 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4493
timestamp 1676037725
transform 1 0 414460 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4505
timestamp 1676037725
transform 1 0 415564 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4509
timestamp 1676037725
transform 1 0 415932 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4521
timestamp 1676037725
transform 1 0 417036 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4533
timestamp 1676037725
transform 1 0 418140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4537
timestamp 1676037725
transform 1 0 418508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4543
timestamp 1676037725
transform 1 0 419060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4547
timestamp 1676037725
transform 1 0 419428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4553
timestamp 1676037725
transform 1 0 419980 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4561
timestamp 1676037725
transform 1 0 420716 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4565
timestamp 1676037725
transform 1 0 421084 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4577
timestamp 1676037725
transform 1 0 422188 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4589
timestamp 1676037725
transform 1 0 423292 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4593
timestamp 1676037725
transform 1 0 423660 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4605
timestamp 1676037725
transform 1 0 424764 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4617
timestamp 1676037725
transform 1 0 425868 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4621
timestamp 1676037725
transform 1 0 426236 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4633
timestamp 1676037725
transform 1 0 427340 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4645
timestamp 1676037725
transform 1 0 428444 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4649
timestamp 1676037725
transform 1 0 428812 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4661
timestamp 1676037725
transform 1 0 429916 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4673
timestamp 1676037725
transform 1 0 431020 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4677
timestamp 1676037725
transform 1 0 431388 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4689
timestamp 1676037725
transform 1 0 432492 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4701
timestamp 1676037725
transform 1 0 433596 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4705
timestamp 1676037725
transform 1 0 433964 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4715
timestamp 1676037725
transform 1 0 434884 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4727
timestamp 1676037725
transform 1 0 435988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4731
timestamp 1676037725
transform 1 0 436356 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4733
timestamp 1676037725
transform 1 0 436540 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4745
timestamp 1676037725
transform 1 0 437644 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4757
timestamp 1676037725
transform 1 0 438748 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4761
timestamp 1676037725
transform 1 0 439116 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4773
timestamp 1676037725
transform 1 0 440220 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4785
timestamp 1676037725
transform 1 0 441324 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4789
timestamp 1676037725
transform 1 0 441692 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4801
timestamp 1676037725
transform 1 0 442796 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4813
timestamp 1676037725
transform 1 0 443900 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4817
timestamp 1676037725
transform 1 0 444268 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4829
timestamp 1676037725
transform 1 0 445372 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4841
timestamp 1676037725
transform 1 0 446476 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4845
timestamp 1676037725
transform 1 0 446844 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4857
timestamp 1676037725
transform 1 0 447948 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4869
timestamp 1676037725
transform 1 0 449052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4873
timestamp 1676037725
transform 1 0 449420 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4883
timestamp 1676037725
transform 1 0 450340 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4895
timestamp 1676037725
transform 1 0 451444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4899
timestamp 1676037725
transform 1 0 451812 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4901
timestamp 1676037725
transform 1 0 451996 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4913
timestamp 1676037725
transform 1 0 453100 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4925
timestamp 1676037725
transform 1 0 454204 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4929
timestamp 1676037725
transform 1 0 454572 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4941
timestamp 1676037725
transform 1 0 455676 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4953
timestamp 1676037725
transform 1 0 456780 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4957
timestamp 1676037725
transform 1 0 457148 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4969
timestamp 1676037725
transform 1 0 458252 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4981
timestamp 1676037725
transform 1 0 459356 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4985
timestamp 1676037725
transform 1 0 459724 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4997
timestamp 1676037725
transform 1 0 460828 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5009
timestamp 1676037725
transform 1 0 461932 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5013
timestamp 1676037725
transform 1 0 462300 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5025
timestamp 1676037725
transform 1 0 463404 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5037
timestamp 1676037725
transform 1 0 464508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5041
timestamp 1676037725
transform 1 0 464876 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5051
timestamp 1676037725
transform 1 0 465796 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5063
timestamp 1676037725
transform 1 0 466900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5067
timestamp 1676037725
transform 1 0 467268 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5069
timestamp 1676037725
transform 1 0 467452 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5081
timestamp 1676037725
transform 1 0 468556 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5093
timestamp 1676037725
transform 1 0 469660 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5097
timestamp 1676037725
transform 1 0 470028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5109
timestamp 1676037725
transform 1 0 471132 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5121
timestamp 1676037725
transform 1 0 472236 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5125
timestamp 1676037725
transform 1 0 472604 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5137
timestamp 1676037725
transform 1 0 473708 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5149
timestamp 1676037725
transform 1 0 474812 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5153
timestamp 1676037725
transform 1 0 475180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5165
timestamp 1676037725
transform 1 0 476284 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5177
timestamp 1676037725
transform 1 0 477388 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5181
timestamp 1676037725
transform 1 0 477756 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5193
timestamp 1676037725
transform 1 0 478860 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5205
timestamp 1676037725
transform 1 0 479964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5209
timestamp 1676037725
transform 1 0 480332 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5219
timestamp 1676037725
transform 1 0 481252 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5231
timestamp 1676037725
transform 1 0 482356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5235
timestamp 1676037725
transform 1 0 482724 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5237
timestamp 1676037725
transform 1 0 482908 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5249
timestamp 1676037725
transform 1 0 484012 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5261
timestamp 1676037725
transform 1 0 485116 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5265
timestamp 1676037725
transform 1 0 485484 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5277
timestamp 1676037725
transform 1 0 486588 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5289
timestamp 1676037725
transform 1 0 487692 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5293
timestamp 1676037725
transform 1 0 488060 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5305
timestamp 1676037725
transform 1 0 489164 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5317
timestamp 1676037725
transform 1 0 490268 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5321
timestamp 1676037725
transform 1 0 490636 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5333
timestamp 1676037725
transform 1 0 491740 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5345
timestamp 1676037725
transform 1 0 492844 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5349
timestamp 1676037725
transform 1 0 493212 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5361
timestamp 1676037725
transform 1 0 494316 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5373
timestamp 1676037725
transform 1 0 495420 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5377
timestamp 1676037725
transform 1 0 495788 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5387
timestamp 1676037725
transform 1 0 496708 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5399
timestamp 1676037725
transform 1 0 497812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5403
timestamp 1676037725
transform 1 0 498180 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5405
timestamp 1676037725
transform 1 0 498364 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5417
timestamp 1676037725
transform 1 0 499468 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5429
timestamp 1676037725
transform 1 0 500572 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5433
timestamp 1676037725
transform 1 0 500940 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5445
timestamp 1676037725
transform 1 0 502044 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5457
timestamp 1676037725
transform 1 0 503148 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5461
timestamp 1676037725
transform 1 0 503516 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5473
timestamp 1676037725
transform 1 0 504620 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5485
timestamp 1676037725
transform 1 0 505724 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5489
timestamp 1676037725
transform 1 0 506092 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5501
timestamp 1676037725
transform 1 0 507196 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5513
timestamp 1676037725
transform 1 0 508300 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5517
timestamp 1676037725
transform 1 0 508668 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5529
timestamp 1676037725
transform 1 0 509772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5541
timestamp 1676037725
transform 1 0 510876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5545
timestamp 1676037725
transform 1 0 511244 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5551
timestamp 1676037725
transform 1 0 511796 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5555
timestamp 1676037725
transform 1 0 512164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5561
timestamp 1676037725
transform 1 0 512716 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5569
timestamp 1676037725
transform 1 0 513452 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5573
timestamp 1676037725
transform 1 0 513820 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5585
timestamp 1676037725
transform 1 0 514924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5597
timestamp 1676037725
transform 1 0 516028 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5601
timestamp 1676037725
transform 1 0 516396 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5613
timestamp 1676037725
transform 1 0 517500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5625
timestamp 1676037725
transform 1 0 518604 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5629
timestamp 1676037725
transform 1 0 518972 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5641
timestamp 1676037725
transform 1 0 520076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5653
timestamp 1676037725
transform 1 0 521180 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5657
timestamp 1676037725
transform 1 0 521548 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5669
timestamp 1676037725
transform 1 0 522652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5681
timestamp 1676037725
transform 1 0 523756 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5685
timestamp 1676037725
transform 1 0 524124 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5697
timestamp 1676037725
transform 1 0 525228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5709
timestamp 1676037725
transform 1 0 526332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5713
timestamp 1676037725
transform 1 0 526700 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5723
timestamp 1676037725
transform 1 0 527620 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5735
timestamp 1676037725
transform 1 0 528724 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5739
timestamp 1676037725
transform 1 0 529092 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5741
timestamp 1676037725
transform 1 0 529276 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5753
timestamp 1676037725
transform 1 0 530380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5765
timestamp 1676037725
transform 1 0 531484 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5769
timestamp 1676037725
transform 1 0 531852 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5781
timestamp 1676037725
transform 1 0 532956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5793
timestamp 1676037725
transform 1 0 534060 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5797
timestamp 1676037725
transform 1 0 534428 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5809
timestamp 1676037725
transform 1 0 535532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5821
timestamp 1676037725
transform 1 0 536636 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5825
timestamp 1676037725
transform 1 0 537004 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5837
timestamp 1676037725
transform 1 0 538108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5849
timestamp 1676037725
transform 1 0 539212 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5853
timestamp 1676037725
transform 1 0 539580 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5865
timestamp 1676037725
transform 1 0 540684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5877
timestamp 1676037725
transform 1 0 541788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5881
timestamp 1676037725
transform 1 0 542156 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5891
timestamp 1676037725
transform 1 0 543076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5903
timestamp 1676037725
transform 1 0 544180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5907
timestamp 1676037725
transform 1 0 544548 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5909
timestamp 1676037725
transform 1 0 544732 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5921
timestamp 1676037725
transform 1 0 545836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5933
timestamp 1676037725
transform 1 0 546940 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5937
timestamp 1676037725
transform 1 0 547308 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5949
timestamp 1676037725
transform 1 0 548412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5961
timestamp 1676037725
transform 1 0 549516 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5965
timestamp 1676037725
transform 1 0 549884 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5977
timestamp 1676037725
transform 1 0 550988 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5989
timestamp 1676037725
transform 1 0 552092 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5993
timestamp 1676037725
transform 1 0 552460 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6005
timestamp 1676037725
transform 1 0 553564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6017
timestamp 1676037725
transform 1 0 554668 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6021
timestamp 1676037725
transform 1 0 555036 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6033
timestamp 1676037725
transform 1 0 556140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6045
timestamp 1676037725
transform 1 0 557244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6049
timestamp 1676037725
transform 1 0 557612 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6059
timestamp 1676037725
transform 1 0 558532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6071
timestamp 1676037725
transform 1 0 559636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6075
timestamp 1676037725
transform 1 0 560004 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6077
timestamp 1676037725
transform 1 0 560188 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6089
timestamp 1676037725
transform 1 0 561292 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6101
timestamp 1676037725
transform 1 0 562396 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6105
timestamp 1676037725
transform 1 0 562764 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6117
timestamp 1676037725
transform 1 0 563868 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6129
timestamp 1676037725
transform 1 0 564972 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6133
timestamp 1676037725
transform 1 0 565340 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6145
timestamp 1676037725
transform 1 0 566444 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6157
timestamp 1676037725
transform 1 0 567548 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6161
timestamp 1676037725
transform 1 0 567916 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6173
timestamp 1676037725
transform 1 0 569020 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6185
timestamp 1676037725
transform 1 0 570124 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6189
timestamp 1676037725
transform 1 0 570492 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6201
timestamp 1676037725
transform 1 0 571596 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6213
timestamp 1676037725
transform 1 0 572700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6217
timestamp 1676037725
transform 1 0 573068 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6227
timestamp 1676037725
transform 1 0 573988 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6239
timestamp 1676037725
transform 1 0 575092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6243
timestamp 1676037725
transform 1 0 575460 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6245
timestamp 1676037725
transform 1 0 575644 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6257
timestamp 1676037725
transform 1 0 576748 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6269
timestamp 1676037725
transform 1 0 577852 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6273
timestamp 1676037725
transform 1 0 578220 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6285
timestamp 1676037725
transform 1 0 579324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6297
timestamp 1676037725
transform 1 0 580428 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6301
timestamp 1676037725
transform 1 0 580796 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6313
timestamp 1676037725
transform 1 0 581900 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6325
timestamp 1676037725
transform 1 0 583004 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6329
timestamp 1676037725
transform 1 0 583372 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6341
timestamp 1676037725
transform 1 0 584476 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6353
timestamp 1676037725
transform 1 0 585580 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6357
timestamp 1676037725
transform 1 0 585948 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6369
timestamp 1676037725
transform 1 0 587052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6381
timestamp 1676037725
transform 1 0 588156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6385
timestamp 1676037725
transform 1 0 588524 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6395
timestamp 1676037725
transform 1 0 589444 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6407
timestamp 1676037725
transform 1 0 590548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6411
timestamp 1676037725
transform 1 0 590916 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6413
timestamp 1676037725
transform 1 0 591100 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6425
timestamp 1676037725
transform 1 0 592204 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6437
timestamp 1676037725
transform 1 0 593308 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6441
timestamp 1676037725
transform 1 0 593676 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6453
timestamp 1676037725
transform 1 0 594780 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6465
timestamp 1676037725
transform 1 0 595884 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6469
timestamp 1676037725
transform 1 0 596252 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6481
timestamp 1676037725
transform 1 0 597356 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6493
timestamp 1676037725
transform 1 0 598460 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6497
timestamp 1676037725
transform 1 0 598828 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6509
timestamp 1676037725
transform 1 0 599932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6521
timestamp 1676037725
transform 1 0 601036 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6525
timestamp 1676037725
transform 1 0 601404 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6537
timestamp 1676037725
transform 1 0 602508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6549
timestamp 1676037725
transform 1 0 603612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6553
timestamp 1676037725
transform 1 0 603980 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6559
timestamp 1676037725
transform 1 0 604532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6563
timestamp 1676037725
transform 1 0 604900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6569
timestamp 1676037725
transform 1 0 605452 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6577
timestamp 1676037725
transform 1 0 606188 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6581
timestamp 1676037725
transform 1 0 606556 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6593
timestamp 1676037725
transform 1 0 607660 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6605
timestamp 1676037725
transform 1 0 608764 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6609
timestamp 1676037725
transform 1 0 609132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6621
timestamp 1676037725
transform 1 0 610236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6633
timestamp 1676037725
transform 1 0 611340 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6637
timestamp 1676037725
transform 1 0 611708 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6649
timestamp 1676037725
transform 1 0 612812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6661
timestamp 1676037725
transform 1 0 613916 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6665
timestamp 1676037725
transform 1 0 614284 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6677
timestamp 1676037725
transform 1 0 615388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6689
timestamp 1676037725
transform 1 0 616492 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6693
timestamp 1676037725
transform 1 0 616860 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6705
timestamp 1676037725
transform 1 0 617964 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6717
timestamp 1676037725
transform 1 0 619068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6721
timestamp 1676037725
transform 1 0 619436 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6731
timestamp 1676037725
transform 1 0 620356 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6743
timestamp 1676037725
transform 1 0 621460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6747
timestamp 1676037725
transform 1 0 621828 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6749
timestamp 1676037725
transform 1 0 622012 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6761
timestamp 1676037725
transform 1 0 623116 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6773
timestamp 1676037725
transform 1 0 624220 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6777
timestamp 1676037725
transform 1 0 624588 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6789
timestamp 1676037725
transform 1 0 625692 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6801
timestamp 1676037725
transform 1 0 626796 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6805
timestamp 1676037725
transform 1 0 627164 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6817
timestamp 1676037725
transform 1 0 628268 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6829
timestamp 1676037725
transform 1 0 629372 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6833
timestamp 1676037725
transform 1 0 629740 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6845
timestamp 1676037725
transform 1 0 630844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6857
timestamp 1676037725
transform 1 0 631948 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6861
timestamp 1676037725
transform 1 0 632316 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6873
timestamp 1676037725
transform 1 0 633420 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6885
timestamp 1676037725
transform 1 0 634524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6889
timestamp 1676037725
transform 1 0 634892 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6899
timestamp 1676037725
transform 1 0 635812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6911
timestamp 1676037725
transform 1 0 636916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6915
timestamp 1676037725
transform 1 0 637284 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6917
timestamp 1676037725
transform 1 0 637468 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6929
timestamp 1676037725
transform 1 0 638572 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6941
timestamp 1676037725
transform 1 0 639676 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6945
timestamp 1676037725
transform 1 0 640044 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6957
timestamp 1676037725
transform 1 0 641148 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6969
timestamp 1676037725
transform 1 0 642252 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6973
timestamp 1676037725
transform 1 0 642620 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6985
timestamp 1676037725
transform 1 0 643724 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6997
timestamp 1676037725
transform 1 0 644828 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7001
timestamp 1676037725
transform 1 0 645196 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7013
timestamp 1676037725
transform 1 0 646300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7025
timestamp 1676037725
transform 1 0 647404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7029
timestamp 1676037725
transform 1 0 647772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7037
timestamp 1676037725
transform 1 0 648508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7
timestamp 1676037725
transform 1 0 1748 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_19
timestamp 1676037725
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_31
timestamp 1676037725
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_43
timestamp 1676037725
transform 1 0 5060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1676037725
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1676037725
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1676037725
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1676037725
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_343
timestamp 1676037725
transform 1 0 32660 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_355
timestamp 1676037725
transform 1 0 33764 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_367
timestamp 1676037725
transform 1 0 34868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_379
timestamp 1676037725
transform 1 0 35972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1676037725
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1676037725
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1676037725
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1676037725
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1676037725
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1676037725
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1676037725
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1676037725
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_511
timestamp 1676037725
transform 1 0 48116 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_523
timestamp 1676037725
transform 1 0 49220 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_535
timestamp 1676037725
transform 1 0 50324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_547
timestamp 1676037725
transform 1 0 51428 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1676037725
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1676037725
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1676037725
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1676037725
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1676037725
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1676037725
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1676037725
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_617
timestamp 1676037725
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_629
timestamp 1676037725
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_641
timestamp 1676037725
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_653
timestamp 1676037725
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 1676037725
transform 1 0 62284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1676037725
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_673
timestamp 1676037725
transform 1 0 63020 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_679
timestamp 1676037725
transform 1 0 63572 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_691
timestamp 1676037725
transform 1 0 64676 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_703
timestamp 1676037725
transform 1 0 65780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_715
timestamp 1676037725
transform 1 0 66884 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1676037725
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_729
timestamp 1676037725
transform 1 0 68172 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_741
timestamp 1676037725
transform 1 0 69276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_753
timestamp 1676037725
transform 1 0 70380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_765
timestamp 1676037725
transform 1 0 71484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_777
timestamp 1676037725
transform 1 0 72588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 1676037725
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_785
timestamp 1676037725
transform 1 0 73324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_797
timestamp 1676037725
transform 1 0 74428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_809
timestamp 1676037725
transform 1 0 75532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_821
timestamp 1676037725
transform 1 0 76636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_833
timestamp 1676037725
transform 1 0 77740 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_839
timestamp 1676037725
transform 1 0 78292 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_841
timestamp 1676037725
transform 1 0 78476 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_847
timestamp 1676037725
transform 1 0 79028 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_859
timestamp 1676037725
transform 1 0 80132 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_871
timestamp 1676037725
transform 1 0 81236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_883
timestamp 1676037725
transform 1 0 82340 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_895
timestamp 1676037725
transform 1 0 83444 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_897
timestamp 1676037725
transform 1 0 83628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_909
timestamp 1676037725
transform 1 0 84732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_921
timestamp 1676037725
transform 1 0 85836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_933
timestamp 1676037725
transform 1 0 86940 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_945
timestamp 1676037725
transform 1 0 88044 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_951
timestamp 1676037725
transform 1 0 88596 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_953
timestamp 1676037725
transform 1 0 88780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_965
timestamp 1676037725
transform 1 0 89884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_977
timestamp 1676037725
transform 1 0 90988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_989
timestamp 1676037725
transform 1 0 92092 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1001
timestamp 1676037725
transform 1 0 93196 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1007
timestamp 1676037725
transform 1 0 93748 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1009
timestamp 1676037725
transform 1 0 93932 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1015
timestamp 1676037725
transform 1 0 94484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1027
timestamp 1676037725
transform 1 0 95588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1039
timestamp 1676037725
transform 1 0 96692 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1051
timestamp 1676037725
transform 1 0 97796 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1063
timestamp 1676037725
transform 1 0 98900 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1065
timestamp 1676037725
transform 1 0 99084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1077
timestamp 1676037725
transform 1 0 100188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1089
timestamp 1676037725
transform 1 0 101292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1101
timestamp 1676037725
transform 1 0 102396 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1113
timestamp 1676037725
transform 1 0 103500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1119
timestamp 1676037725
transform 1 0 104052 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1121
timestamp 1676037725
transform 1 0 104236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1133
timestamp 1676037725
transform 1 0 105340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1145
timestamp 1676037725
transform 1 0 106444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1157
timestamp 1676037725
transform 1 0 107548 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1169
timestamp 1676037725
transform 1 0 108652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1175
timestamp 1676037725
transform 1 0 109204 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1177
timestamp 1676037725
transform 1 0 109388 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1183
timestamp 1676037725
transform 1 0 109940 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1195
timestamp 1676037725
transform 1 0 111044 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1207
timestamp 1676037725
transform 1 0 112148 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1219
timestamp 1676037725
transform 1 0 113252 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1231
timestamp 1676037725
transform 1 0 114356 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1233
timestamp 1676037725
transform 1 0 114540 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1245
timestamp 1676037725
transform 1 0 115644 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1257
timestamp 1676037725
transform 1 0 116748 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1269
timestamp 1676037725
transform 1 0 117852 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1281
timestamp 1676037725
transform 1 0 118956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1287
timestamp 1676037725
transform 1 0 119508 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1289
timestamp 1676037725
transform 1 0 119692 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1301
timestamp 1676037725
transform 1 0 120796 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1313
timestamp 1676037725
transform 1 0 121900 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1325
timestamp 1676037725
transform 1 0 123004 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1337
timestamp 1676037725
transform 1 0 124108 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1343
timestamp 1676037725
transform 1 0 124660 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1345
timestamp 1676037725
transform 1 0 124844 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1351
timestamp 1676037725
transform 1 0 125396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1363
timestamp 1676037725
transform 1 0 126500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1375
timestamp 1676037725
transform 1 0 127604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1387
timestamp 1676037725
transform 1 0 128708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1399
timestamp 1676037725
transform 1 0 129812 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1401
timestamp 1676037725
transform 1 0 129996 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1413
timestamp 1676037725
transform 1 0 131100 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1425
timestamp 1676037725
transform 1 0 132204 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1437
timestamp 1676037725
transform 1 0 133308 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1449
timestamp 1676037725
transform 1 0 134412 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1455
timestamp 1676037725
transform 1 0 134964 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1457
timestamp 1676037725
transform 1 0 135148 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1469
timestamp 1676037725
transform 1 0 136252 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1481
timestamp 1676037725
transform 1 0 137356 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1493
timestamp 1676037725
transform 1 0 138460 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1505
timestamp 1676037725
transform 1 0 139564 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1511
timestamp 1676037725
transform 1 0 140116 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1513
timestamp 1676037725
transform 1 0 140300 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1519
timestamp 1676037725
transform 1 0 140852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1531
timestamp 1676037725
transform 1 0 141956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1543
timestamp 1676037725
transform 1 0 143060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1555
timestamp 1676037725
transform 1 0 144164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1567
timestamp 1676037725
transform 1 0 145268 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1569
timestamp 1676037725
transform 1 0 145452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1581
timestamp 1676037725
transform 1 0 146556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1593
timestamp 1676037725
transform 1 0 147660 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1605
timestamp 1676037725
transform 1 0 148764 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1617
timestamp 1676037725
transform 1 0 149868 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1623
timestamp 1676037725
transform 1 0 150420 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1625
timestamp 1676037725
transform 1 0 150604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1637
timestamp 1676037725
transform 1 0 151708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1649
timestamp 1676037725
transform 1 0 152812 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1661
timestamp 1676037725
transform 1 0 153916 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1673
timestamp 1676037725
transform 1 0 155020 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1679
timestamp 1676037725
transform 1 0 155572 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1681
timestamp 1676037725
transform 1 0 155756 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1687
timestamp 1676037725
transform 1 0 156308 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1699
timestamp 1676037725
transform 1 0 157412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1711
timestamp 1676037725
transform 1 0 158516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1723
timestamp 1676037725
transform 1 0 159620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1735
timestamp 1676037725
transform 1 0 160724 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1737
timestamp 1676037725
transform 1 0 160908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1749
timestamp 1676037725
transform 1 0 162012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1761
timestamp 1676037725
transform 1 0 163116 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1773
timestamp 1676037725
transform 1 0 164220 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1785
timestamp 1676037725
transform 1 0 165324 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1791
timestamp 1676037725
transform 1 0 165876 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1793
timestamp 1676037725
transform 1 0 166060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1805
timestamp 1676037725
transform 1 0 167164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1817
timestamp 1676037725
transform 1 0 168268 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1829
timestamp 1676037725
transform 1 0 169372 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1841
timestamp 1676037725
transform 1 0 170476 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1847
timestamp 1676037725
transform 1 0 171028 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1849
timestamp 1676037725
transform 1 0 171212 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1855
timestamp 1676037725
transform 1 0 171764 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1867
timestamp 1676037725
transform 1 0 172868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1879
timestamp 1676037725
transform 1 0 173972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1891
timestamp 1676037725
transform 1 0 175076 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1903
timestamp 1676037725
transform 1 0 176180 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1905
timestamp 1676037725
transform 1 0 176364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1917
timestamp 1676037725
transform 1 0 177468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1929
timestamp 1676037725
transform 1 0 178572 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1941
timestamp 1676037725
transform 1 0 179676 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1953
timestamp 1676037725
transform 1 0 180780 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1959
timestamp 1676037725
transform 1 0 181332 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1961
timestamp 1676037725
transform 1 0 181516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1973
timestamp 1676037725
transform 1 0 182620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1985
timestamp 1676037725
transform 1 0 183724 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1997
timestamp 1676037725
transform 1 0 184828 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2009
timestamp 1676037725
transform 1 0 185932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2015
timestamp 1676037725
transform 1 0 186484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_2017
timestamp 1676037725
transform 1 0 186668 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2021
timestamp 1676037725
transform 1 0 187036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2033
timestamp 1676037725
transform 1 0 188140 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2045
timestamp 1676037725
transform 1 0 189244 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2057
timestamp 1676037725
transform 1 0 190348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_2069
timestamp 1676037725
transform 1 0 191452 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2073
timestamp 1676037725
transform 1 0 191820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2085
timestamp 1676037725
transform 1 0 192924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2097
timestamp 1676037725
transform 1 0 194028 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2109
timestamp 1676037725
transform 1 0 195132 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2121
timestamp 1676037725
transform 1 0 196236 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2127
timestamp 1676037725
transform 1 0 196788 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2129
timestamp 1676037725
transform 1 0 196972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2141
timestamp 1676037725
transform 1 0 198076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2153
timestamp 1676037725
transform 1 0 199180 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2165
timestamp 1676037725
transform 1 0 200284 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2177
timestamp 1676037725
transform 1 0 201388 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2183
timestamp 1676037725
transform 1 0 201940 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2185
timestamp 1676037725
transform 1 0 202124 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2191
timestamp 1676037725
transform 1 0 202676 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2203
timestamp 1676037725
transform 1 0 203780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2215
timestamp 1676037725
transform 1 0 204884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2227
timestamp 1676037725
transform 1 0 205988 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2239
timestamp 1676037725
transform 1 0 207092 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2241
timestamp 1676037725
transform 1 0 207276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2253
timestamp 1676037725
transform 1 0 208380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2265
timestamp 1676037725
transform 1 0 209484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2277
timestamp 1676037725
transform 1 0 210588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2289
timestamp 1676037725
transform 1 0 211692 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2295
timestamp 1676037725
transform 1 0 212244 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2297
timestamp 1676037725
transform 1 0 212428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2309
timestamp 1676037725
transform 1 0 213532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2321
timestamp 1676037725
transform 1 0 214636 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2333
timestamp 1676037725
transform 1 0 215740 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2345
timestamp 1676037725
transform 1 0 216844 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2351
timestamp 1676037725
transform 1 0 217396 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2353
timestamp 1676037725
transform 1 0 217580 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2359
timestamp 1676037725
transform 1 0 218132 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2371
timestamp 1676037725
transform 1 0 219236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2383
timestamp 1676037725
transform 1 0 220340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2395
timestamp 1676037725
transform 1 0 221444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2407
timestamp 1676037725
transform 1 0 222548 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2409
timestamp 1676037725
transform 1 0 222732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2421
timestamp 1676037725
transform 1 0 223836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2433
timestamp 1676037725
transform 1 0 224940 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2445
timestamp 1676037725
transform 1 0 226044 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2457
timestamp 1676037725
transform 1 0 227148 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2463
timestamp 1676037725
transform 1 0 227700 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2465
timestamp 1676037725
transform 1 0 227884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2477
timestamp 1676037725
transform 1 0 228988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2489
timestamp 1676037725
transform 1 0 230092 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2501
timestamp 1676037725
transform 1 0 231196 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2513
timestamp 1676037725
transform 1 0 232300 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2519
timestamp 1676037725
transform 1 0 232852 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2521
timestamp 1676037725
transform 1 0 233036 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2527
timestamp 1676037725
transform 1 0 233588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2539
timestamp 1676037725
transform 1 0 234692 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2551
timestamp 1676037725
transform 1 0 235796 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2563
timestamp 1676037725
transform 1 0 236900 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2575
timestamp 1676037725
transform 1 0 238004 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2577
timestamp 1676037725
transform 1 0 238188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2589
timestamp 1676037725
transform 1 0 239292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2601
timestamp 1676037725
transform 1 0 240396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2613
timestamp 1676037725
transform 1 0 241500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2625
timestamp 1676037725
transform 1 0 242604 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2631
timestamp 1676037725
transform 1 0 243156 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2633
timestamp 1676037725
transform 1 0 243340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2645
timestamp 1676037725
transform 1 0 244444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2657
timestamp 1676037725
transform 1 0 245548 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2669
timestamp 1676037725
transform 1 0 246652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2681
timestamp 1676037725
transform 1 0 247756 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2687
timestamp 1676037725
transform 1 0 248308 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2689
timestamp 1676037725
transform 1 0 248492 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2695
timestamp 1676037725
transform 1 0 249044 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2707
timestamp 1676037725
transform 1 0 250148 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2719
timestamp 1676037725
transform 1 0 251252 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2731
timestamp 1676037725
transform 1 0 252356 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2743
timestamp 1676037725
transform 1 0 253460 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2745
timestamp 1676037725
transform 1 0 253644 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2757
timestamp 1676037725
transform 1 0 254748 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2769
timestamp 1676037725
transform 1 0 255852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2781
timestamp 1676037725
transform 1 0 256956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2793
timestamp 1676037725
transform 1 0 258060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2799
timestamp 1676037725
transform 1 0 258612 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2801
timestamp 1676037725
transform 1 0 258796 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2813
timestamp 1676037725
transform 1 0 259900 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2825
timestamp 1676037725
transform 1 0 261004 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2837
timestamp 1676037725
transform 1 0 262108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2849
timestamp 1676037725
transform 1 0 263212 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2855
timestamp 1676037725
transform 1 0 263764 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2857
timestamp 1676037725
transform 1 0 263948 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2863
timestamp 1676037725
transform 1 0 264500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2875
timestamp 1676037725
transform 1 0 265604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2887
timestamp 1676037725
transform 1 0 266708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2899
timestamp 1676037725
transform 1 0 267812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2911
timestamp 1676037725
transform 1 0 268916 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2913
timestamp 1676037725
transform 1 0 269100 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2925
timestamp 1676037725
transform 1 0 270204 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2937
timestamp 1676037725
transform 1 0 271308 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2949
timestamp 1676037725
transform 1 0 272412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2961
timestamp 1676037725
transform 1 0 273516 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2967
timestamp 1676037725
transform 1 0 274068 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2969
timestamp 1676037725
transform 1 0 274252 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2981
timestamp 1676037725
transform 1 0 275356 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2993
timestamp 1676037725
transform 1 0 276460 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3005
timestamp 1676037725
transform 1 0 277564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3017
timestamp 1676037725
transform 1 0 278668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3023
timestamp 1676037725
transform 1 0 279220 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3025
timestamp 1676037725
transform 1 0 279404 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3029
timestamp 1676037725
transform 1 0 279772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3041
timestamp 1676037725
transform 1 0 280876 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3053
timestamp 1676037725
transform 1 0 281980 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3065
timestamp 1676037725
transform 1 0 283084 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3077
timestamp 1676037725
transform 1 0 284188 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3081
timestamp 1676037725
transform 1 0 284556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3093
timestamp 1676037725
transform 1 0 285660 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3105
timestamp 1676037725
transform 1 0 286764 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3117
timestamp 1676037725
transform 1 0 287868 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3129
timestamp 1676037725
transform 1 0 288972 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3135
timestamp 1676037725
transform 1 0 289524 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3137
timestamp 1676037725
transform 1 0 289708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3149
timestamp 1676037725
transform 1 0 290812 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3161
timestamp 1676037725
transform 1 0 291916 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3173
timestamp 1676037725
transform 1 0 293020 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3185
timestamp 1676037725
transform 1 0 294124 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3191
timestamp 1676037725
transform 1 0 294676 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3193
timestamp 1676037725
transform 1 0 294860 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3199
timestamp 1676037725
transform 1 0 295412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3211
timestamp 1676037725
transform 1 0 296516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3223
timestamp 1676037725
transform 1 0 297620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3235
timestamp 1676037725
transform 1 0 298724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3247
timestamp 1676037725
transform 1 0 299828 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3249
timestamp 1676037725
transform 1 0 300012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3261
timestamp 1676037725
transform 1 0 301116 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3273
timestamp 1676037725
transform 1 0 302220 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3285
timestamp 1676037725
transform 1 0 303324 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3293
timestamp 1676037725
transform 1 0 304060 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3300
timestamp 1676037725
transform 1 0 304704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3305
timestamp 1676037725
transform 1 0 305164 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3309
timestamp 1676037725
transform 1 0 305532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3321
timestamp 1676037725
transform 1 0 306636 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3333
timestamp 1676037725
transform 1 0 307740 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3345
timestamp 1676037725
transform 1 0 308844 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3357
timestamp 1676037725
transform 1 0 309948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3361
timestamp 1676037725
transform 1 0 310316 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3367
timestamp 1676037725
transform 1 0 310868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3379
timestamp 1676037725
transform 1 0 311972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3391
timestamp 1676037725
transform 1 0 313076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3403
timestamp 1676037725
transform 1 0 314180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3415
timestamp 1676037725
transform 1 0 315284 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3417
timestamp 1676037725
transform 1 0 315468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3429
timestamp 1676037725
transform 1 0 316572 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3441
timestamp 1676037725
transform 1 0 317676 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3453
timestamp 1676037725
transform 1 0 318780 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3465
timestamp 1676037725
transform 1 0 319884 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3471
timestamp 1676037725
transform 1 0 320436 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3473
timestamp 1676037725
transform 1 0 320620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3485
timestamp 1676037725
transform 1 0 321724 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3497
timestamp 1676037725
transform 1 0 322828 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3509
timestamp 1676037725
transform 1 0 323932 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3521
timestamp 1676037725
transform 1 0 325036 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3527
timestamp 1676037725
transform 1 0 325588 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3529
timestamp 1676037725
transform 1 0 325772 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3535
timestamp 1676037725
transform 1 0 326324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3547
timestamp 1676037725
transform 1 0 327428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3559
timestamp 1676037725
transform 1 0 328532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3571
timestamp 1676037725
transform 1 0 329636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3583
timestamp 1676037725
transform 1 0 330740 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3585
timestamp 1676037725
transform 1 0 330924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3597
timestamp 1676037725
transform 1 0 332028 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3609
timestamp 1676037725
transform 1 0 333132 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3621
timestamp 1676037725
transform 1 0 334236 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3633
timestamp 1676037725
transform 1 0 335340 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3639
timestamp 1676037725
transform 1 0 335892 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3641
timestamp 1676037725
transform 1 0 336076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3653
timestamp 1676037725
transform 1 0 337180 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3665
timestamp 1676037725
transform 1 0 338284 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3677
timestamp 1676037725
transform 1 0 339388 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3689
timestamp 1676037725
transform 1 0 340492 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3695
timestamp 1676037725
transform 1 0 341044 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3697
timestamp 1676037725
transform 1 0 341228 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3703
timestamp 1676037725
transform 1 0 341780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3715
timestamp 1676037725
transform 1 0 342884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3727
timestamp 1676037725
transform 1 0 343988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3739
timestamp 1676037725
transform 1 0 345092 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3751
timestamp 1676037725
transform 1 0 346196 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3753
timestamp 1676037725
transform 1 0 346380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3765
timestamp 1676037725
transform 1 0 347484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3777
timestamp 1676037725
transform 1 0 348588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3789
timestamp 1676037725
transform 1 0 349692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3801
timestamp 1676037725
transform 1 0 350796 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3807
timestamp 1676037725
transform 1 0 351348 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3809
timestamp 1676037725
transform 1 0 351532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3821
timestamp 1676037725
transform 1 0 352636 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3833
timestamp 1676037725
transform 1 0 353740 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3845
timestamp 1676037725
transform 1 0 354844 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3857
timestamp 1676037725
transform 1 0 355948 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3863
timestamp 1676037725
transform 1 0 356500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3865
timestamp 1676037725
transform 1 0 356684 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3871
timestamp 1676037725
transform 1 0 357236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3883
timestamp 1676037725
transform 1 0 358340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3895
timestamp 1676037725
transform 1 0 359444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3907
timestamp 1676037725
transform 1 0 360548 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3919
timestamp 1676037725
transform 1 0 361652 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3921
timestamp 1676037725
transform 1 0 361836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3933
timestamp 1676037725
transform 1 0 362940 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3945
timestamp 1676037725
transform 1 0 364044 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3957
timestamp 1676037725
transform 1 0 365148 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3969
timestamp 1676037725
transform 1 0 366252 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3975
timestamp 1676037725
transform 1 0 366804 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3977
timestamp 1676037725
transform 1 0 366988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3989
timestamp 1676037725
transform 1 0 368092 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4001
timestamp 1676037725
transform 1 0 369196 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4013
timestamp 1676037725
transform 1 0 370300 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4025
timestamp 1676037725
transform 1 0 371404 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4031
timestamp 1676037725
transform 1 0 371956 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_4033
timestamp 1676037725
transform 1 0 372140 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4039
timestamp 1676037725
transform 1 0 372692 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4051
timestamp 1676037725
transform 1 0 373796 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4063
timestamp 1676037725
transform 1 0 374900 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4075
timestamp 1676037725
transform 1 0 376004 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4087
timestamp 1676037725
transform 1 0 377108 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4089
timestamp 1676037725
transform 1 0 377292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4101
timestamp 1676037725
transform 1 0 378396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4113
timestamp 1676037725
transform 1 0 379500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4125
timestamp 1676037725
transform 1 0 380604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4137
timestamp 1676037725
transform 1 0 381708 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4143
timestamp 1676037725
transform 1 0 382260 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4145
timestamp 1676037725
transform 1 0 382444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4157
timestamp 1676037725
transform 1 0 383548 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4169
timestamp 1676037725
transform 1 0 384652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4181
timestamp 1676037725
transform 1 0 385756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4193
timestamp 1676037725
transform 1 0 386860 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4199
timestamp 1676037725
transform 1 0 387412 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_4201
timestamp 1676037725
transform 1 0 387596 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4207
timestamp 1676037725
transform 1 0 388148 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4219
timestamp 1676037725
transform 1 0 389252 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4231
timestamp 1676037725
transform 1 0 390356 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4243
timestamp 1676037725
transform 1 0 391460 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4255
timestamp 1676037725
transform 1 0 392564 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4257
timestamp 1676037725
transform 1 0 392748 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4269
timestamp 1676037725
transform 1 0 393852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4281
timestamp 1676037725
transform 1 0 394956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4293
timestamp 1676037725
transform 1 0 396060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4305
timestamp 1676037725
transform 1 0 397164 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4311
timestamp 1676037725
transform 1 0 397716 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4313
timestamp 1676037725
transform 1 0 397900 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4325
timestamp 1676037725
transform 1 0 399004 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_4337
timestamp 1676037725
transform 1 0 400108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4341
timestamp 1676037725
transform 1 0 400476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_4348
timestamp 1676037725
transform 1 0 401120 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4354
timestamp 1676037725
transform 1 0 401672 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_4366
timestamp 1676037725
transform 1 0 402776 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_4369
timestamp 1676037725
transform 1 0 403052 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4373
timestamp 1676037725
transform 1 0 403420 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4385
timestamp 1676037725
transform 1 0 404524 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4397
timestamp 1676037725
transform 1 0 405628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4409
timestamp 1676037725
transform 1 0 406732 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_4421
timestamp 1676037725
transform 1 0 407836 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4425
timestamp 1676037725
transform 1 0 408204 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4437
timestamp 1676037725
transform 1 0 409308 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4449
timestamp 1676037725
transform 1 0 410412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4461
timestamp 1676037725
transform 1 0 411516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4473
timestamp 1676037725
transform 1 0 412620 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4479
timestamp 1676037725
transform 1 0 413172 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4481
timestamp 1676037725
transform 1 0 413356 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4493
timestamp 1676037725
transform 1 0 414460 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4505
timestamp 1676037725
transform 1 0 415564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4517
timestamp 1676037725
transform 1 0 416668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4529
timestamp 1676037725
transform 1 0 417772 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4535
timestamp 1676037725
transform 1 0 418324 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4537
timestamp 1676037725
transform 1 0 418508 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4549
timestamp 1676037725
transform 1 0 419612 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4561
timestamp 1676037725
transform 1 0 420716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4573
timestamp 1676037725
transform 1 0 421820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4585
timestamp 1676037725
transform 1 0 422924 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4591
timestamp 1676037725
transform 1 0 423476 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4593
timestamp 1676037725
transform 1 0 423660 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4605
timestamp 1676037725
transform 1 0 424764 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4617
timestamp 1676037725
transform 1 0 425868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4629
timestamp 1676037725
transform 1 0 426972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4641
timestamp 1676037725
transform 1 0 428076 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4647
timestamp 1676037725
transform 1 0 428628 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4649
timestamp 1676037725
transform 1 0 428812 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4661
timestamp 1676037725
transform 1 0 429916 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4673
timestamp 1676037725
transform 1 0 431020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4685
timestamp 1676037725
transform 1 0 432124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4697
timestamp 1676037725
transform 1 0 433228 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4703
timestamp 1676037725
transform 1 0 433780 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_4705
timestamp 1676037725
transform 1 0 433964 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4711
timestamp 1676037725
transform 1 0 434516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4723
timestamp 1676037725
transform 1 0 435620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4735
timestamp 1676037725
transform 1 0 436724 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4747
timestamp 1676037725
transform 1 0 437828 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4759
timestamp 1676037725
transform 1 0 438932 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4761
timestamp 1676037725
transform 1 0 439116 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4773
timestamp 1676037725
transform 1 0 440220 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4785
timestamp 1676037725
transform 1 0 441324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4797
timestamp 1676037725
transform 1 0 442428 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4809
timestamp 1676037725
transform 1 0 443532 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4815
timestamp 1676037725
transform 1 0 444084 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4817
timestamp 1676037725
transform 1 0 444268 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4829
timestamp 1676037725
transform 1 0 445372 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4841
timestamp 1676037725
transform 1 0 446476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4853
timestamp 1676037725
transform 1 0 447580 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4865
timestamp 1676037725
transform 1 0 448684 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4871
timestamp 1676037725
transform 1 0 449236 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_4873
timestamp 1676037725
transform 1 0 449420 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4879
timestamp 1676037725
transform 1 0 449972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4891
timestamp 1676037725
transform 1 0 451076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4903
timestamp 1676037725
transform 1 0 452180 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4915
timestamp 1676037725
transform 1 0 453284 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4927
timestamp 1676037725
transform 1 0 454388 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4929
timestamp 1676037725
transform 1 0 454572 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4941
timestamp 1676037725
transform 1 0 455676 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4953
timestamp 1676037725
transform 1 0 456780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4965
timestamp 1676037725
transform 1 0 457884 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4977
timestamp 1676037725
transform 1 0 458988 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4983
timestamp 1676037725
transform 1 0 459540 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4985
timestamp 1676037725
transform 1 0 459724 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4997
timestamp 1676037725
transform 1 0 460828 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5009
timestamp 1676037725
transform 1 0 461932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5021
timestamp 1676037725
transform 1 0 463036 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5033
timestamp 1676037725
transform 1 0 464140 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5039
timestamp 1676037725
transform 1 0 464692 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5041
timestamp 1676037725
transform 1 0 464876 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5047
timestamp 1676037725
transform 1 0 465428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5059
timestamp 1676037725
transform 1 0 466532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5071
timestamp 1676037725
transform 1 0 467636 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5083
timestamp 1676037725
transform 1 0 468740 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5095
timestamp 1676037725
transform 1 0 469844 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5097
timestamp 1676037725
transform 1 0 470028 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5109
timestamp 1676037725
transform 1 0 471132 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5121
timestamp 1676037725
transform 1 0 472236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5133
timestamp 1676037725
transform 1 0 473340 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5145
timestamp 1676037725
transform 1 0 474444 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5151
timestamp 1676037725
transform 1 0 474996 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5153
timestamp 1676037725
transform 1 0 475180 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5165
timestamp 1676037725
transform 1 0 476284 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5177
timestamp 1676037725
transform 1 0 477388 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5189
timestamp 1676037725
transform 1 0 478492 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5201
timestamp 1676037725
transform 1 0 479596 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5207
timestamp 1676037725
transform 1 0 480148 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5209
timestamp 1676037725
transform 1 0 480332 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5215
timestamp 1676037725
transform 1 0 480884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5227
timestamp 1676037725
transform 1 0 481988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5239
timestamp 1676037725
transform 1 0 483092 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5251
timestamp 1676037725
transform 1 0 484196 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5263
timestamp 1676037725
transform 1 0 485300 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5265
timestamp 1676037725
transform 1 0 485484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5277
timestamp 1676037725
transform 1 0 486588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5289
timestamp 1676037725
transform 1 0 487692 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5301
timestamp 1676037725
transform 1 0 488796 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5313
timestamp 1676037725
transform 1 0 489900 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5319
timestamp 1676037725
transform 1 0 490452 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5321
timestamp 1676037725
transform 1 0 490636 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5333
timestamp 1676037725
transform 1 0 491740 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5345
timestamp 1676037725
transform 1 0 492844 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5357
timestamp 1676037725
transform 1 0 493948 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5369
timestamp 1676037725
transform 1 0 495052 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5375
timestamp 1676037725
transform 1 0 495604 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5377
timestamp 1676037725
transform 1 0 495788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_5383
timestamp 1676037725
transform 1 0 496340 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5397
timestamp 1676037725
transform 1 0 497628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5409
timestamp 1676037725
transform 1 0 498732 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_5421
timestamp 1676037725
transform 1 0 499836 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_5429
timestamp 1676037725
transform 1 0 500572 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5433
timestamp 1676037725
transform 1 0 500940 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5445
timestamp 1676037725
transform 1 0 502044 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5457
timestamp 1676037725
transform 1 0 503148 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5469
timestamp 1676037725
transform 1 0 504252 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5481
timestamp 1676037725
transform 1 0 505356 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5487
timestamp 1676037725
transform 1 0 505908 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5489
timestamp 1676037725
transform 1 0 506092 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5501
timestamp 1676037725
transform 1 0 507196 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5513
timestamp 1676037725
transform 1 0 508300 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5525
timestamp 1676037725
transform 1 0 509404 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5537
timestamp 1676037725
transform 1 0 510508 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5543
timestamp 1676037725
transform 1 0 511060 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5545
timestamp 1676037725
transform 1 0 511244 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5557
timestamp 1676037725
transform 1 0 512348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5569
timestamp 1676037725
transform 1 0 513452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5581
timestamp 1676037725
transform 1 0 514556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5593
timestamp 1676037725
transform 1 0 515660 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5599
timestamp 1676037725
transform 1 0 516212 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5601
timestamp 1676037725
transform 1 0 516396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5613
timestamp 1676037725
transform 1 0 517500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5625
timestamp 1676037725
transform 1 0 518604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5637
timestamp 1676037725
transform 1 0 519708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5649
timestamp 1676037725
transform 1 0 520812 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5655
timestamp 1676037725
transform 1 0 521364 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5657
timestamp 1676037725
transform 1 0 521548 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5669
timestamp 1676037725
transform 1 0 522652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5681
timestamp 1676037725
transform 1 0 523756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5693
timestamp 1676037725
transform 1 0 524860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5705
timestamp 1676037725
transform 1 0 525964 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5711
timestamp 1676037725
transform 1 0 526516 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5713
timestamp 1676037725
transform 1 0 526700 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5719
timestamp 1676037725
transform 1 0 527252 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5731
timestamp 1676037725
transform 1 0 528356 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5743
timestamp 1676037725
transform 1 0 529460 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5755
timestamp 1676037725
transform 1 0 530564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5767
timestamp 1676037725
transform 1 0 531668 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5769
timestamp 1676037725
transform 1 0 531852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5781
timestamp 1676037725
transform 1 0 532956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5793
timestamp 1676037725
transform 1 0 534060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5805
timestamp 1676037725
transform 1 0 535164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5817
timestamp 1676037725
transform 1 0 536268 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5823
timestamp 1676037725
transform 1 0 536820 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5825
timestamp 1676037725
transform 1 0 537004 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5837
timestamp 1676037725
transform 1 0 538108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5849
timestamp 1676037725
transform 1 0 539212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5861
timestamp 1676037725
transform 1 0 540316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5873
timestamp 1676037725
transform 1 0 541420 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5879
timestamp 1676037725
transform 1 0 541972 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5881
timestamp 1676037725
transform 1 0 542156 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5887
timestamp 1676037725
transform 1 0 542708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5899
timestamp 1676037725
transform 1 0 543812 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5911
timestamp 1676037725
transform 1 0 544916 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5923
timestamp 1676037725
transform 1 0 546020 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5935
timestamp 1676037725
transform 1 0 547124 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5937
timestamp 1676037725
transform 1 0 547308 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5949
timestamp 1676037725
transform 1 0 548412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5961
timestamp 1676037725
transform 1 0 549516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5973
timestamp 1676037725
transform 1 0 550620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5985
timestamp 1676037725
transform 1 0 551724 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5991
timestamp 1676037725
transform 1 0 552276 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5993
timestamp 1676037725
transform 1 0 552460 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6005
timestamp 1676037725
transform 1 0 553564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6017
timestamp 1676037725
transform 1 0 554668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6029
timestamp 1676037725
transform 1 0 555772 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6041
timestamp 1676037725
transform 1 0 556876 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6047
timestamp 1676037725
transform 1 0 557428 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_6049
timestamp 1676037725
transform 1 0 557612 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6055
timestamp 1676037725
transform 1 0 558164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6067
timestamp 1676037725
transform 1 0 559268 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6079
timestamp 1676037725
transform 1 0 560372 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6091
timestamp 1676037725
transform 1 0 561476 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6103
timestamp 1676037725
transform 1 0 562580 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6105
timestamp 1676037725
transform 1 0 562764 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6117
timestamp 1676037725
transform 1 0 563868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6129
timestamp 1676037725
transform 1 0 564972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6141
timestamp 1676037725
transform 1 0 566076 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6153
timestamp 1676037725
transform 1 0 567180 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6159
timestamp 1676037725
transform 1 0 567732 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6161
timestamp 1676037725
transform 1 0 567916 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6173
timestamp 1676037725
transform 1 0 569020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6185
timestamp 1676037725
transform 1 0 570124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6197
timestamp 1676037725
transform 1 0 571228 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6209
timestamp 1676037725
transform 1 0 572332 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6215
timestamp 1676037725
transform 1 0 572884 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_6217
timestamp 1676037725
transform 1 0 573068 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6223
timestamp 1676037725
transform 1 0 573620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6235
timestamp 1676037725
transform 1 0 574724 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6247
timestamp 1676037725
transform 1 0 575828 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6259
timestamp 1676037725
transform 1 0 576932 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6271
timestamp 1676037725
transform 1 0 578036 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6273
timestamp 1676037725
transform 1 0 578220 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6285
timestamp 1676037725
transform 1 0 579324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6297
timestamp 1676037725
transform 1 0 580428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6309
timestamp 1676037725
transform 1 0 581532 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6321
timestamp 1676037725
transform 1 0 582636 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6327
timestamp 1676037725
transform 1 0 583188 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6329
timestamp 1676037725
transform 1 0 583372 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6341
timestamp 1676037725
transform 1 0 584476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6353
timestamp 1676037725
transform 1 0 585580 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6365
timestamp 1676037725
transform 1 0 586684 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6377
timestamp 1676037725
transform 1 0 587788 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6383
timestamp 1676037725
transform 1 0 588340 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_6385
timestamp 1676037725
transform 1 0 588524 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6391
timestamp 1676037725
transform 1 0 589076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6403
timestamp 1676037725
transform 1 0 590180 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6415
timestamp 1676037725
transform 1 0 591284 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6427
timestamp 1676037725
transform 1 0 592388 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6439
timestamp 1676037725
transform 1 0 593492 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_6441
timestamp 1676037725
transform 1 0 593676 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6449
timestamp 1676037725
transform 1 0 594412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6461
timestamp 1676037725
transform 1 0 595516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6473
timestamp 1676037725
transform 1 0 596620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_6485
timestamp 1676037725
transform 1 0 597724 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_6493
timestamp 1676037725
transform 1 0 598460 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6497
timestamp 1676037725
transform 1 0 598828 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6509
timestamp 1676037725
transform 1 0 599932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6521
timestamp 1676037725
transform 1 0 601036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6533
timestamp 1676037725
transform 1 0 602140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6545
timestamp 1676037725
transform 1 0 603244 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6551
timestamp 1676037725
transform 1 0 603796 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6553
timestamp 1676037725
transform 1 0 603980 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6565
timestamp 1676037725
transform 1 0 605084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6577
timestamp 1676037725
transform 1 0 606188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6589
timestamp 1676037725
transform 1 0 607292 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6601
timestamp 1676037725
transform 1 0 608396 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6607
timestamp 1676037725
transform 1 0 608948 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6609
timestamp 1676037725
transform 1 0 609132 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6621
timestamp 1676037725
transform 1 0 610236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6633
timestamp 1676037725
transform 1 0 611340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6645
timestamp 1676037725
transform 1 0 612444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6657
timestamp 1676037725
transform 1 0 613548 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6663
timestamp 1676037725
transform 1 0 614100 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6665
timestamp 1676037725
transform 1 0 614284 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6677
timestamp 1676037725
transform 1 0 615388 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6689
timestamp 1676037725
transform 1 0 616492 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6701
timestamp 1676037725
transform 1 0 617596 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6713
timestamp 1676037725
transform 1 0 618700 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6719
timestamp 1676037725
transform 1 0 619252 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_6721
timestamp 1676037725
transform 1 0 619436 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6727
timestamp 1676037725
transform 1 0 619988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6739
timestamp 1676037725
transform 1 0 621092 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6751
timestamp 1676037725
transform 1 0 622196 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6763
timestamp 1676037725
transform 1 0 623300 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6775
timestamp 1676037725
transform 1 0 624404 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6777
timestamp 1676037725
transform 1 0 624588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6789
timestamp 1676037725
transform 1 0 625692 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6801
timestamp 1676037725
transform 1 0 626796 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6813
timestamp 1676037725
transform 1 0 627900 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6825
timestamp 1676037725
transform 1 0 629004 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6831
timestamp 1676037725
transform 1 0 629556 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6833
timestamp 1676037725
transform 1 0 629740 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6845
timestamp 1676037725
transform 1 0 630844 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6857
timestamp 1676037725
transform 1 0 631948 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6869
timestamp 1676037725
transform 1 0 633052 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6881
timestamp 1676037725
transform 1 0 634156 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6887
timestamp 1676037725
transform 1 0 634708 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_6889
timestamp 1676037725
transform 1 0 634892 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6895
timestamp 1676037725
transform 1 0 635444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6907
timestamp 1676037725
transform 1 0 636548 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6919
timestamp 1676037725
transform 1 0 637652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6931
timestamp 1676037725
transform 1 0 638756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6943
timestamp 1676037725
transform 1 0 639860 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6945
timestamp 1676037725
transform 1 0 640044 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6957
timestamp 1676037725
transform 1 0 641148 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6969
timestamp 1676037725
transform 1 0 642252 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6981
timestamp 1676037725
transform 1 0 643356 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6993
timestamp 1676037725
transform 1 0 644460 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6999
timestamp 1676037725
transform 1 0 645012 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7001
timestamp 1676037725
transform 1 0 645196 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7013
timestamp 1676037725
transform 1 0 646300 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7025
timestamp 1676037725
transform 1 0 647404 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7037
timestamp 1676037725
transform 1 0 648508 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1676037725
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1676037725
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1676037725
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1676037725
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1676037725
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1676037725
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1676037725
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1676037725
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1676037725
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1676037725
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1676037725
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1676037725
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1676037725
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1676037725
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1676037725
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1676037725
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1676037725
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1676037725
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1676037725
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1676037725
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1676037725
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1676037725
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1676037725
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_625
timestamp 1676037725
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1676037725
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1676037725
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1676037725
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1676037725
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1676037725
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1676037725
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 1676037725
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1676037725
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1676037725
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1676037725
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1676037725
transform 1 0 67804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_737
timestamp 1676037725
transform 1 0 68908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 1676037725
transform 1 0 70012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1676037725
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_757
timestamp 1676037725
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_769
timestamp 1676037725
transform 1 0 71852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_781
timestamp 1676037725
transform 1 0 72956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_793
timestamp 1676037725
transform 1 0 74060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 1676037725
transform 1 0 75164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 1676037725
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_813
timestamp 1676037725
transform 1 0 75900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_825
timestamp 1676037725
transform 1 0 77004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_837
timestamp 1676037725
transform 1 0 78108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_849
timestamp 1676037725
transform 1 0 79212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_861
timestamp 1676037725
transform 1 0 80316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_867
timestamp 1676037725
transform 1 0 80868 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_869
timestamp 1676037725
transform 1 0 81052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_881
timestamp 1676037725
transform 1 0 82156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_893
timestamp 1676037725
transform 1 0 83260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_905
timestamp 1676037725
transform 1 0 84364 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_917
timestamp 1676037725
transform 1 0 85468 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_923
timestamp 1676037725
transform 1 0 86020 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_925
timestamp 1676037725
transform 1 0 86204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_937
timestamp 1676037725
transform 1 0 87308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_949
timestamp 1676037725
transform 1 0 88412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_961
timestamp 1676037725
transform 1 0 89516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_973
timestamp 1676037725
transform 1 0 90620 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_979
timestamp 1676037725
transform 1 0 91172 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_981
timestamp 1676037725
transform 1 0 91356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_993
timestamp 1676037725
transform 1 0 92460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1005
timestamp 1676037725
transform 1 0 93564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1017
timestamp 1676037725
transform 1 0 94668 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1029
timestamp 1676037725
transform 1 0 95772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1035
timestamp 1676037725
transform 1 0 96324 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1037
timestamp 1676037725
transform 1 0 96508 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1049
timestamp 1676037725
transform 1 0 97612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1061
timestamp 1676037725
transform 1 0 98716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1073
timestamp 1676037725
transform 1 0 99820 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1085
timestamp 1676037725
transform 1 0 100924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1091
timestamp 1676037725
transform 1 0 101476 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1093
timestamp 1676037725
transform 1 0 101660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1105
timestamp 1676037725
transform 1 0 102764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1117
timestamp 1676037725
transform 1 0 103868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1129
timestamp 1676037725
transform 1 0 104972 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1141
timestamp 1676037725
transform 1 0 106076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1147
timestamp 1676037725
transform 1 0 106628 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1149
timestamp 1676037725
transform 1 0 106812 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1161
timestamp 1676037725
transform 1 0 107916 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1173
timestamp 1676037725
transform 1 0 109020 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1185
timestamp 1676037725
transform 1 0 110124 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1197
timestamp 1676037725
transform 1 0 111228 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1203
timestamp 1676037725
transform 1 0 111780 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1205
timestamp 1676037725
transform 1 0 111964 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1217
timestamp 1676037725
transform 1 0 113068 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1229
timestamp 1676037725
transform 1 0 114172 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1241
timestamp 1676037725
transform 1 0 115276 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1253
timestamp 1676037725
transform 1 0 116380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1259
timestamp 1676037725
transform 1 0 116932 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1261
timestamp 1676037725
transform 1 0 117116 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1273
timestamp 1676037725
transform 1 0 118220 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1285
timestamp 1676037725
transform 1 0 119324 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1297
timestamp 1676037725
transform 1 0 120428 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1309
timestamp 1676037725
transform 1 0 121532 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1315
timestamp 1676037725
transform 1 0 122084 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1317
timestamp 1676037725
transform 1 0 122268 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1329
timestamp 1676037725
transform 1 0 123372 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1341
timestamp 1676037725
transform 1 0 124476 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1353
timestamp 1676037725
transform 1 0 125580 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1365
timestamp 1676037725
transform 1 0 126684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1371
timestamp 1676037725
transform 1 0 127236 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1373
timestamp 1676037725
transform 1 0 127420 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1385
timestamp 1676037725
transform 1 0 128524 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1397
timestamp 1676037725
transform 1 0 129628 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1409
timestamp 1676037725
transform 1 0 130732 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1421
timestamp 1676037725
transform 1 0 131836 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1427
timestamp 1676037725
transform 1 0 132388 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1429
timestamp 1676037725
transform 1 0 132572 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1441
timestamp 1676037725
transform 1 0 133676 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1453
timestamp 1676037725
transform 1 0 134780 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1465
timestamp 1676037725
transform 1 0 135884 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1477
timestamp 1676037725
transform 1 0 136988 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1483
timestamp 1676037725
transform 1 0 137540 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1485
timestamp 1676037725
transform 1 0 137724 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1497
timestamp 1676037725
transform 1 0 138828 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1509
timestamp 1676037725
transform 1 0 139932 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1521
timestamp 1676037725
transform 1 0 141036 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1533
timestamp 1676037725
transform 1 0 142140 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1539
timestamp 1676037725
transform 1 0 142692 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1541
timestamp 1676037725
transform 1 0 142876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1553
timestamp 1676037725
transform 1 0 143980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1565
timestamp 1676037725
transform 1 0 145084 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1577
timestamp 1676037725
transform 1 0 146188 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1589
timestamp 1676037725
transform 1 0 147292 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1595
timestamp 1676037725
transform 1 0 147844 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1597
timestamp 1676037725
transform 1 0 148028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1609
timestamp 1676037725
transform 1 0 149132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1621
timestamp 1676037725
transform 1 0 150236 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1633
timestamp 1676037725
transform 1 0 151340 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1645
timestamp 1676037725
transform 1 0 152444 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1651
timestamp 1676037725
transform 1 0 152996 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1653
timestamp 1676037725
transform 1 0 153180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1665
timestamp 1676037725
transform 1 0 154284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1677
timestamp 1676037725
transform 1 0 155388 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1689
timestamp 1676037725
transform 1 0 156492 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1701
timestamp 1676037725
transform 1 0 157596 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1707
timestamp 1676037725
transform 1 0 158148 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1709
timestamp 1676037725
transform 1 0 158332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1721
timestamp 1676037725
transform 1 0 159436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1733
timestamp 1676037725
transform 1 0 160540 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1745
timestamp 1676037725
transform 1 0 161644 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1757
timestamp 1676037725
transform 1 0 162748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1763
timestamp 1676037725
transform 1 0 163300 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1765
timestamp 1676037725
transform 1 0 163484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1777
timestamp 1676037725
transform 1 0 164588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1789
timestamp 1676037725
transform 1 0 165692 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1801
timestamp 1676037725
transform 1 0 166796 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1813
timestamp 1676037725
transform 1 0 167900 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1819
timestamp 1676037725
transform 1 0 168452 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1821
timestamp 1676037725
transform 1 0 168636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1833
timestamp 1676037725
transform 1 0 169740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1845
timestamp 1676037725
transform 1 0 170844 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1857
timestamp 1676037725
transform 1 0 171948 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1869
timestamp 1676037725
transform 1 0 173052 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1875
timestamp 1676037725
transform 1 0 173604 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1877
timestamp 1676037725
transform 1 0 173788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1889
timestamp 1676037725
transform 1 0 174892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1901
timestamp 1676037725
transform 1 0 175996 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1913
timestamp 1676037725
transform 1 0 177100 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1925
timestamp 1676037725
transform 1 0 178204 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1931
timestamp 1676037725
transform 1 0 178756 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1933
timestamp 1676037725
transform 1 0 178940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1945
timestamp 1676037725
transform 1 0 180044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1957
timestamp 1676037725
transform 1 0 181148 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1969
timestamp 1676037725
transform 1 0 182252 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1981
timestamp 1676037725
transform 1 0 183356 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1987
timestamp 1676037725
transform 1 0 183908 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1989
timestamp 1676037725
transform 1 0 184092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2001
timestamp 1676037725
transform 1 0 185196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2013
timestamp 1676037725
transform 1 0 186300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2025
timestamp 1676037725
transform 1 0 187404 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2037
timestamp 1676037725
transform 1 0 188508 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2043
timestamp 1676037725
transform 1 0 189060 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2045
timestamp 1676037725
transform 1 0 189244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2057
timestamp 1676037725
transform 1 0 190348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2069
timestamp 1676037725
transform 1 0 191452 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2081
timestamp 1676037725
transform 1 0 192556 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2093
timestamp 1676037725
transform 1 0 193660 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2099
timestamp 1676037725
transform 1 0 194212 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2101
timestamp 1676037725
transform 1 0 194396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2113
timestamp 1676037725
transform 1 0 195500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2125
timestamp 1676037725
transform 1 0 196604 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2137
timestamp 1676037725
transform 1 0 197708 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2149
timestamp 1676037725
transform 1 0 198812 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2155
timestamp 1676037725
transform 1 0 199364 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2157
timestamp 1676037725
transform 1 0 199548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2169
timestamp 1676037725
transform 1 0 200652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2181
timestamp 1676037725
transform 1 0 201756 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2193
timestamp 1676037725
transform 1 0 202860 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2205
timestamp 1676037725
transform 1 0 203964 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2211
timestamp 1676037725
transform 1 0 204516 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2213
timestamp 1676037725
transform 1 0 204700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2225
timestamp 1676037725
transform 1 0 205804 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_2237
timestamp 1676037725
transform 1 0 206908 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_2245
timestamp 1676037725
transform 1 0 207644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_2254
timestamp 1676037725
transform 1 0 208472 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_2260
timestamp 1676037725
transform 1 0 209024 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2269
timestamp 1676037725
transform 1 0 209852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2281
timestamp 1676037725
transform 1 0 210956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2293
timestamp 1676037725
transform 1 0 212060 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2305
timestamp 1676037725
transform 1 0 213164 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2317
timestamp 1676037725
transform 1 0 214268 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2323
timestamp 1676037725
transform 1 0 214820 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2325
timestamp 1676037725
transform 1 0 215004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2337
timestamp 1676037725
transform 1 0 216108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2349
timestamp 1676037725
transform 1 0 217212 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2361
timestamp 1676037725
transform 1 0 218316 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2373
timestamp 1676037725
transform 1 0 219420 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2379
timestamp 1676037725
transform 1 0 219972 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2381
timestamp 1676037725
transform 1 0 220156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2393
timestamp 1676037725
transform 1 0 221260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2405
timestamp 1676037725
transform 1 0 222364 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2417
timestamp 1676037725
transform 1 0 223468 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2429
timestamp 1676037725
transform 1 0 224572 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2435
timestamp 1676037725
transform 1 0 225124 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2437
timestamp 1676037725
transform 1 0 225308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2449
timestamp 1676037725
transform 1 0 226412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2461
timestamp 1676037725
transform 1 0 227516 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2473
timestamp 1676037725
transform 1 0 228620 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2485
timestamp 1676037725
transform 1 0 229724 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2491
timestamp 1676037725
transform 1 0 230276 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2493
timestamp 1676037725
transform 1 0 230460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2505
timestamp 1676037725
transform 1 0 231564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2517
timestamp 1676037725
transform 1 0 232668 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2529
timestamp 1676037725
transform 1 0 233772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2541
timestamp 1676037725
transform 1 0 234876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2547
timestamp 1676037725
transform 1 0 235428 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2549
timestamp 1676037725
transform 1 0 235612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2561
timestamp 1676037725
transform 1 0 236716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2573
timestamp 1676037725
transform 1 0 237820 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2585
timestamp 1676037725
transform 1 0 238924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2597
timestamp 1676037725
transform 1 0 240028 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2603
timestamp 1676037725
transform 1 0 240580 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2605
timestamp 1676037725
transform 1 0 240764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2617
timestamp 1676037725
transform 1 0 241868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2629
timestamp 1676037725
transform 1 0 242972 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2641
timestamp 1676037725
transform 1 0 244076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2653
timestamp 1676037725
transform 1 0 245180 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2659
timestamp 1676037725
transform 1 0 245732 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2661
timestamp 1676037725
transform 1 0 245916 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2673
timestamp 1676037725
transform 1 0 247020 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2685
timestamp 1676037725
transform 1 0 248124 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2697
timestamp 1676037725
transform 1 0 249228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2709
timestamp 1676037725
transform 1 0 250332 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2715
timestamp 1676037725
transform 1 0 250884 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2717
timestamp 1676037725
transform 1 0 251068 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2729
timestamp 1676037725
transform 1 0 252172 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2741
timestamp 1676037725
transform 1 0 253276 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2753
timestamp 1676037725
transform 1 0 254380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2765
timestamp 1676037725
transform 1 0 255484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2771
timestamp 1676037725
transform 1 0 256036 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2773
timestamp 1676037725
transform 1 0 256220 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2785
timestamp 1676037725
transform 1 0 257324 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2797
timestamp 1676037725
transform 1 0 258428 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2809
timestamp 1676037725
transform 1 0 259532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2821
timestamp 1676037725
transform 1 0 260636 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2827
timestamp 1676037725
transform 1 0 261188 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2829
timestamp 1676037725
transform 1 0 261372 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2841
timestamp 1676037725
transform 1 0 262476 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2853
timestamp 1676037725
transform 1 0 263580 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2865
timestamp 1676037725
transform 1 0 264684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2877
timestamp 1676037725
transform 1 0 265788 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2883
timestamp 1676037725
transform 1 0 266340 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2885
timestamp 1676037725
transform 1 0 266524 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2897
timestamp 1676037725
transform 1 0 267628 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2909
timestamp 1676037725
transform 1 0 268732 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2921
timestamp 1676037725
transform 1 0 269836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2933
timestamp 1676037725
transform 1 0 270940 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2939
timestamp 1676037725
transform 1 0 271492 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2941
timestamp 1676037725
transform 1 0 271676 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2953
timestamp 1676037725
transform 1 0 272780 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2965
timestamp 1676037725
transform 1 0 273884 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2977
timestamp 1676037725
transform 1 0 274988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2989
timestamp 1676037725
transform 1 0 276092 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2995
timestamp 1676037725
transform 1 0 276644 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2997
timestamp 1676037725
transform 1 0 276828 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3009
timestamp 1676037725
transform 1 0 277932 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3021
timestamp 1676037725
transform 1 0 279036 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3033
timestamp 1676037725
transform 1 0 280140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3045
timestamp 1676037725
transform 1 0 281244 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3051
timestamp 1676037725
transform 1 0 281796 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3053
timestamp 1676037725
transform 1 0 281980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3065
timestamp 1676037725
transform 1 0 283084 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3077
timestamp 1676037725
transform 1 0 284188 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3089
timestamp 1676037725
transform 1 0 285292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3101
timestamp 1676037725
transform 1 0 286396 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3107
timestamp 1676037725
transform 1 0 286948 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3109
timestamp 1676037725
transform 1 0 287132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3121
timestamp 1676037725
transform 1 0 288236 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3133
timestamp 1676037725
transform 1 0 289340 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3145
timestamp 1676037725
transform 1 0 290444 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3157
timestamp 1676037725
transform 1 0 291548 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3163
timestamp 1676037725
transform 1 0 292100 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3165
timestamp 1676037725
transform 1 0 292284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3177
timestamp 1676037725
transform 1 0 293388 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3189
timestamp 1676037725
transform 1 0 294492 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3201
timestamp 1676037725
transform 1 0 295596 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3213
timestamp 1676037725
transform 1 0 296700 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3219
timestamp 1676037725
transform 1 0 297252 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3221
timestamp 1676037725
transform 1 0 297436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3233
timestamp 1676037725
transform 1 0 298540 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3245
timestamp 1676037725
transform 1 0 299644 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3257
timestamp 1676037725
transform 1 0 300748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3269
timestamp 1676037725
transform 1 0 301852 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3275
timestamp 1676037725
transform 1 0 302404 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3277
timestamp 1676037725
transform 1 0 302588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3289
timestamp 1676037725
transform 1 0 303692 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3301
timestamp 1676037725
transform 1 0 304796 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3313
timestamp 1676037725
transform 1 0 305900 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3325
timestamp 1676037725
transform 1 0 307004 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3331
timestamp 1676037725
transform 1 0 307556 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3333
timestamp 1676037725
transform 1 0 307740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3345
timestamp 1676037725
transform 1 0 308844 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3357
timestamp 1676037725
transform 1 0 309948 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3369
timestamp 1676037725
transform 1 0 311052 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3381
timestamp 1676037725
transform 1 0 312156 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3387
timestamp 1676037725
transform 1 0 312708 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3389
timestamp 1676037725
transform 1 0 312892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3401
timestamp 1676037725
transform 1 0 313996 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3413
timestamp 1676037725
transform 1 0 315100 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3425
timestamp 1676037725
transform 1 0 316204 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3437
timestamp 1676037725
transform 1 0 317308 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3443
timestamp 1676037725
transform 1 0 317860 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3445
timestamp 1676037725
transform 1 0 318044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3457
timestamp 1676037725
transform 1 0 319148 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3469
timestamp 1676037725
transform 1 0 320252 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3481
timestamp 1676037725
transform 1 0 321356 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3493
timestamp 1676037725
transform 1 0 322460 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3499
timestamp 1676037725
transform 1 0 323012 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3501
timestamp 1676037725
transform 1 0 323196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3513
timestamp 1676037725
transform 1 0 324300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3525
timestamp 1676037725
transform 1 0 325404 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3537
timestamp 1676037725
transform 1 0 326508 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3549
timestamp 1676037725
transform 1 0 327612 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3555
timestamp 1676037725
transform 1 0 328164 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3557
timestamp 1676037725
transform 1 0 328348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3569
timestamp 1676037725
transform 1 0 329452 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3581
timestamp 1676037725
transform 1 0 330556 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3593
timestamp 1676037725
transform 1 0 331660 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3605
timestamp 1676037725
transform 1 0 332764 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3611
timestamp 1676037725
transform 1 0 333316 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3613
timestamp 1676037725
transform 1 0 333500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3625
timestamp 1676037725
transform 1 0 334604 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3637
timestamp 1676037725
transform 1 0 335708 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3649
timestamp 1676037725
transform 1 0 336812 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3661
timestamp 1676037725
transform 1 0 337916 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3667
timestamp 1676037725
transform 1 0 338468 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3669
timestamp 1676037725
transform 1 0 338652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3681
timestamp 1676037725
transform 1 0 339756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3693
timestamp 1676037725
transform 1 0 340860 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3697
timestamp 1676037725
transform 1 0 341228 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3700
timestamp 1676037725
transform 1 0 341504 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3712
timestamp 1676037725
transform 1 0 342608 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3725
timestamp 1676037725
transform 1 0 343804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3737
timestamp 1676037725
transform 1 0 344908 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3749
timestamp 1676037725
transform 1 0 346012 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3761
timestamp 1676037725
transform 1 0 347116 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3773
timestamp 1676037725
transform 1 0 348220 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3779
timestamp 1676037725
transform 1 0 348772 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3781
timestamp 1676037725
transform 1 0 348956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3793
timestamp 1676037725
transform 1 0 350060 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3805
timestamp 1676037725
transform 1 0 351164 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3817
timestamp 1676037725
transform 1 0 352268 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3829
timestamp 1676037725
transform 1 0 353372 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3835
timestamp 1676037725
transform 1 0 353924 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3837
timestamp 1676037725
transform 1 0 354108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3849
timestamp 1676037725
transform 1 0 355212 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3861
timestamp 1676037725
transform 1 0 356316 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3873
timestamp 1676037725
transform 1 0 357420 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3885
timestamp 1676037725
transform 1 0 358524 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3891
timestamp 1676037725
transform 1 0 359076 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3893
timestamp 1676037725
transform 1 0 359260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3905
timestamp 1676037725
transform 1 0 360364 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3917
timestamp 1676037725
transform 1 0 361468 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3929
timestamp 1676037725
transform 1 0 362572 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3941
timestamp 1676037725
transform 1 0 363676 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3947
timestamp 1676037725
transform 1 0 364228 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3949
timestamp 1676037725
transform 1 0 364412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3961
timestamp 1676037725
transform 1 0 365516 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3973
timestamp 1676037725
transform 1 0 366620 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3985
timestamp 1676037725
transform 1 0 367724 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3997
timestamp 1676037725
transform 1 0 368828 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4003
timestamp 1676037725
transform 1 0 369380 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4005
timestamp 1676037725
transform 1 0 369564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4017
timestamp 1676037725
transform 1 0 370668 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4029
timestamp 1676037725
transform 1 0 371772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4041
timestamp 1676037725
transform 1 0 372876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4053
timestamp 1676037725
transform 1 0 373980 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4059
timestamp 1676037725
transform 1 0 374532 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4061
timestamp 1676037725
transform 1 0 374716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4073
timestamp 1676037725
transform 1 0 375820 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4085
timestamp 1676037725
transform 1 0 376924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4097
timestamp 1676037725
transform 1 0 378028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4109
timestamp 1676037725
transform 1 0 379132 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4115
timestamp 1676037725
transform 1 0 379684 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4117
timestamp 1676037725
transform 1 0 379868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4129
timestamp 1676037725
transform 1 0 380972 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4141
timestamp 1676037725
transform 1 0 382076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4153
timestamp 1676037725
transform 1 0 383180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4165
timestamp 1676037725
transform 1 0 384284 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4171
timestamp 1676037725
transform 1 0 384836 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4173
timestamp 1676037725
transform 1 0 385020 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4185
timestamp 1676037725
transform 1 0 386124 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4197
timestamp 1676037725
transform 1 0 387228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4209
timestamp 1676037725
transform 1 0 388332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4221
timestamp 1676037725
transform 1 0 389436 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4227
timestamp 1676037725
transform 1 0 389988 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4229
timestamp 1676037725
transform 1 0 390172 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4241
timestamp 1676037725
transform 1 0 391276 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4253
timestamp 1676037725
transform 1 0 392380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4265
timestamp 1676037725
transform 1 0 393484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4277
timestamp 1676037725
transform 1 0 394588 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4283
timestamp 1676037725
transform 1 0 395140 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4285
timestamp 1676037725
transform 1 0 395324 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4297
timestamp 1676037725
transform 1 0 396428 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4309
timestamp 1676037725
transform 1 0 397532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4321
timestamp 1676037725
transform 1 0 398636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4333
timestamp 1676037725
transform 1 0 399740 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4339
timestamp 1676037725
transform 1 0 400292 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4341
timestamp 1676037725
transform 1 0 400476 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4353
timestamp 1676037725
transform 1 0 401580 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4368
timestamp 1676037725
transform 1 0 402960 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_4383
timestamp 1676037725
transform 1 0 404340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4389
timestamp 1676037725
transform 1 0 404892 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4395
timestamp 1676037725
transform 1 0 405444 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4397
timestamp 1676037725
transform 1 0 405628 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4409
timestamp 1676037725
transform 1 0 406732 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4421
timestamp 1676037725
transform 1 0 407836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4433
timestamp 1676037725
transform 1 0 408940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4445
timestamp 1676037725
transform 1 0 410044 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4451
timestamp 1676037725
transform 1 0 410596 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4453
timestamp 1676037725
transform 1 0 410780 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4465
timestamp 1676037725
transform 1 0 411884 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4477
timestamp 1676037725
transform 1 0 412988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4489
timestamp 1676037725
transform 1 0 414092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4501
timestamp 1676037725
transform 1 0 415196 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4507
timestamp 1676037725
transform 1 0 415748 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4509
timestamp 1676037725
transform 1 0 415932 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4521
timestamp 1676037725
transform 1 0 417036 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4533
timestamp 1676037725
transform 1 0 418140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4545
timestamp 1676037725
transform 1 0 419244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4557
timestamp 1676037725
transform 1 0 420348 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4563
timestamp 1676037725
transform 1 0 420900 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4565
timestamp 1676037725
transform 1 0 421084 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4577
timestamp 1676037725
transform 1 0 422188 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4589
timestamp 1676037725
transform 1 0 423292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4601
timestamp 1676037725
transform 1 0 424396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4613
timestamp 1676037725
transform 1 0 425500 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4619
timestamp 1676037725
transform 1 0 426052 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4621
timestamp 1676037725
transform 1 0 426236 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4633
timestamp 1676037725
transform 1 0 427340 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4645
timestamp 1676037725
transform 1 0 428444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4657
timestamp 1676037725
transform 1 0 429548 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4669
timestamp 1676037725
transform 1 0 430652 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4675
timestamp 1676037725
transform 1 0 431204 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4677
timestamp 1676037725
transform 1 0 431388 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4689
timestamp 1676037725
transform 1 0 432492 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4701
timestamp 1676037725
transform 1 0 433596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4713
timestamp 1676037725
transform 1 0 434700 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4725
timestamp 1676037725
transform 1 0 435804 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4731
timestamp 1676037725
transform 1 0 436356 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4733
timestamp 1676037725
transform 1 0 436540 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4745
timestamp 1676037725
transform 1 0 437644 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4757
timestamp 1676037725
transform 1 0 438748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4769
timestamp 1676037725
transform 1 0 439852 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4781
timestamp 1676037725
transform 1 0 440956 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4787
timestamp 1676037725
transform 1 0 441508 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4789
timestamp 1676037725
transform 1 0 441692 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4801
timestamp 1676037725
transform 1 0 442796 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4813
timestamp 1676037725
transform 1 0 443900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4825
timestamp 1676037725
transform 1 0 445004 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4837
timestamp 1676037725
transform 1 0 446108 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4843
timestamp 1676037725
transform 1 0 446660 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4845
timestamp 1676037725
transform 1 0 446844 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4857
timestamp 1676037725
transform 1 0 447948 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4869
timestamp 1676037725
transform 1 0 449052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4881
timestamp 1676037725
transform 1 0 450156 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4893
timestamp 1676037725
transform 1 0 451260 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4899
timestamp 1676037725
transform 1 0 451812 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4901
timestamp 1676037725
transform 1 0 451996 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4913
timestamp 1676037725
transform 1 0 453100 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4925
timestamp 1676037725
transform 1 0 454204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4937
timestamp 1676037725
transform 1 0 455308 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4949
timestamp 1676037725
transform 1 0 456412 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4955
timestamp 1676037725
transform 1 0 456964 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4957
timestamp 1676037725
transform 1 0 457148 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4969
timestamp 1676037725
transform 1 0 458252 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4981
timestamp 1676037725
transform 1 0 459356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4993
timestamp 1676037725
transform 1 0 460460 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5005
timestamp 1676037725
transform 1 0 461564 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5011
timestamp 1676037725
transform 1 0 462116 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5013
timestamp 1676037725
transform 1 0 462300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5025
timestamp 1676037725
transform 1 0 463404 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5037
timestamp 1676037725
transform 1 0 464508 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5049
timestamp 1676037725
transform 1 0 465612 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5061
timestamp 1676037725
transform 1 0 466716 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5067
timestamp 1676037725
transform 1 0 467268 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5069
timestamp 1676037725
transform 1 0 467452 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5081
timestamp 1676037725
transform 1 0 468556 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5093
timestamp 1676037725
transform 1 0 469660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5105
timestamp 1676037725
transform 1 0 470764 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5117
timestamp 1676037725
transform 1 0 471868 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5123
timestamp 1676037725
transform 1 0 472420 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5125
timestamp 1676037725
transform 1 0 472604 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5137
timestamp 1676037725
transform 1 0 473708 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5149
timestamp 1676037725
transform 1 0 474812 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5161
timestamp 1676037725
transform 1 0 475916 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5173
timestamp 1676037725
transform 1 0 477020 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5179
timestamp 1676037725
transform 1 0 477572 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5181
timestamp 1676037725
transform 1 0 477756 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5193
timestamp 1676037725
transform 1 0 478860 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5205
timestamp 1676037725
transform 1 0 479964 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5217
timestamp 1676037725
transform 1 0 481068 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5229
timestamp 1676037725
transform 1 0 482172 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5235
timestamp 1676037725
transform 1 0 482724 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5237
timestamp 1676037725
transform 1 0 482908 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5249
timestamp 1676037725
transform 1 0 484012 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5261
timestamp 1676037725
transform 1 0 485116 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5273
timestamp 1676037725
transform 1 0 486220 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5285
timestamp 1676037725
transform 1 0 487324 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5291
timestamp 1676037725
transform 1 0 487876 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5293
timestamp 1676037725
transform 1 0 488060 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5305
timestamp 1676037725
transform 1 0 489164 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5317
timestamp 1676037725
transform 1 0 490268 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5329
timestamp 1676037725
transform 1 0 491372 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5341
timestamp 1676037725
transform 1 0 492476 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5347
timestamp 1676037725
transform 1 0 493028 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5349
timestamp 1676037725
transform 1 0 493212 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5361
timestamp 1676037725
transform 1 0 494316 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5373
timestamp 1676037725
transform 1 0 495420 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5385
timestamp 1676037725
transform 1 0 496524 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5397
timestamp 1676037725
transform 1 0 497628 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5403
timestamp 1676037725
transform 1 0 498180 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_5405
timestamp 1676037725
transform 1 0 498364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_5416
timestamp 1676037725
transform 1 0 499376 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5422
timestamp 1676037725
transform 1 0 499928 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5434
timestamp 1676037725
transform 1 0 501032 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5446
timestamp 1676037725
transform 1 0 502136 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_5458
timestamp 1676037725
transform 1 0 503240 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5461
timestamp 1676037725
transform 1 0 503516 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5473
timestamp 1676037725
transform 1 0 504620 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5485
timestamp 1676037725
transform 1 0 505724 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5497
timestamp 1676037725
transform 1 0 506828 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5509
timestamp 1676037725
transform 1 0 507932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5515
timestamp 1676037725
transform 1 0 508484 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5517
timestamp 1676037725
transform 1 0 508668 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5529
timestamp 1676037725
transform 1 0 509772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5541
timestamp 1676037725
transform 1 0 510876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5553
timestamp 1676037725
transform 1 0 511980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5565
timestamp 1676037725
transform 1 0 513084 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5571
timestamp 1676037725
transform 1 0 513636 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5573
timestamp 1676037725
transform 1 0 513820 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5585
timestamp 1676037725
transform 1 0 514924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5597
timestamp 1676037725
transform 1 0 516028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5609
timestamp 1676037725
transform 1 0 517132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5621
timestamp 1676037725
transform 1 0 518236 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5627
timestamp 1676037725
transform 1 0 518788 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5629
timestamp 1676037725
transform 1 0 518972 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5641
timestamp 1676037725
transform 1 0 520076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5653
timestamp 1676037725
transform 1 0 521180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5665
timestamp 1676037725
transform 1 0 522284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5677
timestamp 1676037725
transform 1 0 523388 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5683
timestamp 1676037725
transform 1 0 523940 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5685
timestamp 1676037725
transform 1 0 524124 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5697
timestamp 1676037725
transform 1 0 525228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5709
timestamp 1676037725
transform 1 0 526332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5721
timestamp 1676037725
transform 1 0 527436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5733
timestamp 1676037725
transform 1 0 528540 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5739
timestamp 1676037725
transform 1 0 529092 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5741
timestamp 1676037725
transform 1 0 529276 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5753
timestamp 1676037725
transform 1 0 530380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5765
timestamp 1676037725
transform 1 0 531484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5777
timestamp 1676037725
transform 1 0 532588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5789
timestamp 1676037725
transform 1 0 533692 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5795
timestamp 1676037725
transform 1 0 534244 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5797
timestamp 1676037725
transform 1 0 534428 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5809
timestamp 1676037725
transform 1 0 535532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5821
timestamp 1676037725
transform 1 0 536636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5833
timestamp 1676037725
transform 1 0 537740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5845
timestamp 1676037725
transform 1 0 538844 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5851
timestamp 1676037725
transform 1 0 539396 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5853
timestamp 1676037725
transform 1 0 539580 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5865
timestamp 1676037725
transform 1 0 540684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5871
timestamp 1676037725
transform 1 0 541236 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_5874
timestamp 1676037725
transform 1 0 541512 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5894
timestamp 1676037725
transform 1 0 543352 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_5906
timestamp 1676037725
transform 1 0 544456 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5909
timestamp 1676037725
transform 1 0 544732 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5921
timestamp 1676037725
transform 1 0 545836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5933
timestamp 1676037725
transform 1 0 546940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5945
timestamp 1676037725
transform 1 0 548044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5957
timestamp 1676037725
transform 1 0 549148 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5963
timestamp 1676037725
transform 1 0 549700 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5965
timestamp 1676037725
transform 1 0 549884 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5977
timestamp 1676037725
transform 1 0 550988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5989
timestamp 1676037725
transform 1 0 552092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6001
timestamp 1676037725
transform 1 0 553196 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6013
timestamp 1676037725
transform 1 0 554300 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6019
timestamp 1676037725
transform 1 0 554852 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6021
timestamp 1676037725
transform 1 0 555036 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6033
timestamp 1676037725
transform 1 0 556140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6045
timestamp 1676037725
transform 1 0 557244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6057
timestamp 1676037725
transform 1 0 558348 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6069
timestamp 1676037725
transform 1 0 559452 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6075
timestamp 1676037725
transform 1 0 560004 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6077
timestamp 1676037725
transform 1 0 560188 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6089
timestamp 1676037725
transform 1 0 561292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6101
timestamp 1676037725
transform 1 0 562396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6113
timestamp 1676037725
transform 1 0 563500 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6125
timestamp 1676037725
transform 1 0 564604 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6131
timestamp 1676037725
transform 1 0 565156 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6133
timestamp 1676037725
transform 1 0 565340 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6145
timestamp 1676037725
transform 1 0 566444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6157
timestamp 1676037725
transform 1 0 567548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6169
timestamp 1676037725
transform 1 0 568652 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6181
timestamp 1676037725
transform 1 0 569756 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6187
timestamp 1676037725
transform 1 0 570308 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6189
timestamp 1676037725
transform 1 0 570492 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6201
timestamp 1676037725
transform 1 0 571596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6213
timestamp 1676037725
transform 1 0 572700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6225
timestamp 1676037725
transform 1 0 573804 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6237
timestamp 1676037725
transform 1 0 574908 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6243
timestamp 1676037725
transform 1 0 575460 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6245
timestamp 1676037725
transform 1 0 575644 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6257
timestamp 1676037725
transform 1 0 576748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6269
timestamp 1676037725
transform 1 0 577852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6281
timestamp 1676037725
transform 1 0 578956 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6293
timestamp 1676037725
transform 1 0 580060 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6299
timestamp 1676037725
transform 1 0 580612 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6301
timestamp 1676037725
transform 1 0 580796 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6313
timestamp 1676037725
transform 1 0 581900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6325
timestamp 1676037725
transform 1 0 583004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6337
timestamp 1676037725
transform 1 0 584108 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6349
timestamp 1676037725
transform 1 0 585212 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6355
timestamp 1676037725
transform 1 0 585764 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6357
timestamp 1676037725
transform 1 0 585948 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6369
timestamp 1676037725
transform 1 0 587052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6381
timestamp 1676037725
transform 1 0 588156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6393
timestamp 1676037725
transform 1 0 589260 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6405
timestamp 1676037725
transform 1 0 590364 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6411
timestamp 1676037725
transform 1 0 590916 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6413
timestamp 1676037725
transform 1 0 591100 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6425
timestamp 1676037725
transform 1 0 592204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6437
timestamp 1676037725
transform 1 0 593308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6449
timestamp 1676037725
transform 1 0 594412 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6461
timestamp 1676037725
transform 1 0 595516 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6467
timestamp 1676037725
transform 1 0 596068 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6469
timestamp 1676037725
transform 1 0 596252 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6481
timestamp 1676037725
transform 1 0 597356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6493
timestamp 1676037725
transform 1 0 598460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6505
timestamp 1676037725
transform 1 0 599564 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6517
timestamp 1676037725
transform 1 0 600668 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6523
timestamp 1676037725
transform 1 0 601220 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6525
timestamp 1676037725
transform 1 0 601404 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6537
timestamp 1676037725
transform 1 0 602508 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6549
timestamp 1676037725
transform 1 0 603612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6561
timestamp 1676037725
transform 1 0 604716 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6573
timestamp 1676037725
transform 1 0 605820 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6579
timestamp 1676037725
transform 1 0 606372 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6581
timestamp 1676037725
transform 1 0 606556 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6593
timestamp 1676037725
transform 1 0 607660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6605
timestamp 1676037725
transform 1 0 608764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6617
timestamp 1676037725
transform 1 0 609868 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6629
timestamp 1676037725
transform 1 0 610972 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6635
timestamp 1676037725
transform 1 0 611524 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6637
timestamp 1676037725
transform 1 0 611708 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6649
timestamp 1676037725
transform 1 0 612812 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6661
timestamp 1676037725
transform 1 0 613916 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6673
timestamp 1676037725
transform 1 0 615020 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6685
timestamp 1676037725
transform 1 0 616124 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6691
timestamp 1676037725
transform 1 0 616676 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6693
timestamp 1676037725
transform 1 0 616860 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6705
timestamp 1676037725
transform 1 0 617964 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6717
timestamp 1676037725
transform 1 0 619068 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6729
timestamp 1676037725
transform 1 0 620172 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6741
timestamp 1676037725
transform 1 0 621276 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6747
timestamp 1676037725
transform 1 0 621828 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6749
timestamp 1676037725
transform 1 0 622012 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6761
timestamp 1676037725
transform 1 0 623116 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6773
timestamp 1676037725
transform 1 0 624220 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6785
timestamp 1676037725
transform 1 0 625324 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6797
timestamp 1676037725
transform 1 0 626428 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6803
timestamp 1676037725
transform 1 0 626980 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6805
timestamp 1676037725
transform 1 0 627164 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6817
timestamp 1676037725
transform 1 0 628268 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6829
timestamp 1676037725
transform 1 0 629372 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6841
timestamp 1676037725
transform 1 0 630476 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6853
timestamp 1676037725
transform 1 0 631580 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6859
timestamp 1676037725
transform 1 0 632132 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6861
timestamp 1676037725
transform 1 0 632316 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6873
timestamp 1676037725
transform 1 0 633420 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6885
timestamp 1676037725
transform 1 0 634524 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6897
timestamp 1676037725
transform 1 0 635628 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6909
timestamp 1676037725
transform 1 0 636732 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6915
timestamp 1676037725
transform 1 0 637284 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6917
timestamp 1676037725
transform 1 0 637468 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6929
timestamp 1676037725
transform 1 0 638572 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6941
timestamp 1676037725
transform 1 0 639676 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6953
timestamp 1676037725
transform 1 0 640780 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6965
timestamp 1676037725
transform 1 0 641884 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6971
timestamp 1676037725
transform 1 0 642436 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6973
timestamp 1676037725
transform 1 0 642620 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6985
timestamp 1676037725
transform 1 0 643724 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6997
timestamp 1676037725
transform 1 0 644828 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7009
timestamp 1676037725
transform 1 0 645932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_7021
timestamp 1676037725
transform 1 0 647036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7027
timestamp 1676037725
transform 1 0 647588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_7029
timestamp 1676037725
transform 1 0 647772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7037
timestamp 1676037725
transform 1 0 648508 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1676037725
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1676037725
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1676037725
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1676037725
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1676037725
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1676037725
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1676037725
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1676037725
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1676037725
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1676037725
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1676037725
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1676037725
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1676037725
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1676037725
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1676037725
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1676037725
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1676037725
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1676037725
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1676037725
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1676037725
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1676037725
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1676037725
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1676037725
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1676037725
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1676037725
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1676037725
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1676037725
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1676037725
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1676037725
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1676037725
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1676037725
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1676037725
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 1676037725
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 1676037725
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1676037725
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1676037725
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1676037725
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_821
timestamp 1676037725
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 1676037725
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 1676037725
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_841
timestamp 1676037725
transform 1 0 78476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_853
timestamp 1676037725
transform 1 0 79580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_865
timestamp 1676037725
transform 1 0 80684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_877
timestamp 1676037725
transform 1 0 81788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_889
timestamp 1676037725
transform 1 0 82892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_895
timestamp 1676037725
transform 1 0 83444 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_897
timestamp 1676037725
transform 1 0 83628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_909
timestamp 1676037725
transform 1 0 84732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_921
timestamp 1676037725
transform 1 0 85836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_933
timestamp 1676037725
transform 1 0 86940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_945
timestamp 1676037725
transform 1 0 88044 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_951
timestamp 1676037725
transform 1 0 88596 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_953
timestamp 1676037725
transform 1 0 88780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_965
timestamp 1676037725
transform 1 0 89884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_977
timestamp 1676037725
transform 1 0 90988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_989
timestamp 1676037725
transform 1 0 92092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1001
timestamp 1676037725
transform 1 0 93196 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1007
timestamp 1676037725
transform 1 0 93748 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1009
timestamp 1676037725
transform 1 0 93932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1021
timestamp 1676037725
transform 1 0 95036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1033
timestamp 1676037725
transform 1 0 96140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1045
timestamp 1676037725
transform 1 0 97244 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1057
timestamp 1676037725
transform 1 0 98348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1063
timestamp 1676037725
transform 1 0 98900 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1065
timestamp 1676037725
transform 1 0 99084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1077
timestamp 1676037725
transform 1 0 100188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1089
timestamp 1676037725
transform 1 0 101292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1101
timestamp 1676037725
transform 1 0 102396 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1113
timestamp 1676037725
transform 1 0 103500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1119
timestamp 1676037725
transform 1 0 104052 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1121
timestamp 1676037725
transform 1 0 104236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1133
timestamp 1676037725
transform 1 0 105340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1145
timestamp 1676037725
transform 1 0 106444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1157
timestamp 1676037725
transform 1 0 107548 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1169
timestamp 1676037725
transform 1 0 108652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1175
timestamp 1676037725
transform 1 0 109204 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1177
timestamp 1676037725
transform 1 0 109388 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1189
timestamp 1676037725
transform 1 0 110492 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1201
timestamp 1676037725
transform 1 0 111596 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1213
timestamp 1676037725
transform 1 0 112700 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1225
timestamp 1676037725
transform 1 0 113804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1231
timestamp 1676037725
transform 1 0 114356 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1233
timestamp 1676037725
transform 1 0 114540 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1245
timestamp 1676037725
transform 1 0 115644 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1257
timestamp 1676037725
transform 1 0 116748 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1269
timestamp 1676037725
transform 1 0 117852 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1281
timestamp 1676037725
transform 1 0 118956 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1287
timestamp 1676037725
transform 1 0 119508 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1289
timestamp 1676037725
transform 1 0 119692 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1301
timestamp 1676037725
transform 1 0 120796 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1313
timestamp 1676037725
transform 1 0 121900 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1325
timestamp 1676037725
transform 1 0 123004 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1337
timestamp 1676037725
transform 1 0 124108 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1343
timestamp 1676037725
transform 1 0 124660 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1345
timestamp 1676037725
transform 1 0 124844 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1357
timestamp 1676037725
transform 1 0 125948 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1369
timestamp 1676037725
transform 1 0 127052 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1381
timestamp 1676037725
transform 1 0 128156 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1393
timestamp 1676037725
transform 1 0 129260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1399
timestamp 1676037725
transform 1 0 129812 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1401
timestamp 1676037725
transform 1 0 129996 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1413
timestamp 1676037725
transform 1 0 131100 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1425
timestamp 1676037725
transform 1 0 132204 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1437
timestamp 1676037725
transform 1 0 133308 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1449
timestamp 1676037725
transform 1 0 134412 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1455
timestamp 1676037725
transform 1 0 134964 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1457
timestamp 1676037725
transform 1 0 135148 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1469
timestamp 1676037725
transform 1 0 136252 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1481
timestamp 1676037725
transform 1 0 137356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1493
timestamp 1676037725
transform 1 0 138460 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1505
timestamp 1676037725
transform 1 0 139564 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1511
timestamp 1676037725
transform 1 0 140116 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1513
timestamp 1676037725
transform 1 0 140300 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1525
timestamp 1676037725
transform 1 0 141404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1537
timestamp 1676037725
transform 1 0 142508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1549
timestamp 1676037725
transform 1 0 143612 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1561
timestamp 1676037725
transform 1 0 144716 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1567
timestamp 1676037725
transform 1 0 145268 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1569
timestamp 1676037725
transform 1 0 145452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1581
timestamp 1676037725
transform 1 0 146556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1593
timestamp 1676037725
transform 1 0 147660 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1605
timestamp 1676037725
transform 1 0 148764 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1617
timestamp 1676037725
transform 1 0 149868 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1623
timestamp 1676037725
transform 1 0 150420 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1625
timestamp 1676037725
transform 1 0 150604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1637
timestamp 1676037725
transform 1 0 151708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1649
timestamp 1676037725
transform 1 0 152812 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1661
timestamp 1676037725
transform 1 0 153916 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1673
timestamp 1676037725
transform 1 0 155020 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1679
timestamp 1676037725
transform 1 0 155572 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1681
timestamp 1676037725
transform 1 0 155756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1693
timestamp 1676037725
transform 1 0 156860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1705
timestamp 1676037725
transform 1 0 157964 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1717
timestamp 1676037725
transform 1 0 159068 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1729
timestamp 1676037725
transform 1 0 160172 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1735
timestamp 1676037725
transform 1 0 160724 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1737
timestamp 1676037725
transform 1 0 160908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1749
timestamp 1676037725
transform 1 0 162012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1761
timestamp 1676037725
transform 1 0 163116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1773
timestamp 1676037725
transform 1 0 164220 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1785
timestamp 1676037725
transform 1 0 165324 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1791
timestamp 1676037725
transform 1 0 165876 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1793
timestamp 1676037725
transform 1 0 166060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1805
timestamp 1676037725
transform 1 0 167164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1817
timestamp 1676037725
transform 1 0 168268 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1829
timestamp 1676037725
transform 1 0 169372 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1841
timestamp 1676037725
transform 1 0 170476 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1847
timestamp 1676037725
transform 1 0 171028 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1849
timestamp 1676037725
transform 1 0 171212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1861
timestamp 1676037725
transform 1 0 172316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1873
timestamp 1676037725
transform 1 0 173420 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1885
timestamp 1676037725
transform 1 0 174524 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1897
timestamp 1676037725
transform 1 0 175628 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1903
timestamp 1676037725
transform 1 0 176180 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1905
timestamp 1676037725
transform 1 0 176364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1917
timestamp 1676037725
transform 1 0 177468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1929
timestamp 1676037725
transform 1 0 178572 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1941
timestamp 1676037725
transform 1 0 179676 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1953
timestamp 1676037725
transform 1 0 180780 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1959
timestamp 1676037725
transform 1 0 181332 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1961
timestamp 1676037725
transform 1 0 181516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1973
timestamp 1676037725
transform 1 0 182620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1985
timestamp 1676037725
transform 1 0 183724 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1997
timestamp 1676037725
transform 1 0 184828 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2009
timestamp 1676037725
transform 1 0 185932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2015
timestamp 1676037725
transform 1 0 186484 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2017
timestamp 1676037725
transform 1 0 186668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2029
timestamp 1676037725
transform 1 0 187772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2041
timestamp 1676037725
transform 1 0 188876 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2053
timestamp 1676037725
transform 1 0 189980 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2065
timestamp 1676037725
transform 1 0 191084 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2071
timestamp 1676037725
transform 1 0 191636 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2073
timestamp 1676037725
transform 1 0 191820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2085
timestamp 1676037725
transform 1 0 192924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2097
timestamp 1676037725
transform 1 0 194028 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2109
timestamp 1676037725
transform 1 0 195132 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2121
timestamp 1676037725
transform 1 0 196236 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2127
timestamp 1676037725
transform 1 0 196788 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2129
timestamp 1676037725
transform 1 0 196972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2141
timestamp 1676037725
transform 1 0 198076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2153
timestamp 1676037725
transform 1 0 199180 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2165
timestamp 1676037725
transform 1 0 200284 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2177
timestamp 1676037725
transform 1 0 201388 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2183
timestamp 1676037725
transform 1 0 201940 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2185
timestamp 1676037725
transform 1 0 202124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2197
timestamp 1676037725
transform 1 0 203228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2209
timestamp 1676037725
transform 1 0 204332 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2221
timestamp 1676037725
transform 1 0 205436 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2233
timestamp 1676037725
transform 1 0 206540 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2239
timestamp 1676037725
transform 1 0 207092 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2241
timestamp 1676037725
transform 1 0 207276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2253
timestamp 1676037725
transform 1 0 208380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2265
timestamp 1676037725
transform 1 0 209484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2277
timestamp 1676037725
transform 1 0 210588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2289
timestamp 1676037725
transform 1 0 211692 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2295
timestamp 1676037725
transform 1 0 212244 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2297
timestamp 1676037725
transform 1 0 212428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2309
timestamp 1676037725
transform 1 0 213532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2321
timestamp 1676037725
transform 1 0 214636 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2333
timestamp 1676037725
transform 1 0 215740 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2345
timestamp 1676037725
transform 1 0 216844 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2351
timestamp 1676037725
transform 1 0 217396 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2353
timestamp 1676037725
transform 1 0 217580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2365
timestamp 1676037725
transform 1 0 218684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2377
timestamp 1676037725
transform 1 0 219788 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2389
timestamp 1676037725
transform 1 0 220892 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2401
timestamp 1676037725
transform 1 0 221996 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2407
timestamp 1676037725
transform 1 0 222548 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2409
timestamp 1676037725
transform 1 0 222732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2421
timestamp 1676037725
transform 1 0 223836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2433
timestamp 1676037725
transform 1 0 224940 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2445
timestamp 1676037725
transform 1 0 226044 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2457
timestamp 1676037725
transform 1 0 227148 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2463
timestamp 1676037725
transform 1 0 227700 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2465
timestamp 1676037725
transform 1 0 227884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2477
timestamp 1676037725
transform 1 0 228988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2489
timestamp 1676037725
transform 1 0 230092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2501
timestamp 1676037725
transform 1 0 231196 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2513
timestamp 1676037725
transform 1 0 232300 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2519
timestamp 1676037725
transform 1 0 232852 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2521
timestamp 1676037725
transform 1 0 233036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2533
timestamp 1676037725
transform 1 0 234140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2545
timestamp 1676037725
transform 1 0 235244 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2557
timestamp 1676037725
transform 1 0 236348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2569
timestamp 1676037725
transform 1 0 237452 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2575
timestamp 1676037725
transform 1 0 238004 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2577
timestamp 1676037725
transform 1 0 238188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2589
timestamp 1676037725
transform 1 0 239292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2601
timestamp 1676037725
transform 1 0 240396 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2613
timestamp 1676037725
transform 1 0 241500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2625
timestamp 1676037725
transform 1 0 242604 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2631
timestamp 1676037725
transform 1 0 243156 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2633
timestamp 1676037725
transform 1 0 243340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2645
timestamp 1676037725
transform 1 0 244444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2657
timestamp 1676037725
transform 1 0 245548 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2669
timestamp 1676037725
transform 1 0 246652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2681
timestamp 1676037725
transform 1 0 247756 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2687
timestamp 1676037725
transform 1 0 248308 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2689
timestamp 1676037725
transform 1 0 248492 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2701
timestamp 1676037725
transform 1 0 249596 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2713
timestamp 1676037725
transform 1 0 250700 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2725
timestamp 1676037725
transform 1 0 251804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2737
timestamp 1676037725
transform 1 0 252908 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2743
timestamp 1676037725
transform 1 0 253460 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2745
timestamp 1676037725
transform 1 0 253644 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2757
timestamp 1676037725
transform 1 0 254748 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2769
timestamp 1676037725
transform 1 0 255852 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2781
timestamp 1676037725
transform 1 0 256956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2793
timestamp 1676037725
transform 1 0 258060 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2799
timestamp 1676037725
transform 1 0 258612 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2801
timestamp 1676037725
transform 1 0 258796 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2813
timestamp 1676037725
transform 1 0 259900 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2825
timestamp 1676037725
transform 1 0 261004 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2837
timestamp 1676037725
transform 1 0 262108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2849
timestamp 1676037725
transform 1 0 263212 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2855
timestamp 1676037725
transform 1 0 263764 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2857
timestamp 1676037725
transform 1 0 263948 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2869
timestamp 1676037725
transform 1 0 265052 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2881
timestamp 1676037725
transform 1 0 266156 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2893
timestamp 1676037725
transform 1 0 267260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2905
timestamp 1676037725
transform 1 0 268364 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2911
timestamp 1676037725
transform 1 0 268916 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2913
timestamp 1676037725
transform 1 0 269100 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2925
timestamp 1676037725
transform 1 0 270204 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2937
timestamp 1676037725
transform 1 0 271308 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2949
timestamp 1676037725
transform 1 0 272412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2961
timestamp 1676037725
transform 1 0 273516 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2967
timestamp 1676037725
transform 1 0 274068 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2969
timestamp 1676037725
transform 1 0 274252 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2981
timestamp 1676037725
transform 1 0 275356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2993
timestamp 1676037725
transform 1 0 276460 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3005
timestamp 1676037725
transform 1 0 277564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3017
timestamp 1676037725
transform 1 0 278668 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3023
timestamp 1676037725
transform 1 0 279220 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3025
timestamp 1676037725
transform 1 0 279404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3037
timestamp 1676037725
transform 1 0 280508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3049
timestamp 1676037725
transform 1 0 281612 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3061
timestamp 1676037725
transform 1 0 282716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3073
timestamp 1676037725
transform 1 0 283820 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3079
timestamp 1676037725
transform 1 0 284372 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3081
timestamp 1676037725
transform 1 0 284556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3093
timestamp 1676037725
transform 1 0 285660 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3105
timestamp 1676037725
transform 1 0 286764 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3117
timestamp 1676037725
transform 1 0 287868 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3129
timestamp 1676037725
transform 1 0 288972 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3135
timestamp 1676037725
transform 1 0 289524 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3137
timestamp 1676037725
transform 1 0 289708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3149
timestamp 1676037725
transform 1 0 290812 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3161
timestamp 1676037725
transform 1 0 291916 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3173
timestamp 1676037725
transform 1 0 293020 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3185
timestamp 1676037725
transform 1 0 294124 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3191
timestamp 1676037725
transform 1 0 294676 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3193
timestamp 1676037725
transform 1 0 294860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3205
timestamp 1676037725
transform 1 0 295964 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3217
timestamp 1676037725
transform 1 0 297068 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3229
timestamp 1676037725
transform 1 0 298172 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3241
timestamp 1676037725
transform 1 0 299276 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3247
timestamp 1676037725
transform 1 0 299828 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3249
timestamp 1676037725
transform 1 0 300012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3261
timestamp 1676037725
transform 1 0 301116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3273
timestamp 1676037725
transform 1 0 302220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3285
timestamp 1676037725
transform 1 0 303324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3297
timestamp 1676037725
transform 1 0 304428 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3303
timestamp 1676037725
transform 1 0 304980 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3305
timestamp 1676037725
transform 1 0 305164 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3311
timestamp 1676037725
transform 1 0 305716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3321
timestamp 1676037725
transform 1 0 306636 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3327
timestamp 1676037725
transform 1 0 307188 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3339
timestamp 1676037725
transform 1 0 308292 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3343
timestamp 1676037725
transform 1 0 308660 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3346
timestamp 1676037725
transform 1 0 308936 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3352
timestamp 1676037725
transform 1 0 309488 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3361
timestamp 1676037725
transform 1 0 310316 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3365
timestamp 1676037725
transform 1 0 310684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3368
timestamp 1676037725
transform 1 0 310960 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3380
timestamp 1676037725
transform 1 0 312064 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3392
timestamp 1676037725
transform 1 0 313168 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3404
timestamp 1676037725
transform 1 0 314272 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3417
timestamp 1676037725
transform 1 0 315468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3429
timestamp 1676037725
transform 1 0 316572 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3441
timestamp 1676037725
transform 1 0 317676 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3453
timestamp 1676037725
transform 1 0 318780 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3465
timestamp 1676037725
transform 1 0 319884 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3471
timestamp 1676037725
transform 1 0 320436 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3473
timestamp 1676037725
transform 1 0 320620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3485
timestamp 1676037725
transform 1 0 321724 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3497
timestamp 1676037725
transform 1 0 322828 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3509
timestamp 1676037725
transform 1 0 323932 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3521
timestamp 1676037725
transform 1 0 325036 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3527
timestamp 1676037725
transform 1 0 325588 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3529
timestamp 1676037725
transform 1 0 325772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3541
timestamp 1676037725
transform 1 0 326876 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3553
timestamp 1676037725
transform 1 0 327980 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3565
timestamp 1676037725
transform 1 0 329084 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3577
timestamp 1676037725
transform 1 0 330188 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3583
timestamp 1676037725
transform 1 0 330740 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3585
timestamp 1676037725
transform 1 0 330924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3597
timestamp 1676037725
transform 1 0 332028 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3609
timestamp 1676037725
transform 1 0 333132 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3621
timestamp 1676037725
transform 1 0 334236 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3633
timestamp 1676037725
transform 1 0 335340 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3639
timestamp 1676037725
transform 1 0 335892 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3641
timestamp 1676037725
transform 1 0 336076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3653
timestamp 1676037725
transform 1 0 337180 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3665
timestamp 1676037725
transform 1 0 338284 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3677
timestamp 1676037725
transform 1 0 339388 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3689
timestamp 1676037725
transform 1 0 340492 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3695
timestamp 1676037725
transform 1 0 341044 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3697
timestamp 1676037725
transform 1 0 341228 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3716
timestamp 1676037725
transform 1 0 342976 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3728
timestamp 1676037725
transform 1 0 344080 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3740
timestamp 1676037725
transform 1 0 345184 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3753
timestamp 1676037725
transform 1 0 346380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3765
timestamp 1676037725
transform 1 0 347484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3777
timestamp 1676037725
transform 1 0 348588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3789
timestamp 1676037725
transform 1 0 349692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3801
timestamp 1676037725
transform 1 0 350796 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3807
timestamp 1676037725
transform 1 0 351348 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3809
timestamp 1676037725
transform 1 0 351532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3821
timestamp 1676037725
transform 1 0 352636 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3833
timestamp 1676037725
transform 1 0 353740 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3845
timestamp 1676037725
transform 1 0 354844 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3857
timestamp 1676037725
transform 1 0 355948 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3862
timestamp 1676037725
transform 1 0 356408 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3865
timestamp 1676037725
transform 1 0 356684 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3883
timestamp 1676037725
transform 1 0 358340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3895
timestamp 1676037725
transform 1 0 359444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3907
timestamp 1676037725
transform 1 0 360548 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3919
timestamp 1676037725
transform 1 0 361652 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3921
timestamp 1676037725
transform 1 0 361836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3933
timestamp 1676037725
transform 1 0 362940 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3945
timestamp 1676037725
transform 1 0 364044 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3957
timestamp 1676037725
transform 1 0 365148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3969
timestamp 1676037725
transform 1 0 366252 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3975
timestamp 1676037725
transform 1 0 366804 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3977
timestamp 1676037725
transform 1 0 366988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3989
timestamp 1676037725
transform 1 0 368092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4001
timestamp 1676037725
transform 1 0 369196 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4013
timestamp 1676037725
transform 1 0 370300 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4025
timestamp 1676037725
transform 1 0 371404 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4031
timestamp 1676037725
transform 1 0 371956 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4033
timestamp 1676037725
transform 1 0 372140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4045
timestamp 1676037725
transform 1 0 373244 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4057
timestamp 1676037725
transform 1 0 374348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4069
timestamp 1676037725
transform 1 0 375452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4081
timestamp 1676037725
transform 1 0 376556 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4087
timestamp 1676037725
transform 1 0 377108 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4089
timestamp 1676037725
transform 1 0 377292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4101
timestamp 1676037725
transform 1 0 378396 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4113
timestamp 1676037725
transform 1 0 379500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4125
timestamp 1676037725
transform 1 0 380604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4137
timestamp 1676037725
transform 1 0 381708 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4143
timestamp 1676037725
transform 1 0 382260 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4145
timestamp 1676037725
transform 1 0 382444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4157
timestamp 1676037725
transform 1 0 383548 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4169
timestamp 1676037725
transform 1 0 384652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4181
timestamp 1676037725
transform 1 0 385756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_4193
timestamp 1676037725
transform 1 0 386860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_4198
timestamp 1676037725
transform 1 0 387320 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_4201
timestamp 1676037725
transform 1 0 387596 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4219
timestamp 1676037725
transform 1 0 389252 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4231
timestamp 1676037725
transform 1 0 390356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4243
timestamp 1676037725
transform 1 0 391460 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4255
timestamp 1676037725
transform 1 0 392564 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4257
timestamp 1676037725
transform 1 0 392748 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4269
timestamp 1676037725
transform 1 0 393852 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4281
timestamp 1676037725
transform 1 0 394956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4293
timestamp 1676037725
transform 1 0 396060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4305
timestamp 1676037725
transform 1 0 397164 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4311
timestamp 1676037725
transform 1 0 397716 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4313
timestamp 1676037725
transform 1 0 397900 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4325
timestamp 1676037725
transform 1 0 399004 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4337
timestamp 1676037725
transform 1 0 400108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4349
timestamp 1676037725
transform 1 0 401212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_4361
timestamp 1676037725
transform 1 0 402316 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_4366
timestamp 1676037725
transform 1 0 402776 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_4369
timestamp 1676037725
transform 1 0 403052 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4387
timestamp 1676037725
transform 1 0 404708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4399
timestamp 1676037725
transform 1 0 405812 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4411
timestamp 1676037725
transform 1 0 406916 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4423
timestamp 1676037725
transform 1 0 408020 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4425
timestamp 1676037725
transform 1 0 408204 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4437
timestamp 1676037725
transform 1 0 409308 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4449
timestamp 1676037725
transform 1 0 410412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4461
timestamp 1676037725
transform 1 0 411516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4473
timestamp 1676037725
transform 1 0 412620 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4479
timestamp 1676037725
transform 1 0 413172 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4481
timestamp 1676037725
transform 1 0 413356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4493
timestamp 1676037725
transform 1 0 414460 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4505
timestamp 1676037725
transform 1 0 415564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4517
timestamp 1676037725
transform 1 0 416668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4529
timestamp 1676037725
transform 1 0 417772 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4535
timestamp 1676037725
transform 1 0 418324 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4537
timestamp 1676037725
transform 1 0 418508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4549
timestamp 1676037725
transform 1 0 419612 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4561
timestamp 1676037725
transform 1 0 420716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4573
timestamp 1676037725
transform 1 0 421820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4585
timestamp 1676037725
transform 1 0 422924 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4591
timestamp 1676037725
transform 1 0 423476 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4593
timestamp 1676037725
transform 1 0 423660 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4605
timestamp 1676037725
transform 1 0 424764 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4617
timestamp 1676037725
transform 1 0 425868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4629
timestamp 1676037725
transform 1 0 426972 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4641
timestamp 1676037725
transform 1 0 428076 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4647
timestamp 1676037725
transform 1 0 428628 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4649
timestamp 1676037725
transform 1 0 428812 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4661
timestamp 1676037725
transform 1 0 429916 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4673
timestamp 1676037725
transform 1 0 431020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4685
timestamp 1676037725
transform 1 0 432124 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_4697
timestamp 1676037725
transform 1 0 433228 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_4702
timestamp 1676037725
transform 1 0 433688 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_4705
timestamp 1676037725
transform 1 0 433964 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4723
timestamp 1676037725
transform 1 0 435620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4735
timestamp 1676037725
transform 1 0 436724 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4747
timestamp 1676037725
transform 1 0 437828 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4759
timestamp 1676037725
transform 1 0 438932 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4761
timestamp 1676037725
transform 1 0 439116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4773
timestamp 1676037725
transform 1 0 440220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4785
timestamp 1676037725
transform 1 0 441324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4797
timestamp 1676037725
transform 1 0 442428 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4809
timestamp 1676037725
transform 1 0 443532 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4815
timestamp 1676037725
transform 1 0 444084 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4817
timestamp 1676037725
transform 1 0 444268 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4829
timestamp 1676037725
transform 1 0 445372 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4841
timestamp 1676037725
transform 1 0 446476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4853
timestamp 1676037725
transform 1 0 447580 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_4865
timestamp 1676037725
transform 1 0 448684 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_4870
timestamp 1676037725
transform 1 0 449144 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_4873
timestamp 1676037725
transform 1 0 449420 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4891
timestamp 1676037725
transform 1 0 451076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4903
timestamp 1676037725
transform 1 0 452180 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4915
timestamp 1676037725
transform 1 0 453284 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4927
timestamp 1676037725
transform 1 0 454388 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4929
timestamp 1676037725
transform 1 0 454572 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4941
timestamp 1676037725
transform 1 0 455676 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4953
timestamp 1676037725
transform 1 0 456780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4965
timestamp 1676037725
transform 1 0 457884 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4977
timestamp 1676037725
transform 1 0 458988 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4983
timestamp 1676037725
transform 1 0 459540 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4985
timestamp 1676037725
transform 1 0 459724 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4997
timestamp 1676037725
transform 1 0 460828 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5009
timestamp 1676037725
transform 1 0 461932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5021
timestamp 1676037725
transform 1 0 463036 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5033
timestamp 1676037725
transform 1 0 464140 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5039
timestamp 1676037725
transform 1 0 464692 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5041
timestamp 1676037725
transform 1 0 464876 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5053
timestamp 1676037725
transform 1 0 465980 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5065
timestamp 1676037725
transform 1 0 467084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5077
timestamp 1676037725
transform 1 0 468188 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5089
timestamp 1676037725
transform 1 0 469292 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5095
timestamp 1676037725
transform 1 0 469844 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5097
timestamp 1676037725
transform 1 0 470028 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5109
timestamp 1676037725
transform 1 0 471132 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5121
timestamp 1676037725
transform 1 0 472236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5133
timestamp 1676037725
transform 1 0 473340 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5145
timestamp 1676037725
transform 1 0 474444 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5151
timestamp 1676037725
transform 1 0 474996 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5153
timestamp 1676037725
transform 1 0 475180 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5165
timestamp 1676037725
transform 1 0 476284 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5177
timestamp 1676037725
transform 1 0 477388 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5189
timestamp 1676037725
transform 1 0 478492 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_5201
timestamp 1676037725
transform 1 0 479596 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_5206
timestamp 1676037725
transform 1 0 480056 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_5209
timestamp 1676037725
transform 1 0 480332 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5227
timestamp 1676037725
transform 1 0 481988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5239
timestamp 1676037725
transform 1 0 483092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5251
timestamp 1676037725
transform 1 0 484196 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5263
timestamp 1676037725
transform 1 0 485300 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5265
timestamp 1676037725
transform 1 0 485484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5277
timestamp 1676037725
transform 1 0 486588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5289
timestamp 1676037725
transform 1 0 487692 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5301
timestamp 1676037725
transform 1 0 488796 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5313
timestamp 1676037725
transform 1 0 489900 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5319
timestamp 1676037725
transform 1 0 490452 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5321
timestamp 1676037725
transform 1 0 490636 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5333
timestamp 1676037725
transform 1 0 491740 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5345
timestamp 1676037725
transform 1 0 492844 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5357
timestamp 1676037725
transform 1 0 493948 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_5369
timestamp 1676037725
transform 1 0 495052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_5374
timestamp 1676037725
transform 1 0 495512 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_5377
timestamp 1676037725
transform 1 0 495788 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5395
timestamp 1676037725
transform 1 0 497444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5407
timestamp 1676037725
transform 1 0 498548 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_5419
timestamp 1676037725
transform 1 0 499652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_5430
timestamp 1676037725
transform 1 0 500664 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_5433
timestamp 1676037725
transform 1 0 500940 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5437
timestamp 1676037725
transform 1 0 501308 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5449
timestamp 1676037725
transform 1 0 502412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5461
timestamp 1676037725
transform 1 0 503516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5473
timestamp 1676037725
transform 1 0 504620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_5485
timestamp 1676037725
transform 1 0 505724 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5489
timestamp 1676037725
transform 1 0 506092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5501
timestamp 1676037725
transform 1 0 507196 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5513
timestamp 1676037725
transform 1 0 508300 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5525
timestamp 1676037725
transform 1 0 509404 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5537
timestamp 1676037725
transform 1 0 510508 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5543
timestamp 1676037725
transform 1 0 511060 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5545
timestamp 1676037725
transform 1 0 511244 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5557
timestamp 1676037725
transform 1 0 512348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5569
timestamp 1676037725
transform 1 0 513452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5581
timestamp 1676037725
transform 1 0 514556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5593
timestamp 1676037725
transform 1 0 515660 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5599
timestamp 1676037725
transform 1 0 516212 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5601
timestamp 1676037725
transform 1 0 516396 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5613
timestamp 1676037725
transform 1 0 517500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5625
timestamp 1676037725
transform 1 0 518604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5637
timestamp 1676037725
transform 1 0 519708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5649
timestamp 1676037725
transform 1 0 520812 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5655
timestamp 1676037725
transform 1 0 521364 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5657
timestamp 1676037725
transform 1 0 521548 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5669
timestamp 1676037725
transform 1 0 522652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5681
timestamp 1676037725
transform 1 0 523756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5693
timestamp 1676037725
transform 1 0 524860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_5705
timestamp 1676037725
transform 1 0 525964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_5710
timestamp 1676037725
transform 1 0 526424 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_5713
timestamp 1676037725
transform 1 0 526700 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5731
timestamp 1676037725
transform 1 0 528356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5743
timestamp 1676037725
transform 1 0 529460 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5755
timestamp 1676037725
transform 1 0 530564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5767
timestamp 1676037725
transform 1 0 531668 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5769
timestamp 1676037725
transform 1 0 531852 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5781
timestamp 1676037725
transform 1 0 532956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5793
timestamp 1676037725
transform 1 0 534060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5805
timestamp 1676037725
transform 1 0 535164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5817
timestamp 1676037725
transform 1 0 536268 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5823
timestamp 1676037725
transform 1 0 536820 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5825
timestamp 1676037725
transform 1 0 537004 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5837
timestamp 1676037725
transform 1 0 538108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5849
timestamp 1676037725
transform 1 0 539212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5861
timestamp 1676037725
transform 1 0 540316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5873
timestamp 1676037725
transform 1 0 541420 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5879
timestamp 1676037725
transform 1 0 541972 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5881
timestamp 1676037725
transform 1 0 542156 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5893
timestamp 1676037725
transform 1 0 543260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5905
timestamp 1676037725
transform 1 0 544364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5917
timestamp 1676037725
transform 1 0 545468 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5929
timestamp 1676037725
transform 1 0 546572 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5935
timestamp 1676037725
transform 1 0 547124 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5937
timestamp 1676037725
transform 1 0 547308 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5949
timestamp 1676037725
transform 1 0 548412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5961
timestamp 1676037725
transform 1 0 549516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5973
timestamp 1676037725
transform 1 0 550620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5985
timestamp 1676037725
transform 1 0 551724 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5991
timestamp 1676037725
transform 1 0 552276 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5993
timestamp 1676037725
transform 1 0 552460 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6005
timestamp 1676037725
transform 1 0 553564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6017
timestamp 1676037725
transform 1 0 554668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6029
timestamp 1676037725
transform 1 0 555772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6041
timestamp 1676037725
transform 1 0 556876 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6047
timestamp 1676037725
transform 1 0 557428 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6049
timestamp 1676037725
transform 1 0 557612 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6061
timestamp 1676037725
transform 1 0 558716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6073
timestamp 1676037725
transform 1 0 559820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6085
timestamp 1676037725
transform 1 0 560924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6097
timestamp 1676037725
transform 1 0 562028 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6103
timestamp 1676037725
transform 1 0 562580 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6105
timestamp 1676037725
transform 1 0 562764 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6117
timestamp 1676037725
transform 1 0 563868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6129
timestamp 1676037725
transform 1 0 564972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6141
timestamp 1676037725
transform 1 0 566076 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6153
timestamp 1676037725
transform 1 0 567180 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6159
timestamp 1676037725
transform 1 0 567732 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6161
timestamp 1676037725
transform 1 0 567916 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6173
timestamp 1676037725
transform 1 0 569020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6185
timestamp 1676037725
transform 1 0 570124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6197
timestamp 1676037725
transform 1 0 571228 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6209
timestamp 1676037725
transform 1 0 572332 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6215
timestamp 1676037725
transform 1 0 572884 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6217
timestamp 1676037725
transform 1 0 573068 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6229
timestamp 1676037725
transform 1 0 574172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6241
timestamp 1676037725
transform 1 0 575276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6253
timestamp 1676037725
transform 1 0 576380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6265
timestamp 1676037725
transform 1 0 577484 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6271
timestamp 1676037725
transform 1 0 578036 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6273
timestamp 1676037725
transform 1 0 578220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6285
timestamp 1676037725
transform 1 0 579324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6297
timestamp 1676037725
transform 1 0 580428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6309
timestamp 1676037725
transform 1 0 581532 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6321
timestamp 1676037725
transform 1 0 582636 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6327
timestamp 1676037725
transform 1 0 583188 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6329
timestamp 1676037725
transform 1 0 583372 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6341
timestamp 1676037725
transform 1 0 584476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6353
timestamp 1676037725
transform 1 0 585580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6365
timestamp 1676037725
transform 1 0 586684 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6377
timestamp 1676037725
transform 1 0 587788 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6383
timestamp 1676037725
transform 1 0 588340 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6385
timestamp 1676037725
transform 1 0 588524 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6397
timestamp 1676037725
transform 1 0 589628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6409
timestamp 1676037725
transform 1 0 590732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6421
timestamp 1676037725
transform 1 0 591836 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6433
timestamp 1676037725
transform 1 0 592940 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6439
timestamp 1676037725
transform 1 0 593492 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6441
timestamp 1676037725
transform 1 0 593676 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6453
timestamp 1676037725
transform 1 0 594780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6465
timestamp 1676037725
transform 1 0 595884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6477
timestamp 1676037725
transform 1 0 596988 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6489
timestamp 1676037725
transform 1 0 598092 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6495
timestamp 1676037725
transform 1 0 598644 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6497
timestamp 1676037725
transform 1 0 598828 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6509
timestamp 1676037725
transform 1 0 599932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6521
timestamp 1676037725
transform 1 0 601036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6533
timestamp 1676037725
transform 1 0 602140 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6545
timestamp 1676037725
transform 1 0 603244 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6551
timestamp 1676037725
transform 1 0 603796 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6553
timestamp 1676037725
transform 1 0 603980 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6565
timestamp 1676037725
transform 1 0 605084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6577
timestamp 1676037725
transform 1 0 606188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6589
timestamp 1676037725
transform 1 0 607292 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6601
timestamp 1676037725
transform 1 0 608396 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6607
timestamp 1676037725
transform 1 0 608948 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6609
timestamp 1676037725
transform 1 0 609132 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6621
timestamp 1676037725
transform 1 0 610236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6633
timestamp 1676037725
transform 1 0 611340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6645
timestamp 1676037725
transform 1 0 612444 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6657
timestamp 1676037725
transform 1 0 613548 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6663
timestamp 1676037725
transform 1 0 614100 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6665
timestamp 1676037725
transform 1 0 614284 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6677
timestamp 1676037725
transform 1 0 615388 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6689
timestamp 1676037725
transform 1 0 616492 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6701
timestamp 1676037725
transform 1 0 617596 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6713
timestamp 1676037725
transform 1 0 618700 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6719
timestamp 1676037725
transform 1 0 619252 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6721
timestamp 1676037725
transform 1 0 619436 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6733
timestamp 1676037725
transform 1 0 620540 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6745
timestamp 1676037725
transform 1 0 621644 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6757
timestamp 1676037725
transform 1 0 622748 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6769
timestamp 1676037725
transform 1 0 623852 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6775
timestamp 1676037725
transform 1 0 624404 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6777
timestamp 1676037725
transform 1 0 624588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6789
timestamp 1676037725
transform 1 0 625692 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6801
timestamp 1676037725
transform 1 0 626796 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6813
timestamp 1676037725
transform 1 0 627900 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6825
timestamp 1676037725
transform 1 0 629004 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6831
timestamp 1676037725
transform 1 0 629556 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6833
timestamp 1676037725
transform 1 0 629740 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6845
timestamp 1676037725
transform 1 0 630844 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6857
timestamp 1676037725
transform 1 0 631948 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6869
timestamp 1676037725
transform 1 0 633052 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6881
timestamp 1676037725
transform 1 0 634156 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6887
timestamp 1676037725
transform 1 0 634708 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6889
timestamp 1676037725
transform 1 0 634892 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6901
timestamp 1676037725
transform 1 0 635996 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6913
timestamp 1676037725
transform 1 0 637100 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6925
timestamp 1676037725
transform 1 0 638204 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6937
timestamp 1676037725
transform 1 0 639308 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6943
timestamp 1676037725
transform 1 0 639860 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6945
timestamp 1676037725
transform 1 0 640044 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6957
timestamp 1676037725
transform 1 0 641148 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6969
timestamp 1676037725
transform 1 0 642252 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6981
timestamp 1676037725
transform 1 0 643356 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6993
timestamp 1676037725
transform 1 0 644460 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6999
timestamp 1676037725
transform 1 0 645012 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7001
timestamp 1676037725
transform 1 0 645196 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7013
timestamp 1676037725
transform 1 0 646300 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7025
timestamp 1676037725
transform 1 0 647404 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7037
timestamp 1676037725
transform 1 0 648508 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1676037725
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1676037725
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1676037725
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1676037725
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1676037725
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1676037725
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1676037725
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1676037725
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1676037725
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1676037725
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1676037725
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1676037725
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1676037725
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1676037725
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1676037725
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1676037725
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1676037725
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1676037725
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1676037725
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1676037725
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1676037725
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1676037725
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1676037725
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1676037725
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1676037725
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1676037725
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1676037725
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1676037725
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1676037725
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1676037725
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1676037725
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1676037725
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1676037725
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1676037725
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1676037725
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1676037725
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1676037725
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1676037725
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_781
timestamp 1676037725
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_793
timestamp 1676037725
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 1676037725
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 1676037725
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1676037725
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_825
timestamp 1676037725
transform 1 0 77004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_837
timestamp 1676037725
transform 1 0 78108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_849
timestamp 1676037725
transform 1 0 79212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_861
timestamp 1676037725
transform 1 0 80316 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_867
timestamp 1676037725
transform 1 0 80868 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_869
timestamp 1676037725
transform 1 0 81052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_881
timestamp 1676037725
transform 1 0 82156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_893
timestamp 1676037725
transform 1 0 83260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_905
timestamp 1676037725
transform 1 0 84364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_917
timestamp 1676037725
transform 1 0 85468 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_923
timestamp 1676037725
transform 1 0 86020 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_925
timestamp 1676037725
transform 1 0 86204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_937
timestamp 1676037725
transform 1 0 87308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_949
timestamp 1676037725
transform 1 0 88412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_961
timestamp 1676037725
transform 1 0 89516 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_973
timestamp 1676037725
transform 1 0 90620 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_979
timestamp 1676037725
transform 1 0 91172 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_981
timestamp 1676037725
transform 1 0 91356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_993
timestamp 1676037725
transform 1 0 92460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1005
timestamp 1676037725
transform 1 0 93564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1017
timestamp 1676037725
transform 1 0 94668 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1029
timestamp 1676037725
transform 1 0 95772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1035
timestamp 1676037725
transform 1 0 96324 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1037
timestamp 1676037725
transform 1 0 96508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1049
timestamp 1676037725
transform 1 0 97612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1061
timestamp 1676037725
transform 1 0 98716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1073
timestamp 1676037725
transform 1 0 99820 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1085
timestamp 1676037725
transform 1 0 100924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1091
timestamp 1676037725
transform 1 0 101476 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1093
timestamp 1676037725
transform 1 0 101660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1105
timestamp 1676037725
transform 1 0 102764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1117
timestamp 1676037725
transform 1 0 103868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1129
timestamp 1676037725
transform 1 0 104972 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1141
timestamp 1676037725
transform 1 0 106076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1147
timestamp 1676037725
transform 1 0 106628 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1149
timestamp 1676037725
transform 1 0 106812 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1161
timestamp 1676037725
transform 1 0 107916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1173
timestamp 1676037725
transform 1 0 109020 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1185
timestamp 1676037725
transform 1 0 110124 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1197
timestamp 1676037725
transform 1 0 111228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1203
timestamp 1676037725
transform 1 0 111780 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1205
timestamp 1676037725
transform 1 0 111964 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1213
timestamp 1676037725
transform 1 0 112700 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1219
timestamp 1676037725
transform 1 0 113252 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1231
timestamp 1676037725
transform 1 0 114356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1243
timestamp 1676037725
transform 1 0 115460 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1255
timestamp 1676037725
transform 1 0 116564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1259
timestamp 1676037725
transform 1 0 116932 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1261
timestamp 1676037725
transform 1 0 117116 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1273
timestamp 1676037725
transform 1 0 118220 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1285
timestamp 1676037725
transform 1 0 119324 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1297
timestamp 1676037725
transform 1 0 120428 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1309
timestamp 1676037725
transform 1 0 121532 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1315
timestamp 1676037725
transform 1 0 122084 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1317
timestamp 1676037725
transform 1 0 122268 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1329
timestamp 1676037725
transform 1 0 123372 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1341
timestamp 1676037725
transform 1 0 124476 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1353
timestamp 1676037725
transform 1 0 125580 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1365
timestamp 1676037725
transform 1 0 126684 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1371
timestamp 1676037725
transform 1 0 127236 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1373
timestamp 1676037725
transform 1 0 127420 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1385
timestamp 1676037725
transform 1 0 128524 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1397
timestamp 1676037725
transform 1 0 129628 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1409
timestamp 1676037725
transform 1 0 130732 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1421
timestamp 1676037725
transform 1 0 131836 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1427
timestamp 1676037725
transform 1 0 132388 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1429
timestamp 1676037725
transform 1 0 132572 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1441
timestamp 1676037725
transform 1 0 133676 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1453
timestamp 1676037725
transform 1 0 134780 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1465
timestamp 1676037725
transform 1 0 135884 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1477
timestamp 1676037725
transform 1 0 136988 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1483
timestamp 1676037725
transform 1 0 137540 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1485
timestamp 1676037725
transform 1 0 137724 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1497
timestamp 1676037725
transform 1 0 138828 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1509
timestamp 1676037725
transform 1 0 139932 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1521
timestamp 1676037725
transform 1 0 141036 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1533
timestamp 1676037725
transform 1 0 142140 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1539
timestamp 1676037725
transform 1 0 142692 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1541
timestamp 1676037725
transform 1 0 142876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1553
timestamp 1676037725
transform 1 0 143980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1565
timestamp 1676037725
transform 1 0 145084 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1577
timestamp 1676037725
transform 1 0 146188 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1589
timestamp 1676037725
transform 1 0 147292 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1595
timestamp 1676037725
transform 1 0 147844 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1597
timestamp 1676037725
transform 1 0 148028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1609
timestamp 1676037725
transform 1 0 149132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1621
timestamp 1676037725
transform 1 0 150236 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1633
timestamp 1676037725
transform 1 0 151340 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1645
timestamp 1676037725
transform 1 0 152444 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1651
timestamp 1676037725
transform 1 0 152996 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1653
timestamp 1676037725
transform 1 0 153180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1665
timestamp 1676037725
transform 1 0 154284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1677
timestamp 1676037725
transform 1 0 155388 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1689
timestamp 1676037725
transform 1 0 156492 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1701
timestamp 1676037725
transform 1 0 157596 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1707
timestamp 1676037725
transform 1 0 158148 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1709
timestamp 1676037725
transform 1 0 158332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1721
timestamp 1676037725
transform 1 0 159436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1733
timestamp 1676037725
transform 1 0 160540 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1745
timestamp 1676037725
transform 1 0 161644 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1757
timestamp 1676037725
transform 1 0 162748 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1763
timestamp 1676037725
transform 1 0 163300 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1765
timestamp 1676037725
transform 1 0 163484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1777
timestamp 1676037725
transform 1 0 164588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1789
timestamp 1676037725
transform 1 0 165692 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1801
timestamp 1676037725
transform 1 0 166796 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1813
timestamp 1676037725
transform 1 0 167900 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1819
timestamp 1676037725
transform 1 0 168452 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1821
timestamp 1676037725
transform 1 0 168636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1833
timestamp 1676037725
transform 1 0 169740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1845
timestamp 1676037725
transform 1 0 170844 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1857
timestamp 1676037725
transform 1 0 171948 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1869
timestamp 1676037725
transform 1 0 173052 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1875
timestamp 1676037725
transform 1 0 173604 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1877
timestamp 1676037725
transform 1 0 173788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1889
timestamp 1676037725
transform 1 0 174892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1901
timestamp 1676037725
transform 1 0 175996 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1913
timestamp 1676037725
transform 1 0 177100 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1925
timestamp 1676037725
transform 1 0 178204 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1931
timestamp 1676037725
transform 1 0 178756 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1933
timestamp 1676037725
transform 1 0 178940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1945
timestamp 1676037725
transform 1 0 180044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1957
timestamp 1676037725
transform 1 0 181148 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1969
timestamp 1676037725
transform 1 0 182252 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1981
timestamp 1676037725
transform 1 0 183356 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1987
timestamp 1676037725
transform 1 0 183908 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1989
timestamp 1676037725
transform 1 0 184092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2001
timestamp 1676037725
transform 1 0 185196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2013
timestamp 1676037725
transform 1 0 186300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2025
timestamp 1676037725
transform 1 0 187404 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2037
timestamp 1676037725
transform 1 0 188508 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2043
timestamp 1676037725
transform 1 0 189060 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2045
timestamp 1676037725
transform 1 0 189244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2057
timestamp 1676037725
transform 1 0 190348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2069
timestamp 1676037725
transform 1 0 191452 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2081
timestamp 1676037725
transform 1 0 192556 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2093
timestamp 1676037725
transform 1 0 193660 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2099
timestamp 1676037725
transform 1 0 194212 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2101
timestamp 1676037725
transform 1 0 194396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2113
timestamp 1676037725
transform 1 0 195500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2125
timestamp 1676037725
transform 1 0 196604 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2137
timestamp 1676037725
transform 1 0 197708 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2149
timestamp 1676037725
transform 1 0 198812 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2155
timestamp 1676037725
transform 1 0 199364 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2157
timestamp 1676037725
transform 1 0 199548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2169
timestamp 1676037725
transform 1 0 200652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2181
timestamp 1676037725
transform 1 0 201756 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2193
timestamp 1676037725
transform 1 0 202860 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2205
timestamp 1676037725
transform 1 0 203964 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2211
timestamp 1676037725
transform 1 0 204516 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2213
timestamp 1676037725
transform 1 0 204700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2225
timestamp 1676037725
transform 1 0 205804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2237
timestamp 1676037725
transform 1 0 206908 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2249
timestamp 1676037725
transform 1 0 208012 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2261
timestamp 1676037725
transform 1 0 209116 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2267
timestamp 1676037725
transform 1 0 209668 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_2269
timestamp 1676037725
transform 1 0 209852 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_2280
timestamp 1676037725
transform 1 0 210864 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2286
timestamp 1676037725
transform 1 0 211416 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2298
timestamp 1676037725
transform 1 0 212520 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2310
timestamp 1676037725
transform 1 0 213624 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_2322
timestamp 1676037725
transform 1 0 214728 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2325
timestamp 1676037725
transform 1 0 215004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2337
timestamp 1676037725
transform 1 0 216108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2349
timestamp 1676037725
transform 1 0 217212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2361
timestamp 1676037725
transform 1 0 218316 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2373
timestamp 1676037725
transform 1 0 219420 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2379
timestamp 1676037725
transform 1 0 219972 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2381
timestamp 1676037725
transform 1 0 220156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2393
timestamp 1676037725
transform 1 0 221260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2405
timestamp 1676037725
transform 1 0 222364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2417
timestamp 1676037725
transform 1 0 223468 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2429
timestamp 1676037725
transform 1 0 224572 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2435
timestamp 1676037725
transform 1 0 225124 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2437
timestamp 1676037725
transform 1 0 225308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2449
timestamp 1676037725
transform 1 0 226412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2461
timestamp 1676037725
transform 1 0 227516 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2473
timestamp 1676037725
transform 1 0 228620 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2485
timestamp 1676037725
transform 1 0 229724 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2491
timestamp 1676037725
transform 1 0 230276 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2493
timestamp 1676037725
transform 1 0 230460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2505
timestamp 1676037725
transform 1 0 231564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2517
timestamp 1676037725
transform 1 0 232668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2529
timestamp 1676037725
transform 1 0 233772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2541
timestamp 1676037725
transform 1 0 234876 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2547
timestamp 1676037725
transform 1 0 235428 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2549
timestamp 1676037725
transform 1 0 235612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2561
timestamp 1676037725
transform 1 0 236716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2573
timestamp 1676037725
transform 1 0 237820 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2585
timestamp 1676037725
transform 1 0 238924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2597
timestamp 1676037725
transform 1 0 240028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2603
timestamp 1676037725
transform 1 0 240580 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2605
timestamp 1676037725
transform 1 0 240764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2617
timestamp 1676037725
transform 1 0 241868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2629
timestamp 1676037725
transform 1 0 242972 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2641
timestamp 1676037725
transform 1 0 244076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2653
timestamp 1676037725
transform 1 0 245180 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2659
timestamp 1676037725
transform 1 0 245732 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2661
timestamp 1676037725
transform 1 0 245916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2673
timestamp 1676037725
transform 1 0 247020 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2685
timestamp 1676037725
transform 1 0 248124 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_2693
timestamp 1676037725
transform 1 0 248860 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_2706
timestamp 1676037725
transform 1 0 250056 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_2714
timestamp 1676037725
transform 1 0 250792 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2717
timestamp 1676037725
transform 1 0 251068 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2729
timestamp 1676037725
transform 1 0 252172 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2741
timestamp 1676037725
transform 1 0 253276 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2753
timestamp 1676037725
transform 1 0 254380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2765
timestamp 1676037725
transform 1 0 255484 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2771
timestamp 1676037725
transform 1 0 256036 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2773
timestamp 1676037725
transform 1 0 256220 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2785
timestamp 1676037725
transform 1 0 257324 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2797
timestamp 1676037725
transform 1 0 258428 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2809
timestamp 1676037725
transform 1 0 259532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2821
timestamp 1676037725
transform 1 0 260636 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2827
timestamp 1676037725
transform 1 0 261188 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2829
timestamp 1676037725
transform 1 0 261372 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2841
timestamp 1676037725
transform 1 0 262476 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_2853
timestamp 1676037725
transform 1 0 263580 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2857
timestamp 1676037725
transform 1 0 263948 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_2860
timestamp 1676037725
transform 1 0 264224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_2873
timestamp 1676037725
transform 1 0 265420 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_2881
timestamp 1676037725
transform 1 0 266156 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2885
timestamp 1676037725
transform 1 0 266524 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2897
timestamp 1676037725
transform 1 0 267628 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2909
timestamp 1676037725
transform 1 0 268732 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2921
timestamp 1676037725
transform 1 0 269836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2933
timestamp 1676037725
transform 1 0 270940 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2939
timestamp 1676037725
transform 1 0 271492 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2941
timestamp 1676037725
transform 1 0 271676 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2953
timestamp 1676037725
transform 1 0 272780 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2965
timestamp 1676037725
transform 1 0 273884 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2977
timestamp 1676037725
transform 1 0 274988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2989
timestamp 1676037725
transform 1 0 276092 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2995
timestamp 1676037725
transform 1 0 276644 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2997
timestamp 1676037725
transform 1 0 276828 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3009
timestamp 1676037725
transform 1 0 277932 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3021
timestamp 1676037725
transform 1 0 279036 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3033
timestamp 1676037725
transform 1 0 280140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3045
timestamp 1676037725
transform 1 0 281244 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3051
timestamp 1676037725
transform 1 0 281796 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3053
timestamp 1676037725
transform 1 0 281980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3065
timestamp 1676037725
transform 1 0 283084 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3077
timestamp 1676037725
transform 1 0 284188 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3089
timestamp 1676037725
transform 1 0 285292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3101
timestamp 1676037725
transform 1 0 286396 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3107
timestamp 1676037725
transform 1 0 286948 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3109
timestamp 1676037725
transform 1 0 287132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3121
timestamp 1676037725
transform 1 0 288236 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3133
timestamp 1676037725
transform 1 0 289340 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3145
timestamp 1676037725
transform 1 0 290444 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3157
timestamp 1676037725
transform 1 0 291548 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3163
timestamp 1676037725
transform 1 0 292100 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3165
timestamp 1676037725
transform 1 0 292284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3177
timestamp 1676037725
transform 1 0 293388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3189
timestamp 1676037725
transform 1 0 294492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3194
timestamp 1676037725
transform 1 0 294952 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3207
timestamp 1676037725
transform 1 0 296148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3219
timestamp 1676037725
transform 1 0 297252 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3221
timestamp 1676037725
transform 1 0 297436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3233
timestamp 1676037725
transform 1 0 298540 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3245
timestamp 1676037725
transform 1 0 299644 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3257
timestamp 1676037725
transform 1 0 300748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3269
timestamp 1676037725
transform 1 0 301852 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3275
timestamp 1676037725
transform 1 0 302404 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3277
timestamp 1676037725
transform 1 0 302588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3289
timestamp 1676037725
transform 1 0 303692 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3301
timestamp 1676037725
transform 1 0 304796 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3313
timestamp 1676037725
transform 1 0 305900 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3325
timestamp 1676037725
transform 1 0 307004 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3331
timestamp 1676037725
transform 1 0 307556 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3333
timestamp 1676037725
transform 1 0 307740 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3344
timestamp 1676037725
transform 1 0 308752 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3364
timestamp 1676037725
transform 1 0 310592 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3377
timestamp 1676037725
transform 1 0 311788 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3385
timestamp 1676037725
transform 1 0 312524 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3389
timestamp 1676037725
transform 1 0 312892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3401
timestamp 1676037725
transform 1 0 313996 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3413
timestamp 1676037725
transform 1 0 315100 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3425
timestamp 1676037725
transform 1 0 316204 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3437
timestamp 1676037725
transform 1 0 317308 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3443
timestamp 1676037725
transform 1 0 317860 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3445
timestamp 1676037725
transform 1 0 318044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3457
timestamp 1676037725
transform 1 0 319148 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3469
timestamp 1676037725
transform 1 0 320252 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3481
timestamp 1676037725
transform 1 0 321356 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3493
timestamp 1676037725
transform 1 0 322460 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3499
timestamp 1676037725
transform 1 0 323012 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3501
timestamp 1676037725
transform 1 0 323196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3513
timestamp 1676037725
transform 1 0 324300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3525
timestamp 1676037725
transform 1 0 325404 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3537
timestamp 1676037725
transform 1 0 326508 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3549
timestamp 1676037725
transform 1 0 327612 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3555
timestamp 1676037725
transform 1 0 328164 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3557
timestamp 1676037725
transform 1 0 328348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3569
timestamp 1676037725
transform 1 0 329452 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3581
timestamp 1676037725
transform 1 0 330556 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3593
timestamp 1676037725
transform 1 0 331660 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3605
timestamp 1676037725
transform 1 0 332764 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3611
timestamp 1676037725
transform 1 0 333316 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3613
timestamp 1676037725
transform 1 0 333500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3625
timestamp 1676037725
transform 1 0 334604 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3637
timestamp 1676037725
transform 1 0 335708 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3649
timestamp 1676037725
transform 1 0 336812 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3661
timestamp 1676037725
transform 1 0 337916 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3667
timestamp 1676037725
transform 1 0 338468 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3669
timestamp 1676037725
transform 1 0 338652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3681
timestamp 1676037725
transform 1 0 339756 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3693
timestamp 1676037725
transform 1 0 340860 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3705
timestamp 1676037725
transform 1 0 341964 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3717
timestamp 1676037725
transform 1 0 343068 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3723
timestamp 1676037725
transform 1 0 343620 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3725
timestamp 1676037725
transform 1 0 343804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3737
timestamp 1676037725
transform 1 0 344908 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3749
timestamp 1676037725
transform 1 0 346012 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3761
timestamp 1676037725
transform 1 0 347116 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3773
timestamp 1676037725
transform 1 0 348220 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3779
timestamp 1676037725
transform 1 0 348772 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3781
timestamp 1676037725
transform 1 0 348956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3793
timestamp 1676037725
transform 1 0 350060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3805
timestamp 1676037725
transform 1 0 351164 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3817
timestamp 1676037725
transform 1 0 352268 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3829
timestamp 1676037725
transform 1 0 353372 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3835
timestamp 1676037725
transform 1 0 353924 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3837
timestamp 1676037725
transform 1 0 354108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3849
timestamp 1676037725
transform 1 0 355212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3861
timestamp 1676037725
transform 1 0 356316 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3873
timestamp 1676037725
transform 1 0 357420 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3885
timestamp 1676037725
transform 1 0 358524 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3891
timestamp 1676037725
transform 1 0 359076 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3893
timestamp 1676037725
transform 1 0 359260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3905
timestamp 1676037725
transform 1 0 360364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3917
timestamp 1676037725
transform 1 0 361468 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3929
timestamp 1676037725
transform 1 0 362572 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3941
timestamp 1676037725
transform 1 0 363676 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3947
timestamp 1676037725
transform 1 0 364228 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3949
timestamp 1676037725
transform 1 0 364412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3961
timestamp 1676037725
transform 1 0 365516 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3973
timestamp 1676037725
transform 1 0 366620 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3985
timestamp 1676037725
transform 1 0 367724 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3997
timestamp 1676037725
transform 1 0 368828 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4003
timestamp 1676037725
transform 1 0 369380 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4005
timestamp 1676037725
transform 1 0 369564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4017
timestamp 1676037725
transform 1 0 370668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4029
timestamp 1676037725
transform 1 0 371772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4041
timestamp 1676037725
transform 1 0 372876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4053
timestamp 1676037725
transform 1 0 373980 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4059
timestamp 1676037725
transform 1 0 374532 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4061
timestamp 1676037725
transform 1 0 374716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4073
timestamp 1676037725
transform 1 0 375820 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4085
timestamp 1676037725
transform 1 0 376924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4097
timestamp 1676037725
transform 1 0 378028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4109
timestamp 1676037725
transform 1 0 379132 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4115
timestamp 1676037725
transform 1 0 379684 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4117
timestamp 1676037725
transform 1 0 379868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4129
timestamp 1676037725
transform 1 0 380972 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4141
timestamp 1676037725
transform 1 0 382076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4153
timestamp 1676037725
transform 1 0 383180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4165
timestamp 1676037725
transform 1 0 384284 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4171
timestamp 1676037725
transform 1 0 384836 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4173
timestamp 1676037725
transform 1 0 385020 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4185
timestamp 1676037725
transform 1 0 386124 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4197
timestamp 1676037725
transform 1 0 387228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4209
timestamp 1676037725
transform 1 0 388332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4221
timestamp 1676037725
transform 1 0 389436 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4227
timestamp 1676037725
transform 1 0 389988 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4229
timestamp 1676037725
transform 1 0 390172 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4241
timestamp 1676037725
transform 1 0 391276 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4253
timestamp 1676037725
transform 1 0 392380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4265
timestamp 1676037725
transform 1 0 393484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4277
timestamp 1676037725
transform 1 0 394588 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4283
timestamp 1676037725
transform 1 0 395140 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4285
timestamp 1676037725
transform 1 0 395324 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4297
timestamp 1676037725
transform 1 0 396428 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4309
timestamp 1676037725
transform 1 0 397532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4321
timestamp 1676037725
transform 1 0 398636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4333
timestamp 1676037725
transform 1 0 399740 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4339
timestamp 1676037725
transform 1 0 400292 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4341
timestamp 1676037725
transform 1 0 400476 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4353
timestamp 1676037725
transform 1 0 401580 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4365
timestamp 1676037725
transform 1 0 402684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_4377
timestamp 1676037725
transform 1 0 403788 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_4394
timestamp 1676037725
transform 1 0 405352 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_4397
timestamp 1676037725
transform 1 0 405628 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4401
timestamp 1676037725
transform 1 0 405996 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4413
timestamp 1676037725
transform 1 0 407100 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4425
timestamp 1676037725
transform 1 0 408204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4437
timestamp 1676037725
transform 1 0 409308 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_4449
timestamp 1676037725
transform 1 0 410412 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4453
timestamp 1676037725
transform 1 0 410780 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4465
timestamp 1676037725
transform 1 0 411884 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4477
timestamp 1676037725
transform 1 0 412988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4489
timestamp 1676037725
transform 1 0 414092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4501
timestamp 1676037725
transform 1 0 415196 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4507
timestamp 1676037725
transform 1 0 415748 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4509
timestamp 1676037725
transform 1 0 415932 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4521
timestamp 1676037725
transform 1 0 417036 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4533
timestamp 1676037725
transform 1 0 418140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4545
timestamp 1676037725
transform 1 0 419244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4557
timestamp 1676037725
transform 1 0 420348 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4563
timestamp 1676037725
transform 1 0 420900 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4565
timestamp 1676037725
transform 1 0 421084 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4577
timestamp 1676037725
transform 1 0 422188 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4589
timestamp 1676037725
transform 1 0 423292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4601
timestamp 1676037725
transform 1 0 424396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4613
timestamp 1676037725
transform 1 0 425500 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4619
timestamp 1676037725
transform 1 0 426052 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4621
timestamp 1676037725
transform 1 0 426236 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4633
timestamp 1676037725
transform 1 0 427340 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4645
timestamp 1676037725
transform 1 0 428444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4657
timestamp 1676037725
transform 1 0 429548 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4669
timestamp 1676037725
transform 1 0 430652 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4675
timestamp 1676037725
transform 1 0 431204 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4677
timestamp 1676037725
transform 1 0 431388 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4689
timestamp 1676037725
transform 1 0 432492 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4701
timestamp 1676037725
transform 1 0 433596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4713
timestamp 1676037725
transform 1 0 434700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4725
timestamp 1676037725
transform 1 0 435804 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4731
timestamp 1676037725
transform 1 0 436356 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4733
timestamp 1676037725
transform 1 0 436540 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4745
timestamp 1676037725
transform 1 0 437644 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4757
timestamp 1676037725
transform 1 0 438748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4769
timestamp 1676037725
transform 1 0 439852 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4781
timestamp 1676037725
transform 1 0 440956 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4787
timestamp 1676037725
transform 1 0 441508 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4789
timestamp 1676037725
transform 1 0 441692 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4801
timestamp 1676037725
transform 1 0 442796 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4813
timestamp 1676037725
transform 1 0 443900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4825
timestamp 1676037725
transform 1 0 445004 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4837
timestamp 1676037725
transform 1 0 446108 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4843
timestamp 1676037725
transform 1 0 446660 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4845
timestamp 1676037725
transform 1 0 446844 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4857
timestamp 1676037725
transform 1 0 447948 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4869
timestamp 1676037725
transform 1 0 449052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4881
timestamp 1676037725
transform 1 0 450156 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4893
timestamp 1676037725
transform 1 0 451260 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4899
timestamp 1676037725
transform 1 0 451812 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4901
timestamp 1676037725
transform 1 0 451996 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4913
timestamp 1676037725
transform 1 0 453100 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4925
timestamp 1676037725
transform 1 0 454204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4937
timestamp 1676037725
transform 1 0 455308 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4949
timestamp 1676037725
transform 1 0 456412 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4955
timestamp 1676037725
transform 1 0 456964 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4957
timestamp 1676037725
transform 1 0 457148 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4969
timestamp 1676037725
transform 1 0 458252 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4981
timestamp 1676037725
transform 1 0 459356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4993
timestamp 1676037725
transform 1 0 460460 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5005
timestamp 1676037725
transform 1 0 461564 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5011
timestamp 1676037725
transform 1 0 462116 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5013
timestamp 1676037725
transform 1 0 462300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5025
timestamp 1676037725
transform 1 0 463404 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5037
timestamp 1676037725
transform 1 0 464508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5049
timestamp 1676037725
transform 1 0 465612 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5061
timestamp 1676037725
transform 1 0 466716 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5067
timestamp 1676037725
transform 1 0 467268 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5069
timestamp 1676037725
transform 1 0 467452 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5081
timestamp 1676037725
transform 1 0 468556 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5093
timestamp 1676037725
transform 1 0 469660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5105
timestamp 1676037725
transform 1 0 470764 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5117
timestamp 1676037725
transform 1 0 471868 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5123
timestamp 1676037725
transform 1 0 472420 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5125
timestamp 1676037725
transform 1 0 472604 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5137
timestamp 1676037725
transform 1 0 473708 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5149
timestamp 1676037725
transform 1 0 474812 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5161
timestamp 1676037725
transform 1 0 475916 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5173
timestamp 1676037725
transform 1 0 477020 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5179
timestamp 1676037725
transform 1 0 477572 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5181
timestamp 1676037725
transform 1 0 477756 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5193
timestamp 1676037725
transform 1 0 478860 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5205
timestamp 1676037725
transform 1 0 479964 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5217
timestamp 1676037725
transform 1 0 481068 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5229
timestamp 1676037725
transform 1 0 482172 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5235
timestamp 1676037725
transform 1 0 482724 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5237
timestamp 1676037725
transform 1 0 482908 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5249
timestamp 1676037725
transform 1 0 484012 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5261
timestamp 1676037725
transform 1 0 485116 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5273
timestamp 1676037725
transform 1 0 486220 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5285
timestamp 1676037725
transform 1 0 487324 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5291
timestamp 1676037725
transform 1 0 487876 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5293
timestamp 1676037725
transform 1 0 488060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5305
timestamp 1676037725
transform 1 0 489164 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5317
timestamp 1676037725
transform 1 0 490268 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5329
timestamp 1676037725
transform 1 0 491372 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5341
timestamp 1676037725
transform 1 0 492476 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5347
timestamp 1676037725
transform 1 0 493028 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5349
timestamp 1676037725
transform 1 0 493212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5361
timestamp 1676037725
transform 1 0 494316 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5373
timestamp 1676037725
transform 1 0 495420 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5385
timestamp 1676037725
transform 1 0 496524 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5397
timestamp 1676037725
transform 1 0 497628 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5403
timestamp 1676037725
transform 1 0 498180 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5405
timestamp 1676037725
transform 1 0 498364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5417
timestamp 1676037725
transform 1 0 499468 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5429
timestamp 1676037725
transform 1 0 500572 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5441
timestamp 1676037725
transform 1 0 501676 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5453
timestamp 1676037725
transform 1 0 502780 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5459
timestamp 1676037725
transform 1 0 503332 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5461
timestamp 1676037725
transform 1 0 503516 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5473
timestamp 1676037725
transform 1 0 504620 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5485
timestamp 1676037725
transform 1 0 505724 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5497
timestamp 1676037725
transform 1 0 506828 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5509
timestamp 1676037725
transform 1 0 507932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5515
timestamp 1676037725
transform 1 0 508484 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5517
timestamp 1676037725
transform 1 0 508668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5529
timestamp 1676037725
transform 1 0 509772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5541
timestamp 1676037725
transform 1 0 510876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5553
timestamp 1676037725
transform 1 0 511980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5565
timestamp 1676037725
transform 1 0 513084 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5571
timestamp 1676037725
transform 1 0 513636 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5573
timestamp 1676037725
transform 1 0 513820 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5585
timestamp 1676037725
transform 1 0 514924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5597
timestamp 1676037725
transform 1 0 516028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5609
timestamp 1676037725
transform 1 0 517132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5621
timestamp 1676037725
transform 1 0 518236 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5627
timestamp 1676037725
transform 1 0 518788 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5629
timestamp 1676037725
transform 1 0 518972 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5641
timestamp 1676037725
transform 1 0 520076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5653
timestamp 1676037725
transform 1 0 521180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5665
timestamp 1676037725
transform 1 0 522284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5677
timestamp 1676037725
transform 1 0 523388 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5683
timestamp 1676037725
transform 1 0 523940 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5685
timestamp 1676037725
transform 1 0 524124 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5697
timestamp 1676037725
transform 1 0 525228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5709
timestamp 1676037725
transform 1 0 526332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5721
timestamp 1676037725
transform 1 0 527436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5733
timestamp 1676037725
transform 1 0 528540 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5739
timestamp 1676037725
transform 1 0 529092 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5741
timestamp 1676037725
transform 1 0 529276 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5753
timestamp 1676037725
transform 1 0 530380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5765
timestamp 1676037725
transform 1 0 531484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5777
timestamp 1676037725
transform 1 0 532588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5789
timestamp 1676037725
transform 1 0 533692 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5795
timestamp 1676037725
transform 1 0 534244 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5797
timestamp 1676037725
transform 1 0 534428 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5809
timestamp 1676037725
transform 1 0 535532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5821
timestamp 1676037725
transform 1 0 536636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5833
timestamp 1676037725
transform 1 0 537740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5845
timestamp 1676037725
transform 1 0 538844 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5851
timestamp 1676037725
transform 1 0 539396 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5853
timestamp 1676037725
transform 1 0 539580 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5865
timestamp 1676037725
transform 1 0 540684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5877
timestamp 1676037725
transform 1 0 541788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5889
timestamp 1676037725
transform 1 0 542892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5901
timestamp 1676037725
transform 1 0 543996 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5907
timestamp 1676037725
transform 1 0 544548 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5909
timestamp 1676037725
transform 1 0 544732 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5921
timestamp 1676037725
transform 1 0 545836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5933
timestamp 1676037725
transform 1 0 546940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5945
timestamp 1676037725
transform 1 0 548044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5957
timestamp 1676037725
transform 1 0 549148 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5963
timestamp 1676037725
transform 1 0 549700 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5965
timestamp 1676037725
transform 1 0 549884 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5977
timestamp 1676037725
transform 1 0 550988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5989
timestamp 1676037725
transform 1 0 552092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6001
timestamp 1676037725
transform 1 0 553196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6013
timestamp 1676037725
transform 1 0 554300 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6019
timestamp 1676037725
transform 1 0 554852 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6021
timestamp 1676037725
transform 1 0 555036 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6033
timestamp 1676037725
transform 1 0 556140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6045
timestamp 1676037725
transform 1 0 557244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6057
timestamp 1676037725
transform 1 0 558348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6069
timestamp 1676037725
transform 1 0 559452 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6075
timestamp 1676037725
transform 1 0 560004 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6077
timestamp 1676037725
transform 1 0 560188 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6089
timestamp 1676037725
transform 1 0 561292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6101
timestamp 1676037725
transform 1 0 562396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6113
timestamp 1676037725
transform 1 0 563500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6125
timestamp 1676037725
transform 1 0 564604 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6131
timestamp 1676037725
transform 1 0 565156 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6133
timestamp 1676037725
transform 1 0 565340 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6145
timestamp 1676037725
transform 1 0 566444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6157
timestamp 1676037725
transform 1 0 567548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6169
timestamp 1676037725
transform 1 0 568652 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6181
timestamp 1676037725
transform 1 0 569756 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6187
timestamp 1676037725
transform 1 0 570308 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6189
timestamp 1676037725
transform 1 0 570492 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6201
timestamp 1676037725
transform 1 0 571596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6213
timestamp 1676037725
transform 1 0 572700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6225
timestamp 1676037725
transform 1 0 573804 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6237
timestamp 1676037725
transform 1 0 574908 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6243
timestamp 1676037725
transform 1 0 575460 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6245
timestamp 1676037725
transform 1 0 575644 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6257
timestamp 1676037725
transform 1 0 576748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6269
timestamp 1676037725
transform 1 0 577852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6281
timestamp 1676037725
transform 1 0 578956 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6293
timestamp 1676037725
transform 1 0 580060 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6299
timestamp 1676037725
transform 1 0 580612 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6301
timestamp 1676037725
transform 1 0 580796 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6313
timestamp 1676037725
transform 1 0 581900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6325
timestamp 1676037725
transform 1 0 583004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6337
timestamp 1676037725
transform 1 0 584108 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6349
timestamp 1676037725
transform 1 0 585212 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6355
timestamp 1676037725
transform 1 0 585764 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6357
timestamp 1676037725
transform 1 0 585948 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6369
timestamp 1676037725
transform 1 0 587052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6381
timestamp 1676037725
transform 1 0 588156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6393
timestamp 1676037725
transform 1 0 589260 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6405
timestamp 1676037725
transform 1 0 590364 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6411
timestamp 1676037725
transform 1 0 590916 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6413
timestamp 1676037725
transform 1 0 591100 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6425
timestamp 1676037725
transform 1 0 592204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6437
timestamp 1676037725
transform 1 0 593308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6449
timestamp 1676037725
transform 1 0 594412 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6461
timestamp 1676037725
transform 1 0 595516 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6467
timestamp 1676037725
transform 1 0 596068 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6469
timestamp 1676037725
transform 1 0 596252 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6481
timestamp 1676037725
transform 1 0 597356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6493
timestamp 1676037725
transform 1 0 598460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6505
timestamp 1676037725
transform 1 0 599564 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6517
timestamp 1676037725
transform 1 0 600668 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6523
timestamp 1676037725
transform 1 0 601220 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6525
timestamp 1676037725
transform 1 0 601404 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6537
timestamp 1676037725
transform 1 0 602508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6549
timestamp 1676037725
transform 1 0 603612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6561
timestamp 1676037725
transform 1 0 604716 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6573
timestamp 1676037725
transform 1 0 605820 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6579
timestamp 1676037725
transform 1 0 606372 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6581
timestamp 1676037725
transform 1 0 606556 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6593
timestamp 1676037725
transform 1 0 607660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6605
timestamp 1676037725
transform 1 0 608764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6617
timestamp 1676037725
transform 1 0 609868 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6629
timestamp 1676037725
transform 1 0 610972 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6635
timestamp 1676037725
transform 1 0 611524 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6637
timestamp 1676037725
transform 1 0 611708 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6649
timestamp 1676037725
transform 1 0 612812 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6661
timestamp 1676037725
transform 1 0 613916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6673
timestamp 1676037725
transform 1 0 615020 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6685
timestamp 1676037725
transform 1 0 616124 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6691
timestamp 1676037725
transform 1 0 616676 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6693
timestamp 1676037725
transform 1 0 616860 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6705
timestamp 1676037725
transform 1 0 617964 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6717
timestamp 1676037725
transform 1 0 619068 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6729
timestamp 1676037725
transform 1 0 620172 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6741
timestamp 1676037725
transform 1 0 621276 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6747
timestamp 1676037725
transform 1 0 621828 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6749
timestamp 1676037725
transform 1 0 622012 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6761
timestamp 1676037725
transform 1 0 623116 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6773
timestamp 1676037725
transform 1 0 624220 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6785
timestamp 1676037725
transform 1 0 625324 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6797
timestamp 1676037725
transform 1 0 626428 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6803
timestamp 1676037725
transform 1 0 626980 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6805
timestamp 1676037725
transform 1 0 627164 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6817
timestamp 1676037725
transform 1 0 628268 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6829
timestamp 1676037725
transform 1 0 629372 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6841
timestamp 1676037725
transform 1 0 630476 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6853
timestamp 1676037725
transform 1 0 631580 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6859
timestamp 1676037725
transform 1 0 632132 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6861
timestamp 1676037725
transform 1 0 632316 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6873
timestamp 1676037725
transform 1 0 633420 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6885
timestamp 1676037725
transform 1 0 634524 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6897
timestamp 1676037725
transform 1 0 635628 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6909
timestamp 1676037725
transform 1 0 636732 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6915
timestamp 1676037725
transform 1 0 637284 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6917
timestamp 1676037725
transform 1 0 637468 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6929
timestamp 1676037725
transform 1 0 638572 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6941
timestamp 1676037725
transform 1 0 639676 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6953
timestamp 1676037725
transform 1 0 640780 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6965
timestamp 1676037725
transform 1 0 641884 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6971
timestamp 1676037725
transform 1 0 642436 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6973
timestamp 1676037725
transform 1 0 642620 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6985
timestamp 1676037725
transform 1 0 643724 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6997
timestamp 1676037725
transform 1 0 644828 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7009
timestamp 1676037725
transform 1 0 645932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_7021
timestamp 1676037725
transform 1 0 647036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7027
timestamp 1676037725
transform 1 0 647588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_7029
timestamp 1676037725
transform 1 0 647772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7037
timestamp 1676037725
transform 1 0 648508 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1676037725
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1676037725
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1676037725
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1676037725
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1676037725
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1676037725
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1676037725
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1676037725
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1676037725
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1676037725
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1676037725
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1676037725
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1676037725
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1676037725
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1676037725
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1676037725
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1676037725
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1676037725
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1676037725
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1676037725
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1676037725
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1676037725
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1676037725
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1676037725
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1676037725
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1676037725
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1676037725
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1676037725
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1676037725
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1676037725
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1676037725
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1676037725
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1676037725
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1676037725
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1676037725
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1676037725
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 1676037725
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1676037725
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1676037725
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1676037725
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_809
timestamp 1676037725
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_821
timestamp 1676037725
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_833
timestamp 1676037725
transform 1 0 77740 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_839
timestamp 1676037725
transform 1 0 78292 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_841
timestamp 1676037725
transform 1 0 78476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_853
timestamp 1676037725
transform 1 0 79580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_865
timestamp 1676037725
transform 1 0 80684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_877
timestamp 1676037725
transform 1 0 81788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_889
timestamp 1676037725
transform 1 0 82892 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_895
timestamp 1676037725
transform 1 0 83444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_897
timestamp 1676037725
transform 1 0 83628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_909
timestamp 1676037725
transform 1 0 84732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_921
timestamp 1676037725
transform 1 0 85836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_933
timestamp 1676037725
transform 1 0 86940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_945
timestamp 1676037725
transform 1 0 88044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_951
timestamp 1676037725
transform 1 0 88596 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_953
timestamp 1676037725
transform 1 0 88780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_965
timestamp 1676037725
transform 1 0 89884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_977
timestamp 1676037725
transform 1 0 90988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_989
timestamp 1676037725
transform 1 0 92092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1001
timestamp 1676037725
transform 1 0 93196 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1007
timestamp 1676037725
transform 1 0 93748 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1009
timestamp 1676037725
transform 1 0 93932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1021
timestamp 1676037725
transform 1 0 95036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1033
timestamp 1676037725
transform 1 0 96140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1045
timestamp 1676037725
transform 1 0 97244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1057
timestamp 1676037725
transform 1 0 98348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1063
timestamp 1676037725
transform 1 0 98900 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1065
timestamp 1676037725
transform 1 0 99084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1077
timestamp 1676037725
transform 1 0 100188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1089
timestamp 1676037725
transform 1 0 101292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1101
timestamp 1676037725
transform 1 0 102396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1113
timestamp 1676037725
transform 1 0 103500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1119
timestamp 1676037725
transform 1 0 104052 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1121
timestamp 1676037725
transform 1 0 104236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1133
timestamp 1676037725
transform 1 0 105340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1145
timestamp 1676037725
transform 1 0 106444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1157
timestamp 1676037725
transform 1 0 107548 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1169
timestamp 1676037725
transform 1 0 108652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1175
timestamp 1676037725
transform 1 0 109204 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1177
timestamp 1676037725
transform 1 0 109388 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1189
timestamp 1676037725
transform 1 0 110492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1201
timestamp 1676037725
transform 1 0 111596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1213
timestamp 1676037725
transform 1 0 112700 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1225
timestamp 1676037725
transform 1 0 113804 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1231
timestamp 1676037725
transform 1 0 114356 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1233
timestamp 1676037725
transform 1 0 114540 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1245
timestamp 1676037725
transform 1 0 115644 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1257
timestamp 1676037725
transform 1 0 116748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1269
timestamp 1676037725
transform 1 0 117852 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1281
timestamp 1676037725
transform 1 0 118956 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1287
timestamp 1676037725
transform 1 0 119508 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1289
timestamp 1676037725
transform 1 0 119692 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1301
timestamp 1676037725
transform 1 0 120796 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1313
timestamp 1676037725
transform 1 0 121900 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1325
timestamp 1676037725
transform 1 0 123004 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1337
timestamp 1676037725
transform 1 0 124108 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1343
timestamp 1676037725
transform 1 0 124660 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1345
timestamp 1676037725
transform 1 0 124844 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1357
timestamp 1676037725
transform 1 0 125948 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1369
timestamp 1676037725
transform 1 0 127052 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1381
timestamp 1676037725
transform 1 0 128156 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1393
timestamp 1676037725
transform 1 0 129260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1399
timestamp 1676037725
transform 1 0 129812 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1401
timestamp 1676037725
transform 1 0 129996 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1413
timestamp 1676037725
transform 1 0 131100 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1425
timestamp 1676037725
transform 1 0 132204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1437
timestamp 1676037725
transform 1 0 133308 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1449
timestamp 1676037725
transform 1 0 134412 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1455
timestamp 1676037725
transform 1 0 134964 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1457
timestamp 1676037725
transform 1 0 135148 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1469
timestamp 1676037725
transform 1 0 136252 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1481
timestamp 1676037725
transform 1 0 137356 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1493
timestamp 1676037725
transform 1 0 138460 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1505
timestamp 1676037725
transform 1 0 139564 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1511
timestamp 1676037725
transform 1 0 140116 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1513
timestamp 1676037725
transform 1 0 140300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1525
timestamp 1676037725
transform 1 0 141404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1537
timestamp 1676037725
transform 1 0 142508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1549
timestamp 1676037725
transform 1 0 143612 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1561
timestamp 1676037725
transform 1 0 144716 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1567
timestamp 1676037725
transform 1 0 145268 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1569
timestamp 1676037725
transform 1 0 145452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1581
timestamp 1676037725
transform 1 0 146556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1593
timestamp 1676037725
transform 1 0 147660 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1605
timestamp 1676037725
transform 1 0 148764 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1617
timestamp 1676037725
transform 1 0 149868 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1623
timestamp 1676037725
transform 1 0 150420 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1625
timestamp 1676037725
transform 1 0 150604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1637
timestamp 1676037725
transform 1 0 151708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1649
timestamp 1676037725
transform 1 0 152812 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1661
timestamp 1676037725
transform 1 0 153916 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1673
timestamp 1676037725
transform 1 0 155020 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1679
timestamp 1676037725
transform 1 0 155572 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1681
timestamp 1676037725
transform 1 0 155756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1693
timestamp 1676037725
transform 1 0 156860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1705
timestamp 1676037725
transform 1 0 157964 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1717
timestamp 1676037725
transform 1 0 159068 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1729
timestamp 1676037725
transform 1 0 160172 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1735
timestamp 1676037725
transform 1 0 160724 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1737
timestamp 1676037725
transform 1 0 160908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1749
timestamp 1676037725
transform 1 0 162012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1761
timestamp 1676037725
transform 1 0 163116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1773
timestamp 1676037725
transform 1 0 164220 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1785
timestamp 1676037725
transform 1 0 165324 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1791
timestamp 1676037725
transform 1 0 165876 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1793
timestamp 1676037725
transform 1 0 166060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1805
timestamp 1676037725
transform 1 0 167164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1817
timestamp 1676037725
transform 1 0 168268 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1829
timestamp 1676037725
transform 1 0 169372 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1841
timestamp 1676037725
transform 1 0 170476 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1847
timestamp 1676037725
transform 1 0 171028 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1849
timestamp 1676037725
transform 1 0 171212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1861
timestamp 1676037725
transform 1 0 172316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1873
timestamp 1676037725
transform 1 0 173420 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1885
timestamp 1676037725
transform 1 0 174524 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1897
timestamp 1676037725
transform 1 0 175628 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1903
timestamp 1676037725
transform 1 0 176180 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1905
timestamp 1676037725
transform 1 0 176364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1917
timestamp 1676037725
transform 1 0 177468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1929
timestamp 1676037725
transform 1 0 178572 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1941
timestamp 1676037725
transform 1 0 179676 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1953
timestamp 1676037725
transform 1 0 180780 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1959
timestamp 1676037725
transform 1 0 181332 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1961
timestamp 1676037725
transform 1 0 181516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1973
timestamp 1676037725
transform 1 0 182620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1985
timestamp 1676037725
transform 1 0 183724 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1997
timestamp 1676037725
transform 1 0 184828 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2009
timestamp 1676037725
transform 1 0 185932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2015
timestamp 1676037725
transform 1 0 186484 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2017
timestamp 1676037725
transform 1 0 186668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2029
timestamp 1676037725
transform 1 0 187772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2041
timestamp 1676037725
transform 1 0 188876 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2053
timestamp 1676037725
transform 1 0 189980 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2065
timestamp 1676037725
transform 1 0 191084 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2071
timestamp 1676037725
transform 1 0 191636 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2073
timestamp 1676037725
transform 1 0 191820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2085
timestamp 1676037725
transform 1 0 192924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2097
timestamp 1676037725
transform 1 0 194028 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2109
timestamp 1676037725
transform 1 0 195132 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2121
timestamp 1676037725
transform 1 0 196236 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2127
timestamp 1676037725
transform 1 0 196788 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2129
timestamp 1676037725
transform 1 0 196972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2141
timestamp 1676037725
transform 1 0 198076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2153
timestamp 1676037725
transform 1 0 199180 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2165
timestamp 1676037725
transform 1 0 200284 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2177
timestamp 1676037725
transform 1 0 201388 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2183
timestamp 1676037725
transform 1 0 201940 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2185
timestamp 1676037725
transform 1 0 202124 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_2193
timestamp 1676037725
transform 1 0 202860 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2206
timestamp 1676037725
transform 1 0 204056 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2218
timestamp 1676037725
transform 1 0 205160 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_2230
timestamp 1676037725
transform 1 0 206264 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_2238
timestamp 1676037725
transform 1 0 207000 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2241
timestamp 1676037725
transform 1 0 207276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2253
timestamp 1676037725
transform 1 0 208380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2265
timestamp 1676037725
transform 1 0 209484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2277
timestamp 1676037725
transform 1 0 210588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2289
timestamp 1676037725
transform 1 0 211692 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2295
timestamp 1676037725
transform 1 0 212244 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2297
timestamp 1676037725
transform 1 0 212428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2309
timestamp 1676037725
transform 1 0 213532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2321
timestamp 1676037725
transform 1 0 214636 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2333
timestamp 1676037725
transform 1 0 215740 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2345
timestamp 1676037725
transform 1 0 216844 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2351
timestamp 1676037725
transform 1 0 217396 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_2353
timestamp 1676037725
transform 1 0 217580 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_2359
timestamp 1676037725
transform 1 0 218132 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2372
timestamp 1676037725
transform 1 0 219328 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2384
timestamp 1676037725
transform 1 0 220432 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2396
timestamp 1676037725
transform 1 0 221536 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2409
timestamp 1676037725
transform 1 0 222732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2421
timestamp 1676037725
transform 1 0 223836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2433
timestamp 1676037725
transform 1 0 224940 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2445
timestamp 1676037725
transform 1 0 226044 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2457
timestamp 1676037725
transform 1 0 227148 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2463
timestamp 1676037725
transform 1 0 227700 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2465
timestamp 1676037725
transform 1 0 227884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2477
timestamp 1676037725
transform 1 0 228988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2489
timestamp 1676037725
transform 1 0 230092 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2501
timestamp 1676037725
transform 1 0 231196 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2513
timestamp 1676037725
transform 1 0 232300 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2519
timestamp 1676037725
transform 1 0 232852 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2521
timestamp 1676037725
transform 1 0 233036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2533
timestamp 1676037725
transform 1 0 234140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2545
timestamp 1676037725
transform 1 0 235244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2557
timestamp 1676037725
transform 1 0 236348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2569
timestamp 1676037725
transform 1 0 237452 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2575
timestamp 1676037725
transform 1 0 238004 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2577
timestamp 1676037725
transform 1 0 238188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2589
timestamp 1676037725
transform 1 0 239292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2601
timestamp 1676037725
transform 1 0 240396 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2613
timestamp 1676037725
transform 1 0 241500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2625
timestamp 1676037725
transform 1 0 242604 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2631
timestamp 1676037725
transform 1 0 243156 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2633
timestamp 1676037725
transform 1 0 243340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2645
timestamp 1676037725
transform 1 0 244444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2657
timestamp 1676037725
transform 1 0 245548 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2669
timestamp 1676037725
transform 1 0 246652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2681
timestamp 1676037725
transform 1 0 247756 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2687
timestamp 1676037725
transform 1 0 248308 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2689
timestamp 1676037725
transform 1 0 248492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2701
timestamp 1676037725
transform 1 0 249596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2713
timestamp 1676037725
transform 1 0 250700 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2725
timestamp 1676037725
transform 1 0 251804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2737
timestamp 1676037725
transform 1 0 252908 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2743
timestamp 1676037725
transform 1 0 253460 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2745
timestamp 1676037725
transform 1 0 253644 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2757
timestamp 1676037725
transform 1 0 254748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2769
timestamp 1676037725
transform 1 0 255852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2781
timestamp 1676037725
transform 1 0 256956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2793
timestamp 1676037725
transform 1 0 258060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2799
timestamp 1676037725
transform 1 0 258612 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2801
timestamp 1676037725
transform 1 0 258796 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2813
timestamp 1676037725
transform 1 0 259900 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2825
timestamp 1676037725
transform 1 0 261004 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2837
timestamp 1676037725
transform 1 0 262108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2849
timestamp 1676037725
transform 1 0 263212 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2855
timestamp 1676037725
transform 1 0 263764 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2857
timestamp 1676037725
transform 1 0 263948 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2869
timestamp 1676037725
transform 1 0 265052 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2881
timestamp 1676037725
transform 1 0 266156 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2893
timestamp 1676037725
transform 1 0 267260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2905
timestamp 1676037725
transform 1 0 268364 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2911
timestamp 1676037725
transform 1 0 268916 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2913
timestamp 1676037725
transform 1 0 269100 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2925
timestamp 1676037725
transform 1 0 270204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2937
timestamp 1676037725
transform 1 0 271308 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2949
timestamp 1676037725
transform 1 0 272412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2961
timestamp 1676037725
transform 1 0 273516 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2967
timestamp 1676037725
transform 1 0 274068 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2969
timestamp 1676037725
transform 1 0 274252 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2981
timestamp 1676037725
transform 1 0 275356 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2993
timestamp 1676037725
transform 1 0 276460 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3005
timestamp 1676037725
transform 1 0 277564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3017
timestamp 1676037725
transform 1 0 278668 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3023
timestamp 1676037725
transform 1 0 279220 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3025
timestamp 1676037725
transform 1 0 279404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3037
timestamp 1676037725
transform 1 0 280508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3049
timestamp 1676037725
transform 1 0 281612 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3061
timestamp 1676037725
transform 1 0 282716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3073
timestamp 1676037725
transform 1 0 283820 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3079
timestamp 1676037725
transform 1 0 284372 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3081
timestamp 1676037725
transform 1 0 284556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3093
timestamp 1676037725
transform 1 0 285660 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3105
timestamp 1676037725
transform 1 0 286764 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3117
timestamp 1676037725
transform 1 0 287868 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3129
timestamp 1676037725
transform 1 0 288972 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3135
timestamp 1676037725
transform 1 0 289524 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3137
timestamp 1676037725
transform 1 0 289708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3149
timestamp 1676037725
transform 1 0 290812 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3161
timestamp 1676037725
transform 1 0 291916 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3173
timestamp 1676037725
transform 1 0 293020 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3185
timestamp 1676037725
transform 1 0 294124 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3191
timestamp 1676037725
transform 1 0 294676 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3193
timestamp 1676037725
transform 1 0 294860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3205
timestamp 1676037725
transform 1 0 295964 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3217
timestamp 1676037725
transform 1 0 297068 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3229
timestamp 1676037725
transform 1 0 298172 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3241
timestamp 1676037725
transform 1 0 299276 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3247
timestamp 1676037725
transform 1 0 299828 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3249
timestamp 1676037725
transform 1 0 300012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3261
timestamp 1676037725
transform 1 0 301116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3273
timestamp 1676037725
transform 1 0 302220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3285
timestamp 1676037725
transform 1 0 303324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3297
timestamp 1676037725
transform 1 0 304428 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3303
timestamp 1676037725
transform 1 0 304980 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3305
timestamp 1676037725
transform 1 0 305164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3317
timestamp 1676037725
transform 1 0 306268 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3329
timestamp 1676037725
transform 1 0 307372 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3341
timestamp 1676037725
transform 1 0 308476 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3352
timestamp 1676037725
transform 1 0 309488 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3358
timestamp 1676037725
transform 1 0 310040 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3361
timestamp 1676037725
transform 1 0 310316 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3367
timestamp 1676037725
transform 1 0 310868 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3370
timestamp 1676037725
transform 1 0 311144 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3382
timestamp 1676037725
transform 1 0 312248 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3394
timestamp 1676037725
transform 1 0 313352 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3406
timestamp 1676037725
transform 1 0 314456 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3414
timestamp 1676037725
transform 1 0 315192 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3417
timestamp 1676037725
transform 1 0 315468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3429
timestamp 1676037725
transform 1 0 316572 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3441
timestamp 1676037725
transform 1 0 317676 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3453
timestamp 1676037725
transform 1 0 318780 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3465
timestamp 1676037725
transform 1 0 319884 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3471
timestamp 1676037725
transform 1 0 320436 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3473
timestamp 1676037725
transform 1 0 320620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3485
timestamp 1676037725
transform 1 0 321724 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3497
timestamp 1676037725
transform 1 0 322828 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3509
timestamp 1676037725
transform 1 0 323932 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3521
timestamp 1676037725
transform 1 0 325036 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3527
timestamp 1676037725
transform 1 0 325588 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3529
timestamp 1676037725
transform 1 0 325772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3541
timestamp 1676037725
transform 1 0 326876 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3553
timestamp 1676037725
transform 1 0 327980 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3565
timestamp 1676037725
transform 1 0 329084 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3577
timestamp 1676037725
transform 1 0 330188 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3583
timestamp 1676037725
transform 1 0 330740 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3585
timestamp 1676037725
transform 1 0 330924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3597
timestamp 1676037725
transform 1 0 332028 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3609
timestamp 1676037725
transform 1 0 333132 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3621
timestamp 1676037725
transform 1 0 334236 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3633
timestamp 1676037725
transform 1 0 335340 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3639
timestamp 1676037725
transform 1 0 335892 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3641
timestamp 1676037725
transform 1 0 336076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3653
timestamp 1676037725
transform 1 0 337180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3665
timestamp 1676037725
transform 1 0 338284 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3673
timestamp 1676037725
transform 1 0 339020 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3678
timestamp 1676037725
transform 1 0 339480 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3694
timestamp 1676037725
transform 1 0 340952 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3697
timestamp 1676037725
transform 1 0 341228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3709
timestamp 1676037725
transform 1 0 342332 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3721
timestamp 1676037725
transform 1 0 343436 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3733
timestamp 1676037725
transform 1 0 344540 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3745
timestamp 1676037725
transform 1 0 345644 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3751
timestamp 1676037725
transform 1 0 346196 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3753
timestamp 1676037725
transform 1 0 346380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3765
timestamp 1676037725
transform 1 0 347484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3777
timestamp 1676037725
transform 1 0 348588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3789
timestamp 1676037725
transform 1 0 349692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3801
timestamp 1676037725
transform 1 0 350796 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3807
timestamp 1676037725
transform 1 0 351348 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3809
timestamp 1676037725
transform 1 0 351532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3821
timestamp 1676037725
transform 1 0 352636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3833
timestamp 1676037725
transform 1 0 353740 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3841
timestamp 1676037725
transform 1 0 354476 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3846
timestamp 1676037725
transform 1 0 354936 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3862
timestamp 1676037725
transform 1 0 356408 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3865
timestamp 1676037725
transform 1 0 356684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3877
timestamp 1676037725
transform 1 0 357788 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3889
timestamp 1676037725
transform 1 0 358892 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3901
timestamp 1676037725
transform 1 0 359996 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3913
timestamp 1676037725
transform 1 0 361100 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3919
timestamp 1676037725
transform 1 0 361652 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3921
timestamp 1676037725
transform 1 0 361836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3933
timestamp 1676037725
transform 1 0 362940 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3945
timestamp 1676037725
transform 1 0 364044 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3957
timestamp 1676037725
transform 1 0 365148 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3969
timestamp 1676037725
transform 1 0 366252 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3975
timestamp 1676037725
transform 1 0 366804 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3977
timestamp 1676037725
transform 1 0 366988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3989
timestamp 1676037725
transform 1 0 368092 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4001
timestamp 1676037725
transform 1 0 369196 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4013
timestamp 1676037725
transform 1 0 370300 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4025
timestamp 1676037725
transform 1 0 371404 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4031
timestamp 1676037725
transform 1 0 371956 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4033
timestamp 1676037725
transform 1 0 372140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4045
timestamp 1676037725
transform 1 0 373244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4057
timestamp 1676037725
transform 1 0 374348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4069
timestamp 1676037725
transform 1 0 375452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4081
timestamp 1676037725
transform 1 0 376556 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4087
timestamp 1676037725
transform 1 0 377108 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4089
timestamp 1676037725
transform 1 0 377292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4101
timestamp 1676037725
transform 1 0 378396 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4113
timestamp 1676037725
transform 1 0 379500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4125
timestamp 1676037725
transform 1 0 380604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4137
timestamp 1676037725
transform 1 0 381708 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4143
timestamp 1676037725
transform 1 0 382260 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4145
timestamp 1676037725
transform 1 0 382444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4157
timestamp 1676037725
transform 1 0 383548 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_4169
timestamp 1676037725
transform 1 0 384652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_4177
timestamp 1676037725
transform 1 0 385388 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_4182
timestamp 1676037725
transform 1 0 385848 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_4198
timestamp 1676037725
transform 1 0 387320 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4201
timestamp 1676037725
transform 1 0 387596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4213
timestamp 1676037725
transform 1 0 388700 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4225
timestamp 1676037725
transform 1 0 389804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4237
timestamp 1676037725
transform 1 0 390908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4249
timestamp 1676037725
transform 1 0 392012 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4255
timestamp 1676037725
transform 1 0 392564 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4257
timestamp 1676037725
transform 1 0 392748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4269
timestamp 1676037725
transform 1 0 393852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4281
timestamp 1676037725
transform 1 0 394956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4293
timestamp 1676037725
transform 1 0 396060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4305
timestamp 1676037725
transform 1 0 397164 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4311
timestamp 1676037725
transform 1 0 397716 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4313
timestamp 1676037725
transform 1 0 397900 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4325
timestamp 1676037725
transform 1 0 399004 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_4337
timestamp 1676037725
transform 1 0 400108 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_4345
timestamp 1676037725
transform 1 0 400844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_4350
timestamp 1676037725
transform 1 0 401304 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_4366
timestamp 1676037725
transform 1 0 402776 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4369
timestamp 1676037725
transform 1 0 403052 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4381
timestamp 1676037725
transform 1 0 404156 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_4393
timestamp 1676037725
transform 1 0 405260 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_4410
timestamp 1676037725
transform 1 0 406824 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_4416
timestamp 1676037725
transform 1 0 407376 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4425
timestamp 1676037725
transform 1 0 408204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4437
timestamp 1676037725
transform 1 0 409308 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4449
timestamp 1676037725
transform 1 0 410412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4461
timestamp 1676037725
transform 1 0 411516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4473
timestamp 1676037725
transform 1 0 412620 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4479
timestamp 1676037725
transform 1 0 413172 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4481
timestamp 1676037725
transform 1 0 413356 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4493
timestamp 1676037725
transform 1 0 414460 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4505
timestamp 1676037725
transform 1 0 415564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4517
timestamp 1676037725
transform 1 0 416668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4529
timestamp 1676037725
transform 1 0 417772 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4535
timestamp 1676037725
transform 1 0 418324 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4537
timestamp 1676037725
transform 1 0 418508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4549
timestamp 1676037725
transform 1 0 419612 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4561
timestamp 1676037725
transform 1 0 420716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4573
timestamp 1676037725
transform 1 0 421820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4585
timestamp 1676037725
transform 1 0 422924 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4591
timestamp 1676037725
transform 1 0 423476 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4593
timestamp 1676037725
transform 1 0 423660 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4605
timestamp 1676037725
transform 1 0 424764 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4617
timestamp 1676037725
transform 1 0 425868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4629
timestamp 1676037725
transform 1 0 426972 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4641
timestamp 1676037725
transform 1 0 428076 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4647
timestamp 1676037725
transform 1 0 428628 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4649
timestamp 1676037725
transform 1 0 428812 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4661
timestamp 1676037725
transform 1 0 429916 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_4673
timestamp 1676037725
transform 1 0 431020 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_4681
timestamp 1676037725
transform 1 0 431756 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_4686
timestamp 1676037725
transform 1 0 432216 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_4702
timestamp 1676037725
transform 1 0 433688 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4705
timestamp 1676037725
transform 1 0 433964 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4717
timestamp 1676037725
transform 1 0 435068 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4729
timestamp 1676037725
transform 1 0 436172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4741
timestamp 1676037725
transform 1 0 437276 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4753
timestamp 1676037725
transform 1 0 438380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4759
timestamp 1676037725
transform 1 0 438932 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4761
timestamp 1676037725
transform 1 0 439116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4773
timestamp 1676037725
transform 1 0 440220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4785
timestamp 1676037725
transform 1 0 441324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4797
timestamp 1676037725
transform 1 0 442428 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4809
timestamp 1676037725
transform 1 0 443532 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4815
timestamp 1676037725
transform 1 0 444084 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4817
timestamp 1676037725
transform 1 0 444268 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4829
timestamp 1676037725
transform 1 0 445372 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_4841
timestamp 1676037725
transform 1 0 446476 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_4849
timestamp 1676037725
transform 1 0 447212 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_4853
timestamp 1676037725
transform 1 0 447580 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_4869
timestamp 1676037725
transform 1 0 449052 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4873
timestamp 1676037725
transform 1 0 449420 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4885
timestamp 1676037725
transform 1 0 450524 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4897
timestamp 1676037725
transform 1 0 451628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4909
timestamp 1676037725
transform 1 0 452732 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4921
timestamp 1676037725
transform 1 0 453836 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4927
timestamp 1676037725
transform 1 0 454388 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4929
timestamp 1676037725
transform 1 0 454572 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4941
timestamp 1676037725
transform 1 0 455676 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4953
timestamp 1676037725
transform 1 0 456780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4965
timestamp 1676037725
transform 1 0 457884 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4977
timestamp 1676037725
transform 1 0 458988 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4983
timestamp 1676037725
transform 1 0 459540 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4985
timestamp 1676037725
transform 1 0 459724 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4997
timestamp 1676037725
transform 1 0 460828 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5009
timestamp 1676037725
transform 1 0 461932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5021
timestamp 1676037725
transform 1 0 463036 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5033
timestamp 1676037725
transform 1 0 464140 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5039
timestamp 1676037725
transform 1 0 464692 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5041
timestamp 1676037725
transform 1 0 464876 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5053
timestamp 1676037725
transform 1 0 465980 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5065
timestamp 1676037725
transform 1 0 467084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5077
timestamp 1676037725
transform 1 0 468188 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5089
timestamp 1676037725
transform 1 0 469292 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5095
timestamp 1676037725
transform 1 0 469844 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5097
timestamp 1676037725
transform 1 0 470028 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5109
timestamp 1676037725
transform 1 0 471132 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5121
timestamp 1676037725
transform 1 0 472236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5133
timestamp 1676037725
transform 1 0 473340 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5145
timestamp 1676037725
transform 1 0 474444 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5151
timestamp 1676037725
transform 1 0 474996 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5153
timestamp 1676037725
transform 1 0 475180 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5165
timestamp 1676037725
transform 1 0 476284 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5177
timestamp 1676037725
transform 1 0 477388 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5189
timestamp 1676037725
transform 1 0 478492 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5201
timestamp 1676037725
transform 1 0 479596 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5207
timestamp 1676037725
transform 1 0 480148 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5209
timestamp 1676037725
transform 1 0 480332 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5221
timestamp 1676037725
transform 1 0 481436 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5233
timestamp 1676037725
transform 1 0 482540 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5245
timestamp 1676037725
transform 1 0 483644 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5257
timestamp 1676037725
transform 1 0 484748 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5263
timestamp 1676037725
transform 1 0 485300 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5265
timestamp 1676037725
transform 1 0 485484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5277
timestamp 1676037725
transform 1 0 486588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5289
timestamp 1676037725
transform 1 0 487692 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5301
timestamp 1676037725
transform 1 0 488796 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5313
timestamp 1676037725
transform 1 0 489900 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5319
timestamp 1676037725
transform 1 0 490452 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5321
timestamp 1676037725
transform 1 0 490636 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5333
timestamp 1676037725
transform 1 0 491740 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5345
timestamp 1676037725
transform 1 0 492844 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5357
timestamp 1676037725
transform 1 0 493948 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5369
timestamp 1676037725
transform 1 0 495052 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5375
timestamp 1676037725
transform 1 0 495604 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5377
timestamp 1676037725
transform 1 0 495788 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5389
timestamp 1676037725
transform 1 0 496892 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5401
timestamp 1676037725
transform 1 0 497996 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5413
timestamp 1676037725
transform 1 0 499100 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5425
timestamp 1676037725
transform 1 0 500204 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5431
timestamp 1676037725
transform 1 0 500756 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5433
timestamp 1676037725
transform 1 0 500940 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5445
timestamp 1676037725
transform 1 0 502044 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5457
timestamp 1676037725
transform 1 0 503148 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5469
timestamp 1676037725
transform 1 0 504252 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5481
timestamp 1676037725
transform 1 0 505356 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5487
timestamp 1676037725
transform 1 0 505908 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5489
timestamp 1676037725
transform 1 0 506092 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5501
timestamp 1676037725
transform 1 0 507196 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5513
timestamp 1676037725
transform 1 0 508300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5525
timestamp 1676037725
transform 1 0 509404 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5537
timestamp 1676037725
transform 1 0 510508 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5543
timestamp 1676037725
transform 1 0 511060 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5545
timestamp 1676037725
transform 1 0 511244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5557
timestamp 1676037725
transform 1 0 512348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5569
timestamp 1676037725
transform 1 0 513452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5581
timestamp 1676037725
transform 1 0 514556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5593
timestamp 1676037725
transform 1 0 515660 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5599
timestamp 1676037725
transform 1 0 516212 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5601
timestamp 1676037725
transform 1 0 516396 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5613
timestamp 1676037725
transform 1 0 517500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5625
timestamp 1676037725
transform 1 0 518604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5637
timestamp 1676037725
transform 1 0 519708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5649
timestamp 1676037725
transform 1 0 520812 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5655
timestamp 1676037725
transform 1 0 521364 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5657
timestamp 1676037725
transform 1 0 521548 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5669
timestamp 1676037725
transform 1 0 522652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5681
timestamp 1676037725
transform 1 0 523756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5693
timestamp 1676037725
transform 1 0 524860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5705
timestamp 1676037725
transform 1 0 525964 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5711
timestamp 1676037725
transform 1 0 526516 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5713
timestamp 1676037725
transform 1 0 526700 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5725
timestamp 1676037725
transform 1 0 527804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5737
timestamp 1676037725
transform 1 0 528908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5749
timestamp 1676037725
transform 1 0 530012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5761
timestamp 1676037725
transform 1 0 531116 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5767
timestamp 1676037725
transform 1 0 531668 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5769
timestamp 1676037725
transform 1 0 531852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5781
timestamp 1676037725
transform 1 0 532956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5793
timestamp 1676037725
transform 1 0 534060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5805
timestamp 1676037725
transform 1 0 535164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5817
timestamp 1676037725
transform 1 0 536268 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5823
timestamp 1676037725
transform 1 0 536820 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5825
timestamp 1676037725
transform 1 0 537004 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5837
timestamp 1676037725
transform 1 0 538108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5849
timestamp 1676037725
transform 1 0 539212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5861
timestamp 1676037725
transform 1 0 540316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5873
timestamp 1676037725
transform 1 0 541420 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5879
timestamp 1676037725
transform 1 0 541972 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5881
timestamp 1676037725
transform 1 0 542156 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5893
timestamp 1676037725
transform 1 0 543260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5905
timestamp 1676037725
transform 1 0 544364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5917
timestamp 1676037725
transform 1 0 545468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5929
timestamp 1676037725
transform 1 0 546572 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5935
timestamp 1676037725
transform 1 0 547124 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5937
timestamp 1676037725
transform 1 0 547308 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5949
timestamp 1676037725
transform 1 0 548412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5961
timestamp 1676037725
transform 1 0 549516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5973
timestamp 1676037725
transform 1 0 550620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5985
timestamp 1676037725
transform 1 0 551724 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5991
timestamp 1676037725
transform 1 0 552276 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5993
timestamp 1676037725
transform 1 0 552460 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6005
timestamp 1676037725
transform 1 0 553564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6017
timestamp 1676037725
transform 1 0 554668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6029
timestamp 1676037725
transform 1 0 555772 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6041
timestamp 1676037725
transform 1 0 556876 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6047
timestamp 1676037725
transform 1 0 557428 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6049
timestamp 1676037725
transform 1 0 557612 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6061
timestamp 1676037725
transform 1 0 558716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6073
timestamp 1676037725
transform 1 0 559820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6085
timestamp 1676037725
transform 1 0 560924 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6097
timestamp 1676037725
transform 1 0 562028 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6103
timestamp 1676037725
transform 1 0 562580 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6105
timestamp 1676037725
transform 1 0 562764 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6117
timestamp 1676037725
transform 1 0 563868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6129
timestamp 1676037725
transform 1 0 564972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6141
timestamp 1676037725
transform 1 0 566076 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6153
timestamp 1676037725
transform 1 0 567180 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6159
timestamp 1676037725
transform 1 0 567732 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6161
timestamp 1676037725
transform 1 0 567916 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6173
timestamp 1676037725
transform 1 0 569020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6185
timestamp 1676037725
transform 1 0 570124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6197
timestamp 1676037725
transform 1 0 571228 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6209
timestamp 1676037725
transform 1 0 572332 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6215
timestamp 1676037725
transform 1 0 572884 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6217
timestamp 1676037725
transform 1 0 573068 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6229
timestamp 1676037725
transform 1 0 574172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6241
timestamp 1676037725
transform 1 0 575276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6253
timestamp 1676037725
transform 1 0 576380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6265
timestamp 1676037725
transform 1 0 577484 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6271
timestamp 1676037725
transform 1 0 578036 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6273
timestamp 1676037725
transform 1 0 578220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6285
timestamp 1676037725
transform 1 0 579324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6297
timestamp 1676037725
transform 1 0 580428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6309
timestamp 1676037725
transform 1 0 581532 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6321
timestamp 1676037725
transform 1 0 582636 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6327
timestamp 1676037725
transform 1 0 583188 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6329
timestamp 1676037725
transform 1 0 583372 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6341
timestamp 1676037725
transform 1 0 584476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6353
timestamp 1676037725
transform 1 0 585580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6365
timestamp 1676037725
transform 1 0 586684 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6377
timestamp 1676037725
transform 1 0 587788 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6383
timestamp 1676037725
transform 1 0 588340 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6385
timestamp 1676037725
transform 1 0 588524 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6397
timestamp 1676037725
transform 1 0 589628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6409
timestamp 1676037725
transform 1 0 590732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6421
timestamp 1676037725
transform 1 0 591836 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6433
timestamp 1676037725
transform 1 0 592940 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6439
timestamp 1676037725
transform 1 0 593492 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6441
timestamp 1676037725
transform 1 0 593676 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6453
timestamp 1676037725
transform 1 0 594780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6465
timestamp 1676037725
transform 1 0 595884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6477
timestamp 1676037725
transform 1 0 596988 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6489
timestamp 1676037725
transform 1 0 598092 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6495
timestamp 1676037725
transform 1 0 598644 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6497
timestamp 1676037725
transform 1 0 598828 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6509
timestamp 1676037725
transform 1 0 599932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6521
timestamp 1676037725
transform 1 0 601036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6533
timestamp 1676037725
transform 1 0 602140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6545
timestamp 1676037725
transform 1 0 603244 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6551
timestamp 1676037725
transform 1 0 603796 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6553
timestamp 1676037725
transform 1 0 603980 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6565
timestamp 1676037725
transform 1 0 605084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6577
timestamp 1676037725
transform 1 0 606188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6589
timestamp 1676037725
transform 1 0 607292 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6601
timestamp 1676037725
transform 1 0 608396 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6607
timestamp 1676037725
transform 1 0 608948 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6609
timestamp 1676037725
transform 1 0 609132 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6621
timestamp 1676037725
transform 1 0 610236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6633
timestamp 1676037725
transform 1 0 611340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6645
timestamp 1676037725
transform 1 0 612444 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6657
timestamp 1676037725
transform 1 0 613548 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6663
timestamp 1676037725
transform 1 0 614100 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6665
timestamp 1676037725
transform 1 0 614284 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6677
timestamp 1676037725
transform 1 0 615388 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6689
timestamp 1676037725
transform 1 0 616492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6701
timestamp 1676037725
transform 1 0 617596 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6713
timestamp 1676037725
transform 1 0 618700 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6719
timestamp 1676037725
transform 1 0 619252 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6721
timestamp 1676037725
transform 1 0 619436 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6733
timestamp 1676037725
transform 1 0 620540 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6745
timestamp 1676037725
transform 1 0 621644 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6757
timestamp 1676037725
transform 1 0 622748 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6769
timestamp 1676037725
transform 1 0 623852 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6775
timestamp 1676037725
transform 1 0 624404 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6777
timestamp 1676037725
transform 1 0 624588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6789
timestamp 1676037725
transform 1 0 625692 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6801
timestamp 1676037725
transform 1 0 626796 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6813
timestamp 1676037725
transform 1 0 627900 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6825
timestamp 1676037725
transform 1 0 629004 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6831
timestamp 1676037725
transform 1 0 629556 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6833
timestamp 1676037725
transform 1 0 629740 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6845
timestamp 1676037725
transform 1 0 630844 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6857
timestamp 1676037725
transform 1 0 631948 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6869
timestamp 1676037725
transform 1 0 633052 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6881
timestamp 1676037725
transform 1 0 634156 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6887
timestamp 1676037725
transform 1 0 634708 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6889
timestamp 1676037725
transform 1 0 634892 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6901
timestamp 1676037725
transform 1 0 635996 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6913
timestamp 1676037725
transform 1 0 637100 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6925
timestamp 1676037725
transform 1 0 638204 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6937
timestamp 1676037725
transform 1 0 639308 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6943
timestamp 1676037725
transform 1 0 639860 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6945
timestamp 1676037725
transform 1 0 640044 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6957
timestamp 1676037725
transform 1 0 641148 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6969
timestamp 1676037725
transform 1 0 642252 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6981
timestamp 1676037725
transform 1 0 643356 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6993
timestamp 1676037725
transform 1 0 644460 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6999
timestamp 1676037725
transform 1 0 645012 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7001
timestamp 1676037725
transform 1 0 645196 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7013
timestamp 1676037725
transform 1 0 646300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7025
timestamp 1676037725
transform 1 0 647404 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7037
timestamp 1676037725
transform 1 0 648508 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1676037725
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1676037725
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1676037725
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1676037725
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1676037725
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1676037725
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1676037725
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1676037725
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1676037725
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1676037725
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1676037725
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1676037725
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1676037725
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1676037725
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1676037725
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1676037725
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1676037725
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1676037725
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1676037725
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1676037725
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1676037725
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1676037725
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1676037725
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1676037725
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1676037725
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1676037725
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1676037725
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1676037725
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1676037725
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1676037725
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1676037725
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_725
timestamp 1676037725
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_737
timestamp 1676037725
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 1676037725
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1676037725
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1676037725
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1676037725
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_781
timestamp 1676037725
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_793
timestamp 1676037725
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1676037725
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1676037725
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_813
timestamp 1676037725
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_825
timestamp 1676037725
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_837
timestamp 1676037725
transform 1 0 78108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_849
timestamp 1676037725
transform 1 0 79212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_861
timestamp 1676037725
transform 1 0 80316 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_867
timestamp 1676037725
transform 1 0 80868 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_869
timestamp 1676037725
transform 1 0 81052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_881
timestamp 1676037725
transform 1 0 82156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_893
timestamp 1676037725
transform 1 0 83260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_905
timestamp 1676037725
transform 1 0 84364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_917
timestamp 1676037725
transform 1 0 85468 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_923
timestamp 1676037725
transform 1 0 86020 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_925
timestamp 1676037725
transform 1 0 86204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_937
timestamp 1676037725
transform 1 0 87308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_949
timestamp 1676037725
transform 1 0 88412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_961
timestamp 1676037725
transform 1 0 89516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_973
timestamp 1676037725
transform 1 0 90620 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_979
timestamp 1676037725
transform 1 0 91172 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_981
timestamp 1676037725
transform 1 0 91356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_993
timestamp 1676037725
transform 1 0 92460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1005
timestamp 1676037725
transform 1 0 93564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1017
timestamp 1676037725
transform 1 0 94668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1029
timestamp 1676037725
transform 1 0 95772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1035
timestamp 1676037725
transform 1 0 96324 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1037
timestamp 1676037725
transform 1 0 96508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1049
timestamp 1676037725
transform 1 0 97612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1061
timestamp 1676037725
transform 1 0 98716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1073
timestamp 1676037725
transform 1 0 99820 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1085
timestamp 1676037725
transform 1 0 100924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1091
timestamp 1676037725
transform 1 0 101476 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1093
timestamp 1676037725
transform 1 0 101660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1105
timestamp 1676037725
transform 1 0 102764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1117
timestamp 1676037725
transform 1 0 103868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1129
timestamp 1676037725
transform 1 0 104972 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1141
timestamp 1676037725
transform 1 0 106076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1147
timestamp 1676037725
transform 1 0 106628 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1149
timestamp 1676037725
transform 1 0 106812 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1161
timestamp 1676037725
transform 1 0 107916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1173
timestamp 1676037725
transform 1 0 109020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1185
timestamp 1676037725
transform 1 0 110124 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1197
timestamp 1676037725
transform 1 0 111228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1203
timestamp 1676037725
transform 1 0 111780 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1205
timestamp 1676037725
transform 1 0 111964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1217
timestamp 1676037725
transform 1 0 113068 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1229
timestamp 1676037725
transform 1 0 114172 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1240
timestamp 1676037725
transform 1 0 115184 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1246
timestamp 1676037725
transform 1 0 115736 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1258
timestamp 1676037725
transform 1 0 116840 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1261
timestamp 1676037725
transform 1 0 117116 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1273
timestamp 1676037725
transform 1 0 118220 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1285
timestamp 1676037725
transform 1 0 119324 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1297
timestamp 1676037725
transform 1 0 120428 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1309
timestamp 1676037725
transform 1 0 121532 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1315
timestamp 1676037725
transform 1 0 122084 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1317
timestamp 1676037725
transform 1 0 122268 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1321
timestamp 1676037725
transform 1 0 122636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1333
timestamp 1676037725
transform 1 0 123740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1345
timestamp 1676037725
transform 1 0 124844 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1357
timestamp 1676037725
transform 1 0 125948 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_1369
timestamp 1676037725
transform 1 0 127052 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1373
timestamp 1676037725
transform 1 0 127420 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1385
timestamp 1676037725
transform 1 0 128524 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1397
timestamp 1676037725
transform 1 0 129628 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1409
timestamp 1676037725
transform 1 0 130732 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1421
timestamp 1676037725
transform 1 0 131836 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1427
timestamp 1676037725
transform 1 0 132388 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1429
timestamp 1676037725
transform 1 0 132572 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1441
timestamp 1676037725
transform 1 0 133676 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1453
timestamp 1676037725
transform 1 0 134780 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1465
timestamp 1676037725
transform 1 0 135884 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1477
timestamp 1676037725
transform 1 0 136988 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1483
timestamp 1676037725
transform 1 0 137540 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1485
timestamp 1676037725
transform 1 0 137724 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1497
timestamp 1676037725
transform 1 0 138828 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1509
timestamp 1676037725
transform 1 0 139932 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1521
timestamp 1676037725
transform 1 0 141036 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1533
timestamp 1676037725
transform 1 0 142140 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1539
timestamp 1676037725
transform 1 0 142692 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1541
timestamp 1676037725
transform 1 0 142876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1553
timestamp 1676037725
transform 1 0 143980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1565
timestamp 1676037725
transform 1 0 145084 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1577
timestamp 1676037725
transform 1 0 146188 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1589
timestamp 1676037725
transform 1 0 147292 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1595
timestamp 1676037725
transform 1 0 147844 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1597
timestamp 1676037725
transform 1 0 148028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1609
timestamp 1676037725
transform 1 0 149132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1621
timestamp 1676037725
transform 1 0 150236 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1633
timestamp 1676037725
transform 1 0 151340 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1645
timestamp 1676037725
transform 1 0 152444 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1651
timestamp 1676037725
transform 1 0 152996 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1653
timestamp 1676037725
transform 1 0 153180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1665
timestamp 1676037725
transform 1 0 154284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1677
timestamp 1676037725
transform 1 0 155388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1689
timestamp 1676037725
transform 1 0 156492 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1693
timestamp 1676037725
transform 1 0 156860 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1706
timestamp 1676037725
transform 1 0 158056 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1709
timestamp 1676037725
transform 1 0 158332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1721
timestamp 1676037725
transform 1 0 159436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1733
timestamp 1676037725
transform 1 0 160540 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1745
timestamp 1676037725
transform 1 0 161644 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1757
timestamp 1676037725
transform 1 0 162748 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1763
timestamp 1676037725
transform 1 0 163300 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1765
timestamp 1676037725
transform 1 0 163484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1777
timestamp 1676037725
transform 1 0 164588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1789
timestamp 1676037725
transform 1 0 165692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1801
timestamp 1676037725
transform 1 0 166796 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1813
timestamp 1676037725
transform 1 0 167900 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1819
timestamp 1676037725
transform 1 0 168452 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1821
timestamp 1676037725
transform 1 0 168636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1833
timestamp 1676037725
transform 1 0 169740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1845
timestamp 1676037725
transform 1 0 170844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1857
timestamp 1676037725
transform 1 0 171948 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1860
timestamp 1676037725
transform 1 0 172224 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_1873
timestamp 1676037725
transform 1 0 173420 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1877
timestamp 1676037725
transform 1 0 173788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1889
timestamp 1676037725
transform 1 0 174892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1901
timestamp 1676037725
transform 1 0 175996 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1913
timestamp 1676037725
transform 1 0 177100 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1925
timestamp 1676037725
transform 1 0 178204 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1931
timestamp 1676037725
transform 1 0 178756 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1933
timestamp 1676037725
transform 1 0 178940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1945
timestamp 1676037725
transform 1 0 180044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1957
timestamp 1676037725
transform 1 0 181148 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1969
timestamp 1676037725
transform 1 0 182252 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1981
timestamp 1676037725
transform 1 0 183356 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1987
timestamp 1676037725
transform 1 0 183908 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1989
timestamp 1676037725
transform 1 0 184092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2001
timestamp 1676037725
transform 1 0 185196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2013
timestamp 1676037725
transform 1 0 186300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2025
timestamp 1676037725
transform 1 0 187404 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2037
timestamp 1676037725
transform 1 0 188508 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2043
timestamp 1676037725
transform 1 0 189060 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2045
timestamp 1676037725
transform 1 0 189244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2057
timestamp 1676037725
transform 1 0 190348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2069
timestamp 1676037725
transform 1 0 191452 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2081
timestamp 1676037725
transform 1 0 192556 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2093
timestamp 1676037725
transform 1 0 193660 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2099
timestamp 1676037725
transform 1 0 194212 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2101
timestamp 1676037725
transform 1 0 194396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2113
timestamp 1676037725
transform 1 0 195500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2125
timestamp 1676037725
transform 1 0 196604 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2137
timestamp 1676037725
transform 1 0 197708 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2149
timestamp 1676037725
transform 1 0 198812 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2155
timestamp 1676037725
transform 1 0 199364 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2157
timestamp 1676037725
transform 1 0 199548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2169
timestamp 1676037725
transform 1 0 200652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2181
timestamp 1676037725
transform 1 0 201756 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2193
timestamp 1676037725
transform 1 0 202860 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2205
timestamp 1676037725
transform 1 0 203964 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2211
timestamp 1676037725
transform 1 0 204516 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2213
timestamp 1676037725
transform 1 0 204700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2225
timestamp 1676037725
transform 1 0 205804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2237
timestamp 1676037725
transform 1 0 206908 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2249
timestamp 1676037725
transform 1 0 208012 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2261
timestamp 1676037725
transform 1 0 209116 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2267
timestamp 1676037725
transform 1 0 209668 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2269
timestamp 1676037725
transform 1 0 209852 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_2281
timestamp 1676037725
transform 1 0 210956 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2285
timestamp 1676037725
transform 1 0 211324 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_2295
timestamp 1676037725
transform 1 0 212244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_2301
timestamp 1676037725
transform 1 0 212796 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2309
timestamp 1676037725
transform 1 0 213532 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2312
timestamp 1676037725
transform 1 0 213808 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_2325
timestamp 1676037725
transform 1 0 215004 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2329
timestamp 1676037725
transform 1 0 215372 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2341
timestamp 1676037725
transform 1 0 216476 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2353
timestamp 1676037725
transform 1 0 217580 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2365
timestamp 1676037725
transform 1 0 218684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_2377
timestamp 1676037725
transform 1 0 219788 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2381
timestamp 1676037725
transform 1 0 220156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2393
timestamp 1676037725
transform 1 0 221260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2405
timestamp 1676037725
transform 1 0 222364 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2417
timestamp 1676037725
transform 1 0 223468 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2429
timestamp 1676037725
transform 1 0 224572 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2435
timestamp 1676037725
transform 1 0 225124 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2437
timestamp 1676037725
transform 1 0 225308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2449
timestamp 1676037725
transform 1 0 226412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2461
timestamp 1676037725
transform 1 0 227516 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2473
timestamp 1676037725
transform 1 0 228620 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2485
timestamp 1676037725
transform 1 0 229724 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2491
timestamp 1676037725
transform 1 0 230276 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2493
timestamp 1676037725
transform 1 0 230460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2505
timestamp 1676037725
transform 1 0 231564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2517
timestamp 1676037725
transform 1 0 232668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2529
timestamp 1676037725
transform 1 0 233772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2541
timestamp 1676037725
transform 1 0 234876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2547
timestamp 1676037725
transform 1 0 235428 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2549
timestamp 1676037725
transform 1 0 235612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2561
timestamp 1676037725
transform 1 0 236716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2573
timestamp 1676037725
transform 1 0 237820 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2585
timestamp 1676037725
transform 1 0 238924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2597
timestamp 1676037725
transform 1 0 240028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2603
timestamp 1676037725
transform 1 0 240580 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2605
timestamp 1676037725
transform 1 0 240764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2617
timestamp 1676037725
transform 1 0 241868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2629
timestamp 1676037725
transform 1 0 242972 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2641
timestamp 1676037725
transform 1 0 244076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2653
timestamp 1676037725
transform 1 0 245180 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2659
timestamp 1676037725
transform 1 0 245732 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2661
timestamp 1676037725
transform 1 0 245916 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2673
timestamp 1676037725
transform 1 0 247020 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_2681
timestamp 1676037725
transform 1 0 247756 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2697
timestamp 1676037725
transform 1 0 249228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2709
timestamp 1676037725
transform 1 0 250332 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2715
timestamp 1676037725
transform 1 0 250884 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2717
timestamp 1676037725
transform 1 0 251068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2729
timestamp 1676037725
transform 1 0 252172 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2741
timestamp 1676037725
transform 1 0 253276 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2753
timestamp 1676037725
transform 1 0 254380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2765
timestamp 1676037725
transform 1 0 255484 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2771
timestamp 1676037725
transform 1 0 256036 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2773
timestamp 1676037725
transform 1 0 256220 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2785
timestamp 1676037725
transform 1 0 257324 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2797
timestamp 1676037725
transform 1 0 258428 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2809
timestamp 1676037725
transform 1 0 259532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2821
timestamp 1676037725
transform 1 0 260636 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2827
timestamp 1676037725
transform 1 0 261188 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2829
timestamp 1676037725
transform 1 0 261372 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_2841
timestamp 1676037725
transform 1 0 262476 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2845
timestamp 1676037725
transform 1 0 262844 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_2848
timestamp 1676037725
transform 1 0 263120 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2864
timestamp 1676037725
transform 1 0 264592 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_2876
timestamp 1676037725
transform 1 0 265696 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2885
timestamp 1676037725
transform 1 0 266524 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2897
timestamp 1676037725
transform 1 0 267628 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2909
timestamp 1676037725
transform 1 0 268732 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2921
timestamp 1676037725
transform 1 0 269836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2933
timestamp 1676037725
transform 1 0 270940 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2939
timestamp 1676037725
transform 1 0 271492 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2941
timestamp 1676037725
transform 1 0 271676 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2953
timestamp 1676037725
transform 1 0 272780 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2965
timestamp 1676037725
transform 1 0 273884 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2977
timestamp 1676037725
transform 1 0 274988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2989
timestamp 1676037725
transform 1 0 276092 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2995
timestamp 1676037725
transform 1 0 276644 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2997
timestamp 1676037725
transform 1 0 276828 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3009
timestamp 1676037725
transform 1 0 277932 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3021
timestamp 1676037725
transform 1 0 279036 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3033
timestamp 1676037725
transform 1 0 280140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3045
timestamp 1676037725
transform 1 0 281244 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3051
timestamp 1676037725
transform 1 0 281796 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3053
timestamp 1676037725
transform 1 0 281980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3065
timestamp 1676037725
transform 1 0 283084 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3077
timestamp 1676037725
transform 1 0 284188 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3089
timestamp 1676037725
transform 1 0 285292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3101
timestamp 1676037725
transform 1 0 286396 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3107
timestamp 1676037725
transform 1 0 286948 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3109
timestamp 1676037725
transform 1 0 287132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3121
timestamp 1676037725
transform 1 0 288236 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3133
timestamp 1676037725
transform 1 0 289340 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3145
timestamp 1676037725
transform 1 0 290444 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3157
timestamp 1676037725
transform 1 0 291548 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3163
timestamp 1676037725
transform 1 0 292100 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3165
timestamp 1676037725
transform 1 0 292284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3177
timestamp 1676037725
transform 1 0 293388 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3182
timestamp 1676037725
transform 1 0 293848 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3198
timestamp 1676037725
transform 1 0 295320 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3210
timestamp 1676037725
transform 1 0 296424 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3218
timestamp 1676037725
transform 1 0 297160 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3221
timestamp 1676037725
transform 1 0 297436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3233
timestamp 1676037725
transform 1 0 298540 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3245
timestamp 1676037725
transform 1 0 299644 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3257
timestamp 1676037725
transform 1 0 300748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3269
timestamp 1676037725
transform 1 0 301852 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3275
timestamp 1676037725
transform 1 0 302404 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3277
timestamp 1676037725
transform 1 0 302588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3289
timestamp 1676037725
transform 1 0 303692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3301
timestamp 1676037725
transform 1 0 304796 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3313
timestamp 1676037725
transform 1 0 305900 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3325
timestamp 1676037725
transform 1 0 307004 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3331
timestamp 1676037725
transform 1 0 307556 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3333
timestamp 1676037725
transform 1 0 307740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3345
timestamp 1676037725
transform 1 0 308844 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3353
timestamp 1676037725
transform 1 0 309580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3368
timestamp 1676037725
transform 1 0 310960 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3376
timestamp 1676037725
transform 1 0 311696 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3379
timestamp 1676037725
transform 1 0 311972 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3387
timestamp 1676037725
transform 1 0 312708 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3389
timestamp 1676037725
transform 1 0 312892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3401
timestamp 1676037725
transform 1 0 313996 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3413
timestamp 1676037725
transform 1 0 315100 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3425
timestamp 1676037725
transform 1 0 316204 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3437
timestamp 1676037725
transform 1 0 317308 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3443
timestamp 1676037725
transform 1 0 317860 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3445
timestamp 1676037725
transform 1 0 318044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3457
timestamp 1676037725
transform 1 0 319148 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3469
timestamp 1676037725
transform 1 0 320252 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3481
timestamp 1676037725
transform 1 0 321356 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3493
timestamp 1676037725
transform 1 0 322460 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3499
timestamp 1676037725
transform 1 0 323012 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3501
timestamp 1676037725
transform 1 0 323196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3513
timestamp 1676037725
transform 1 0 324300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3525
timestamp 1676037725
transform 1 0 325404 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3537
timestamp 1676037725
transform 1 0 326508 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3549
timestamp 1676037725
transform 1 0 327612 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3555
timestamp 1676037725
transform 1 0 328164 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3557
timestamp 1676037725
transform 1 0 328348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3569
timestamp 1676037725
transform 1 0 329452 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3581
timestamp 1676037725
transform 1 0 330556 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3593
timestamp 1676037725
transform 1 0 331660 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3605
timestamp 1676037725
transform 1 0 332764 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3611
timestamp 1676037725
transform 1 0 333316 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3613
timestamp 1676037725
transform 1 0 333500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3625
timestamp 1676037725
transform 1 0 334604 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3637
timestamp 1676037725
transform 1 0 335708 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3649
timestamp 1676037725
transform 1 0 336812 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3661
timestamp 1676037725
transform 1 0 337916 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3667
timestamp 1676037725
transform 1 0 338468 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3669
timestamp 1676037725
transform 1 0 338652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3681
timestamp 1676037725
transform 1 0 339756 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3693
timestamp 1676037725
transform 1 0 340860 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3705
timestamp 1676037725
transform 1 0 341964 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3717
timestamp 1676037725
transform 1 0 343068 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3723
timestamp 1676037725
transform 1 0 343620 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3725
timestamp 1676037725
transform 1 0 343804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3737
timestamp 1676037725
transform 1 0 344908 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3749
timestamp 1676037725
transform 1 0 346012 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3761
timestamp 1676037725
transform 1 0 347116 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3773
timestamp 1676037725
transform 1 0 348220 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3779
timestamp 1676037725
transform 1 0 348772 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3781
timestamp 1676037725
transform 1 0 348956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3793
timestamp 1676037725
transform 1 0 350060 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3805
timestamp 1676037725
transform 1 0 351164 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3817
timestamp 1676037725
transform 1 0 352268 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3829
timestamp 1676037725
transform 1 0 353372 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3835
timestamp 1676037725
transform 1 0 353924 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3837
timestamp 1676037725
transform 1 0 354108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3849
timestamp 1676037725
transform 1 0 355212 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3861
timestamp 1676037725
transform 1 0 356316 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3873
timestamp 1676037725
transform 1 0 357420 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3885
timestamp 1676037725
transform 1 0 358524 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3891
timestamp 1676037725
transform 1 0 359076 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3893
timestamp 1676037725
transform 1 0 359260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3905
timestamp 1676037725
transform 1 0 360364 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3917
timestamp 1676037725
transform 1 0 361468 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3929
timestamp 1676037725
transform 1 0 362572 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3941
timestamp 1676037725
transform 1 0 363676 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3947
timestamp 1676037725
transform 1 0 364228 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3949
timestamp 1676037725
transform 1 0 364412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3961
timestamp 1676037725
transform 1 0 365516 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3973
timestamp 1676037725
transform 1 0 366620 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3985
timestamp 1676037725
transform 1 0 367724 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3997
timestamp 1676037725
transform 1 0 368828 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4003
timestamp 1676037725
transform 1 0 369380 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4005
timestamp 1676037725
transform 1 0 369564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4017
timestamp 1676037725
transform 1 0 370668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4029
timestamp 1676037725
transform 1 0 371772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4041
timestamp 1676037725
transform 1 0 372876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4053
timestamp 1676037725
transform 1 0 373980 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4059
timestamp 1676037725
transform 1 0 374532 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4061
timestamp 1676037725
transform 1 0 374716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4073
timestamp 1676037725
transform 1 0 375820 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4085
timestamp 1676037725
transform 1 0 376924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4097
timestamp 1676037725
transform 1 0 378028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4109
timestamp 1676037725
transform 1 0 379132 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4115
timestamp 1676037725
transform 1 0 379684 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4117
timestamp 1676037725
transform 1 0 379868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4129
timestamp 1676037725
transform 1 0 380972 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4141
timestamp 1676037725
transform 1 0 382076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4153
timestamp 1676037725
transform 1 0 383180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4165
timestamp 1676037725
transform 1 0 384284 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4171
timestamp 1676037725
transform 1 0 384836 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4173
timestamp 1676037725
transform 1 0 385020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4185
timestamp 1676037725
transform 1 0 386124 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4197
timestamp 1676037725
transform 1 0 387228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4209
timestamp 1676037725
transform 1 0 388332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4221
timestamp 1676037725
transform 1 0 389436 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4227
timestamp 1676037725
transform 1 0 389988 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4229
timestamp 1676037725
transform 1 0 390172 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4241
timestamp 1676037725
transform 1 0 391276 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4253
timestamp 1676037725
transform 1 0 392380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4265
timestamp 1676037725
transform 1 0 393484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4277
timestamp 1676037725
transform 1 0 394588 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4283
timestamp 1676037725
transform 1 0 395140 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4285
timestamp 1676037725
transform 1 0 395324 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4297
timestamp 1676037725
transform 1 0 396428 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4309
timestamp 1676037725
transform 1 0 397532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4321
timestamp 1676037725
transform 1 0 398636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4333
timestamp 1676037725
transform 1 0 399740 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4339
timestamp 1676037725
transform 1 0 400292 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4341
timestamp 1676037725
transform 1 0 400476 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4353
timestamp 1676037725
transform 1 0 401580 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4365
timestamp 1676037725
transform 1 0 402684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4377
timestamp 1676037725
transform 1 0 403788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4389
timestamp 1676037725
transform 1 0 404892 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4395
timestamp 1676037725
transform 1 0 405444 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4397
timestamp 1676037725
transform 1 0 405628 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4409
timestamp 1676037725
transform 1 0 406732 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4421
timestamp 1676037725
transform 1 0 407836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4433
timestamp 1676037725
transform 1 0 408940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4445
timestamp 1676037725
transform 1 0 410044 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4451
timestamp 1676037725
transform 1 0 410596 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4453
timestamp 1676037725
transform 1 0 410780 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4465
timestamp 1676037725
transform 1 0 411884 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4477
timestamp 1676037725
transform 1 0 412988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4489
timestamp 1676037725
transform 1 0 414092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4501
timestamp 1676037725
transform 1 0 415196 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4507
timestamp 1676037725
transform 1 0 415748 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4509
timestamp 1676037725
transform 1 0 415932 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4521
timestamp 1676037725
transform 1 0 417036 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4533
timestamp 1676037725
transform 1 0 418140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4545
timestamp 1676037725
transform 1 0 419244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4557
timestamp 1676037725
transform 1 0 420348 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4563
timestamp 1676037725
transform 1 0 420900 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4565
timestamp 1676037725
transform 1 0 421084 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4577
timestamp 1676037725
transform 1 0 422188 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4589
timestamp 1676037725
transform 1 0 423292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4601
timestamp 1676037725
transform 1 0 424396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4613
timestamp 1676037725
transform 1 0 425500 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4619
timestamp 1676037725
transform 1 0 426052 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4621
timestamp 1676037725
transform 1 0 426236 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4633
timestamp 1676037725
transform 1 0 427340 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4645
timestamp 1676037725
transform 1 0 428444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4657
timestamp 1676037725
transform 1 0 429548 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4669
timestamp 1676037725
transform 1 0 430652 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4675
timestamp 1676037725
transform 1 0 431204 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4677
timestamp 1676037725
transform 1 0 431388 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4689
timestamp 1676037725
transform 1 0 432492 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4701
timestamp 1676037725
transform 1 0 433596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4713
timestamp 1676037725
transform 1 0 434700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4725
timestamp 1676037725
transform 1 0 435804 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4731
timestamp 1676037725
transform 1 0 436356 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4733
timestamp 1676037725
transform 1 0 436540 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4745
timestamp 1676037725
transform 1 0 437644 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4757
timestamp 1676037725
transform 1 0 438748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4769
timestamp 1676037725
transform 1 0 439852 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4781
timestamp 1676037725
transform 1 0 440956 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4787
timestamp 1676037725
transform 1 0 441508 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4789
timestamp 1676037725
transform 1 0 441692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4801
timestamp 1676037725
transform 1 0 442796 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4813
timestamp 1676037725
transform 1 0 443900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4825
timestamp 1676037725
transform 1 0 445004 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4837
timestamp 1676037725
transform 1 0 446108 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4843
timestamp 1676037725
transform 1 0 446660 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4845
timestamp 1676037725
transform 1 0 446844 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4857
timestamp 1676037725
transform 1 0 447948 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4869
timestamp 1676037725
transform 1 0 449052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4881
timestamp 1676037725
transform 1 0 450156 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4893
timestamp 1676037725
transform 1 0 451260 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4899
timestamp 1676037725
transform 1 0 451812 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4901
timestamp 1676037725
transform 1 0 451996 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4913
timestamp 1676037725
transform 1 0 453100 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4925
timestamp 1676037725
transform 1 0 454204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4937
timestamp 1676037725
transform 1 0 455308 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4949
timestamp 1676037725
transform 1 0 456412 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4955
timestamp 1676037725
transform 1 0 456964 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4957
timestamp 1676037725
transform 1 0 457148 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4969
timestamp 1676037725
transform 1 0 458252 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4981
timestamp 1676037725
transform 1 0 459356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4993
timestamp 1676037725
transform 1 0 460460 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5005
timestamp 1676037725
transform 1 0 461564 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5011
timestamp 1676037725
transform 1 0 462116 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5013
timestamp 1676037725
transform 1 0 462300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5025
timestamp 1676037725
transform 1 0 463404 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5037
timestamp 1676037725
transform 1 0 464508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5049
timestamp 1676037725
transform 1 0 465612 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5061
timestamp 1676037725
transform 1 0 466716 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5067
timestamp 1676037725
transform 1 0 467268 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5069
timestamp 1676037725
transform 1 0 467452 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5081
timestamp 1676037725
transform 1 0 468556 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5093
timestamp 1676037725
transform 1 0 469660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5105
timestamp 1676037725
transform 1 0 470764 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5117
timestamp 1676037725
transform 1 0 471868 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5123
timestamp 1676037725
transform 1 0 472420 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5125
timestamp 1676037725
transform 1 0 472604 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5137
timestamp 1676037725
transform 1 0 473708 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5149
timestamp 1676037725
transform 1 0 474812 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5161
timestamp 1676037725
transform 1 0 475916 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5173
timestamp 1676037725
transform 1 0 477020 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5179
timestamp 1676037725
transform 1 0 477572 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5181
timestamp 1676037725
transform 1 0 477756 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5193
timestamp 1676037725
transform 1 0 478860 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5205
timestamp 1676037725
transform 1 0 479964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5217
timestamp 1676037725
transform 1 0 481068 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5229
timestamp 1676037725
transform 1 0 482172 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5235
timestamp 1676037725
transform 1 0 482724 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5237
timestamp 1676037725
transform 1 0 482908 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5249
timestamp 1676037725
transform 1 0 484012 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5261
timestamp 1676037725
transform 1 0 485116 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5273
timestamp 1676037725
transform 1 0 486220 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5285
timestamp 1676037725
transform 1 0 487324 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5291
timestamp 1676037725
transform 1 0 487876 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5293
timestamp 1676037725
transform 1 0 488060 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5305
timestamp 1676037725
transform 1 0 489164 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5317
timestamp 1676037725
transform 1 0 490268 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5329
timestamp 1676037725
transform 1 0 491372 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5341
timestamp 1676037725
transform 1 0 492476 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5347
timestamp 1676037725
transform 1 0 493028 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5349
timestamp 1676037725
transform 1 0 493212 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5361
timestamp 1676037725
transform 1 0 494316 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5373
timestamp 1676037725
transform 1 0 495420 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5385
timestamp 1676037725
transform 1 0 496524 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5397
timestamp 1676037725
transform 1 0 497628 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5403
timestamp 1676037725
transform 1 0 498180 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5405
timestamp 1676037725
transform 1 0 498364 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5417
timestamp 1676037725
transform 1 0 499468 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5429
timestamp 1676037725
transform 1 0 500572 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5441
timestamp 1676037725
transform 1 0 501676 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5453
timestamp 1676037725
transform 1 0 502780 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5459
timestamp 1676037725
transform 1 0 503332 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5461
timestamp 1676037725
transform 1 0 503516 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5473
timestamp 1676037725
transform 1 0 504620 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5485
timestamp 1676037725
transform 1 0 505724 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5497
timestamp 1676037725
transform 1 0 506828 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5509
timestamp 1676037725
transform 1 0 507932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5515
timestamp 1676037725
transform 1 0 508484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5517
timestamp 1676037725
transform 1 0 508668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5529
timestamp 1676037725
transform 1 0 509772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5541
timestamp 1676037725
transform 1 0 510876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5553
timestamp 1676037725
transform 1 0 511980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5565
timestamp 1676037725
transform 1 0 513084 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5571
timestamp 1676037725
transform 1 0 513636 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5573
timestamp 1676037725
transform 1 0 513820 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5585
timestamp 1676037725
transform 1 0 514924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5597
timestamp 1676037725
transform 1 0 516028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5609
timestamp 1676037725
transform 1 0 517132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5621
timestamp 1676037725
transform 1 0 518236 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5627
timestamp 1676037725
transform 1 0 518788 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5629
timestamp 1676037725
transform 1 0 518972 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5641
timestamp 1676037725
transform 1 0 520076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5653
timestamp 1676037725
transform 1 0 521180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5665
timestamp 1676037725
transform 1 0 522284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5677
timestamp 1676037725
transform 1 0 523388 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5683
timestamp 1676037725
transform 1 0 523940 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5685
timestamp 1676037725
transform 1 0 524124 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5697
timestamp 1676037725
transform 1 0 525228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5709
timestamp 1676037725
transform 1 0 526332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5721
timestamp 1676037725
transform 1 0 527436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5733
timestamp 1676037725
transform 1 0 528540 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5739
timestamp 1676037725
transform 1 0 529092 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5741
timestamp 1676037725
transform 1 0 529276 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5753
timestamp 1676037725
transform 1 0 530380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5765
timestamp 1676037725
transform 1 0 531484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5777
timestamp 1676037725
transform 1 0 532588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5789
timestamp 1676037725
transform 1 0 533692 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5795
timestamp 1676037725
transform 1 0 534244 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5797
timestamp 1676037725
transform 1 0 534428 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5809
timestamp 1676037725
transform 1 0 535532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5821
timestamp 1676037725
transform 1 0 536636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5833
timestamp 1676037725
transform 1 0 537740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5845
timestamp 1676037725
transform 1 0 538844 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5851
timestamp 1676037725
transform 1 0 539396 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5853
timestamp 1676037725
transform 1 0 539580 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5865
timestamp 1676037725
transform 1 0 540684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5877
timestamp 1676037725
transform 1 0 541788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5889
timestamp 1676037725
transform 1 0 542892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5901
timestamp 1676037725
transform 1 0 543996 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5907
timestamp 1676037725
transform 1 0 544548 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5909
timestamp 1676037725
transform 1 0 544732 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5921
timestamp 1676037725
transform 1 0 545836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5933
timestamp 1676037725
transform 1 0 546940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5945
timestamp 1676037725
transform 1 0 548044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5957
timestamp 1676037725
transform 1 0 549148 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5963
timestamp 1676037725
transform 1 0 549700 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5965
timestamp 1676037725
transform 1 0 549884 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5977
timestamp 1676037725
transform 1 0 550988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5989
timestamp 1676037725
transform 1 0 552092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6001
timestamp 1676037725
transform 1 0 553196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6013
timestamp 1676037725
transform 1 0 554300 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6019
timestamp 1676037725
transform 1 0 554852 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6021
timestamp 1676037725
transform 1 0 555036 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6033
timestamp 1676037725
transform 1 0 556140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6045
timestamp 1676037725
transform 1 0 557244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6057
timestamp 1676037725
transform 1 0 558348 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6069
timestamp 1676037725
transform 1 0 559452 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6075
timestamp 1676037725
transform 1 0 560004 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6077
timestamp 1676037725
transform 1 0 560188 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6089
timestamp 1676037725
transform 1 0 561292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6101
timestamp 1676037725
transform 1 0 562396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6113
timestamp 1676037725
transform 1 0 563500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6125
timestamp 1676037725
transform 1 0 564604 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6131
timestamp 1676037725
transform 1 0 565156 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6133
timestamp 1676037725
transform 1 0 565340 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6145
timestamp 1676037725
transform 1 0 566444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6157
timestamp 1676037725
transform 1 0 567548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6169
timestamp 1676037725
transform 1 0 568652 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6181
timestamp 1676037725
transform 1 0 569756 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6187
timestamp 1676037725
transform 1 0 570308 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6189
timestamp 1676037725
transform 1 0 570492 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6201
timestamp 1676037725
transform 1 0 571596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6213
timestamp 1676037725
transform 1 0 572700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6225
timestamp 1676037725
transform 1 0 573804 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6237
timestamp 1676037725
transform 1 0 574908 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6243
timestamp 1676037725
transform 1 0 575460 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6245
timestamp 1676037725
transform 1 0 575644 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6257
timestamp 1676037725
transform 1 0 576748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6269
timestamp 1676037725
transform 1 0 577852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6281
timestamp 1676037725
transform 1 0 578956 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6293
timestamp 1676037725
transform 1 0 580060 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6299
timestamp 1676037725
transform 1 0 580612 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6301
timestamp 1676037725
transform 1 0 580796 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6313
timestamp 1676037725
transform 1 0 581900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6325
timestamp 1676037725
transform 1 0 583004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6337
timestamp 1676037725
transform 1 0 584108 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6349
timestamp 1676037725
transform 1 0 585212 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6355
timestamp 1676037725
transform 1 0 585764 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6357
timestamp 1676037725
transform 1 0 585948 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6369
timestamp 1676037725
transform 1 0 587052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6381
timestamp 1676037725
transform 1 0 588156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6393
timestamp 1676037725
transform 1 0 589260 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6405
timestamp 1676037725
transform 1 0 590364 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6411
timestamp 1676037725
transform 1 0 590916 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6413
timestamp 1676037725
transform 1 0 591100 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6425
timestamp 1676037725
transform 1 0 592204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6437
timestamp 1676037725
transform 1 0 593308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6449
timestamp 1676037725
transform 1 0 594412 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6461
timestamp 1676037725
transform 1 0 595516 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6467
timestamp 1676037725
transform 1 0 596068 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6469
timestamp 1676037725
transform 1 0 596252 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6481
timestamp 1676037725
transform 1 0 597356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6493
timestamp 1676037725
transform 1 0 598460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6505
timestamp 1676037725
transform 1 0 599564 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6517
timestamp 1676037725
transform 1 0 600668 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6523
timestamp 1676037725
transform 1 0 601220 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6525
timestamp 1676037725
transform 1 0 601404 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6537
timestamp 1676037725
transform 1 0 602508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6549
timestamp 1676037725
transform 1 0 603612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6561
timestamp 1676037725
transform 1 0 604716 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6573
timestamp 1676037725
transform 1 0 605820 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6579
timestamp 1676037725
transform 1 0 606372 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6581
timestamp 1676037725
transform 1 0 606556 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6593
timestamp 1676037725
transform 1 0 607660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6605
timestamp 1676037725
transform 1 0 608764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6617
timestamp 1676037725
transform 1 0 609868 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6629
timestamp 1676037725
transform 1 0 610972 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6635
timestamp 1676037725
transform 1 0 611524 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6637
timestamp 1676037725
transform 1 0 611708 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6649
timestamp 1676037725
transform 1 0 612812 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6661
timestamp 1676037725
transform 1 0 613916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6673
timestamp 1676037725
transform 1 0 615020 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6685
timestamp 1676037725
transform 1 0 616124 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6691
timestamp 1676037725
transform 1 0 616676 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6693
timestamp 1676037725
transform 1 0 616860 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6705
timestamp 1676037725
transform 1 0 617964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6717
timestamp 1676037725
transform 1 0 619068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6729
timestamp 1676037725
transform 1 0 620172 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6741
timestamp 1676037725
transform 1 0 621276 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6747
timestamp 1676037725
transform 1 0 621828 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6749
timestamp 1676037725
transform 1 0 622012 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6761
timestamp 1676037725
transform 1 0 623116 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6773
timestamp 1676037725
transform 1 0 624220 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6785
timestamp 1676037725
transform 1 0 625324 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6797
timestamp 1676037725
transform 1 0 626428 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6803
timestamp 1676037725
transform 1 0 626980 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6805
timestamp 1676037725
transform 1 0 627164 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6817
timestamp 1676037725
transform 1 0 628268 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6829
timestamp 1676037725
transform 1 0 629372 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6841
timestamp 1676037725
transform 1 0 630476 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6853
timestamp 1676037725
transform 1 0 631580 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6859
timestamp 1676037725
transform 1 0 632132 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6861
timestamp 1676037725
transform 1 0 632316 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6873
timestamp 1676037725
transform 1 0 633420 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6885
timestamp 1676037725
transform 1 0 634524 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6897
timestamp 1676037725
transform 1 0 635628 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6909
timestamp 1676037725
transform 1 0 636732 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6915
timestamp 1676037725
transform 1 0 637284 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6917
timestamp 1676037725
transform 1 0 637468 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6929
timestamp 1676037725
transform 1 0 638572 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6941
timestamp 1676037725
transform 1 0 639676 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6953
timestamp 1676037725
transform 1 0 640780 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6965
timestamp 1676037725
transform 1 0 641884 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6971
timestamp 1676037725
transform 1 0 642436 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6973
timestamp 1676037725
transform 1 0 642620 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6985
timestamp 1676037725
transform 1 0 643724 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6997
timestamp 1676037725
transform 1 0 644828 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7009
timestamp 1676037725
transform 1 0 645932 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_7021
timestamp 1676037725
transform 1 0 647036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7027
timestamp 1676037725
transform 1 0 647588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_7029
timestamp 1676037725
transform 1 0 647772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7037
timestamp 1676037725
transform 1 0 648508 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1676037725
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1676037725
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1676037725
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1676037725
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1676037725
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1676037725
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1676037725
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1676037725
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1676037725
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1676037725
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1676037725
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1676037725
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1676037725
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1676037725
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1676037725
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1676037725
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1676037725
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1676037725
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1676037725
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1676037725
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1676037725
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1676037725
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1676037725
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1676037725
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1676037725
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1676037725
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1676037725
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1676037725
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1676037725
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1676037725
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_729
timestamp 1676037725
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_741
timestamp 1676037725
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_753
timestamp 1676037725
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_765
timestamp 1676037725
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1676037725
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1676037725
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_785
timestamp 1676037725
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_797
timestamp 1676037725
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_809
timestamp 1676037725
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_821
timestamp 1676037725
transform 1 0 76636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_833
timestamp 1676037725
transform 1 0 77740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_839
timestamp 1676037725
transform 1 0 78292 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_841
timestamp 1676037725
transform 1 0 78476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_853
timestamp 1676037725
transform 1 0 79580 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_865
timestamp 1676037725
transform 1 0 80684 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_873
timestamp 1676037725
transform 1 0 81420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_885
timestamp 1676037725
transform 1 0 82524 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_893
timestamp 1676037725
transform 1 0 83260 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_897
timestamp 1676037725
transform 1 0 83628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_909
timestamp 1676037725
transform 1 0 84732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_921
timestamp 1676037725
transform 1 0 85836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_933
timestamp 1676037725
transform 1 0 86940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_945
timestamp 1676037725
transform 1 0 88044 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_951
timestamp 1676037725
transform 1 0 88596 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_953
timestamp 1676037725
transform 1 0 88780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_965
timestamp 1676037725
transform 1 0 89884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_977
timestamp 1676037725
transform 1 0 90988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_989
timestamp 1676037725
transform 1 0 92092 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1001
timestamp 1676037725
transform 1 0 93196 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1007
timestamp 1676037725
transform 1 0 93748 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1009
timestamp 1676037725
transform 1 0 93932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1021
timestamp 1676037725
transform 1 0 95036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1033
timestamp 1676037725
transform 1 0 96140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1045
timestamp 1676037725
transform 1 0 97244 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1057
timestamp 1676037725
transform 1 0 98348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1063
timestamp 1676037725
transform 1 0 98900 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1065
timestamp 1676037725
transform 1 0 99084 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1077
timestamp 1676037725
transform 1 0 100188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1089
timestamp 1676037725
transform 1 0 101292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1101
timestamp 1676037725
transform 1 0 102396 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1113
timestamp 1676037725
transform 1 0 103500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1119
timestamp 1676037725
transform 1 0 104052 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1121
timestamp 1676037725
transform 1 0 104236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1133
timestamp 1676037725
transform 1 0 105340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1145
timestamp 1676037725
transform 1 0 106444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1157
timestamp 1676037725
transform 1 0 107548 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1169
timestamp 1676037725
transform 1 0 108652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1175
timestamp 1676037725
transform 1 0 109204 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1177
timestamp 1676037725
transform 1 0 109388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1189
timestamp 1676037725
transform 1 0 110492 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1195
timestamp 1676037725
transform 1 0 111044 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1198
timestamp 1676037725
transform 1 0 111320 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1211
timestamp 1676037725
transform 1 0 112516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1223
timestamp 1676037725
transform 1 0 113620 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1231
timestamp 1676037725
transform 1 0 114356 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1233
timestamp 1676037725
transform 1 0 114540 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1245
timestamp 1676037725
transform 1 0 115644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1257
timestamp 1676037725
transform 1 0 116748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1269
timestamp 1676037725
transform 1 0 117852 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_1281
timestamp 1676037725
transform 1 0 118956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1286
timestamp 1676037725
transform 1 0 119416 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1289
timestamp 1676037725
transform 1 0 119692 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1295
timestamp 1676037725
transform 1 0 120244 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1298
timestamp 1676037725
transform 1 0 120520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1306
timestamp 1676037725
transform 1 0 121256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1309
timestamp 1676037725
transform 1 0 121532 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1315
timestamp 1676037725
transform 1 0 122084 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1328
timestamp 1676037725
transform 1 0 123280 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1334
timestamp 1676037725
transform 1 0 123832 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1340
timestamp 1676037725
transform 1 0 124384 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1345
timestamp 1676037725
transform 1 0 124844 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1357
timestamp 1676037725
transform 1 0 125948 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1363
timestamp 1676037725
transform 1 0 126500 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1376
timestamp 1676037725
transform 1 0 127696 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1388
timestamp 1676037725
transform 1 0 128800 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1401
timestamp 1676037725
transform 1 0 129996 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1413
timestamp 1676037725
transform 1 0 131100 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1425
timestamp 1676037725
transform 1 0 132204 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1437
timestamp 1676037725
transform 1 0 133308 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1449
timestamp 1676037725
transform 1 0 134412 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1455
timestamp 1676037725
transform 1 0 134964 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1457
timestamp 1676037725
transform 1 0 135148 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1469
timestamp 1676037725
transform 1 0 136252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1481
timestamp 1676037725
transform 1 0 137356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1493
timestamp 1676037725
transform 1 0 138460 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1505
timestamp 1676037725
transform 1 0 139564 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1511
timestamp 1676037725
transform 1 0 140116 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1513
timestamp 1676037725
transform 1 0 140300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1525
timestamp 1676037725
transform 1 0 141404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1537
timestamp 1676037725
transform 1 0 142508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1549
timestamp 1676037725
transform 1 0 143612 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1561
timestamp 1676037725
transform 1 0 144716 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1567
timestamp 1676037725
transform 1 0 145268 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1569
timestamp 1676037725
transform 1 0 145452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1581
timestamp 1676037725
transform 1 0 146556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1593
timestamp 1676037725
transform 1 0 147660 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1605
timestamp 1676037725
transform 1 0 148764 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1617
timestamp 1676037725
transform 1 0 149868 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1623
timestamp 1676037725
transform 1 0 150420 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1625
timestamp 1676037725
transform 1 0 150604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1637
timestamp 1676037725
transform 1 0 151708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1649
timestamp 1676037725
transform 1 0 152812 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1661
timestamp 1676037725
transform 1 0 153916 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1673
timestamp 1676037725
transform 1 0 155020 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1679
timestamp 1676037725
transform 1 0 155572 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1681
timestamp 1676037725
transform 1 0 155756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1693
timestamp 1676037725
transform 1 0 156860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1705
timestamp 1676037725
transform 1 0 157964 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1717
timestamp 1676037725
transform 1 0 159068 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1729
timestamp 1676037725
transform 1 0 160172 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1735
timestamp 1676037725
transform 1 0 160724 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1737
timestamp 1676037725
transform 1 0 160908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1749
timestamp 1676037725
transform 1 0 162012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1761
timestamp 1676037725
transform 1 0 163116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1773
timestamp 1676037725
transform 1 0 164220 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1785
timestamp 1676037725
transform 1 0 165324 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1791
timestamp 1676037725
transform 1 0 165876 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1793
timestamp 1676037725
transform 1 0 166060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1805
timestamp 1676037725
transform 1 0 167164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1817
timestamp 1676037725
transform 1 0 168268 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1829
timestamp 1676037725
transform 1 0 169372 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1841
timestamp 1676037725
transform 1 0 170476 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1847
timestamp 1676037725
transform 1 0 171028 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1849
timestamp 1676037725
transform 1 0 171212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1861
timestamp 1676037725
transform 1 0 172316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1873
timestamp 1676037725
transform 1 0 173420 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1885
timestamp 1676037725
transform 1 0 174524 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1897
timestamp 1676037725
transform 1 0 175628 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1903
timestamp 1676037725
transform 1 0 176180 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1905
timestamp 1676037725
transform 1 0 176364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1917
timestamp 1676037725
transform 1 0 177468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1929
timestamp 1676037725
transform 1 0 178572 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1941
timestamp 1676037725
transform 1 0 179676 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1953
timestamp 1676037725
transform 1 0 180780 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1959
timestamp 1676037725
transform 1 0 181332 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1961
timestamp 1676037725
transform 1 0 181516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1973
timestamp 1676037725
transform 1 0 182620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1985
timestamp 1676037725
transform 1 0 183724 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1997
timestamp 1676037725
transform 1 0 184828 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2009
timestamp 1676037725
transform 1 0 185932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2015
timestamp 1676037725
transform 1 0 186484 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2017
timestamp 1676037725
transform 1 0 186668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2029
timestamp 1676037725
transform 1 0 187772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2041
timestamp 1676037725
transform 1 0 188876 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2053
timestamp 1676037725
transform 1 0 189980 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2065
timestamp 1676037725
transform 1 0 191084 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2071
timestamp 1676037725
transform 1 0 191636 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2073
timestamp 1676037725
transform 1 0 191820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2085
timestamp 1676037725
transform 1 0 192924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2097
timestamp 1676037725
transform 1 0 194028 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2109
timestamp 1676037725
transform 1 0 195132 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2121
timestamp 1676037725
transform 1 0 196236 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2127
timestamp 1676037725
transform 1 0 196788 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2129
timestamp 1676037725
transform 1 0 196972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2141
timestamp 1676037725
transform 1 0 198076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2153
timestamp 1676037725
transform 1 0 199180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2165
timestamp 1676037725
transform 1 0 200284 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_2177
timestamp 1676037725
transform 1 0 201388 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_2182
timestamp 1676037725
transform 1 0 201848 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_2185
timestamp 1676037725
transform 1 0 202124 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2196
timestamp 1676037725
transform 1 0 203136 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2208
timestamp 1676037725
transform 1 0 204240 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2220
timestamp 1676037725
transform 1 0 205344 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_2232
timestamp 1676037725
transform 1 0 206448 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2241
timestamp 1676037725
transform 1 0 207276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2253
timestamp 1676037725
transform 1 0 208380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2265
timestamp 1676037725
transform 1 0 209484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2277
timestamp 1676037725
transform 1 0 210588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2289
timestamp 1676037725
transform 1 0 211692 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2295
timestamp 1676037725
transform 1 0 212244 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_2297
timestamp 1676037725
transform 1 0 212428 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_2310
timestamp 1676037725
transform 1 0 213624 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_2323
timestamp 1676037725
transform 1 0 214820 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_2336
timestamp 1676037725
transform 1 0 216016 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2342
timestamp 1676037725
transform 1 0 216568 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_2350
timestamp 1676037725
transform 1 0 217304 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_2353
timestamp 1676037725
transform 1 0 217580 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2364
timestamp 1676037725
transform 1 0 218592 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2376
timestamp 1676037725
transform 1 0 219696 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2388
timestamp 1676037725
transform 1 0 220800 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_2400
timestamp 1676037725
transform 1 0 221904 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2409
timestamp 1676037725
transform 1 0 222732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2421
timestamp 1676037725
transform 1 0 223836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2433
timestamp 1676037725
transform 1 0 224940 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2445
timestamp 1676037725
transform 1 0 226044 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2457
timestamp 1676037725
transform 1 0 227148 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2463
timestamp 1676037725
transform 1 0 227700 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2465
timestamp 1676037725
transform 1 0 227884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2477
timestamp 1676037725
transform 1 0 228988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2489
timestamp 1676037725
transform 1 0 230092 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2501
timestamp 1676037725
transform 1 0 231196 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2513
timestamp 1676037725
transform 1 0 232300 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2519
timestamp 1676037725
transform 1 0 232852 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2521
timestamp 1676037725
transform 1 0 233036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2533
timestamp 1676037725
transform 1 0 234140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2545
timestamp 1676037725
transform 1 0 235244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2557
timestamp 1676037725
transform 1 0 236348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2569
timestamp 1676037725
transform 1 0 237452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2575
timestamp 1676037725
transform 1 0 238004 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2577
timestamp 1676037725
transform 1 0 238188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2589
timestamp 1676037725
transform 1 0 239292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2601
timestamp 1676037725
transform 1 0 240396 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2613
timestamp 1676037725
transform 1 0 241500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2625
timestamp 1676037725
transform 1 0 242604 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2631
timestamp 1676037725
transform 1 0 243156 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2633
timestamp 1676037725
transform 1 0 243340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2645
timestamp 1676037725
transform 1 0 244444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2657
timestamp 1676037725
transform 1 0 245548 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2669
timestamp 1676037725
transform 1 0 246652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2681
timestamp 1676037725
transform 1 0 247756 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2687
timestamp 1676037725
transform 1 0 248308 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2689
timestamp 1676037725
transform 1 0 248492 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2701
timestamp 1676037725
transform 1 0 249596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2713
timestamp 1676037725
transform 1 0 250700 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2725
timestamp 1676037725
transform 1 0 251804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2737
timestamp 1676037725
transform 1 0 252908 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2743
timestamp 1676037725
transform 1 0 253460 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2745
timestamp 1676037725
transform 1 0 253644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2757
timestamp 1676037725
transform 1 0 254748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2769
timestamp 1676037725
transform 1 0 255852 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2781
timestamp 1676037725
transform 1 0 256956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2793
timestamp 1676037725
transform 1 0 258060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2799
timestamp 1676037725
transform 1 0 258612 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2801
timestamp 1676037725
transform 1 0 258796 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2813
timestamp 1676037725
transform 1 0 259900 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_2825
timestamp 1676037725
transform 1 0 261004 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2835
timestamp 1676037725
transform 1 0 261924 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_2847
timestamp 1676037725
transform 1 0 263028 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2855
timestamp 1676037725
transform 1 0 263764 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2857
timestamp 1676037725
transform 1 0 263948 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2869
timestamp 1676037725
transform 1 0 265052 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2881
timestamp 1676037725
transform 1 0 266156 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2893
timestamp 1676037725
transform 1 0 267260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2905
timestamp 1676037725
transform 1 0 268364 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2911
timestamp 1676037725
transform 1 0 268916 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2913
timestamp 1676037725
transform 1 0 269100 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2925
timestamp 1676037725
transform 1 0 270204 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2937
timestamp 1676037725
transform 1 0 271308 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2949
timestamp 1676037725
transform 1 0 272412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2961
timestamp 1676037725
transform 1 0 273516 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2967
timestamp 1676037725
transform 1 0 274068 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2969
timestamp 1676037725
transform 1 0 274252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2981
timestamp 1676037725
transform 1 0 275356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2993
timestamp 1676037725
transform 1 0 276460 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3005
timestamp 1676037725
transform 1 0 277564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3017
timestamp 1676037725
transform 1 0 278668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3023
timestamp 1676037725
transform 1 0 279220 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3025
timestamp 1676037725
transform 1 0 279404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3037
timestamp 1676037725
transform 1 0 280508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3049
timestamp 1676037725
transform 1 0 281612 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3061
timestamp 1676037725
transform 1 0 282716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3073
timestamp 1676037725
transform 1 0 283820 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3079
timestamp 1676037725
transform 1 0 284372 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3081
timestamp 1676037725
transform 1 0 284556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3093
timestamp 1676037725
transform 1 0 285660 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3105
timestamp 1676037725
transform 1 0 286764 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3117
timestamp 1676037725
transform 1 0 287868 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3129
timestamp 1676037725
transform 1 0 288972 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3135
timestamp 1676037725
transform 1 0 289524 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3137
timestamp 1676037725
transform 1 0 289708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3149
timestamp 1676037725
transform 1 0 290812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3161
timestamp 1676037725
transform 1 0 291916 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3165
timestamp 1676037725
transform 1 0 292284 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3178
timestamp 1676037725
transform 1 0 293480 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3190
timestamp 1676037725
transform 1 0 294584 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3193
timestamp 1676037725
transform 1 0 294860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3205
timestamp 1676037725
transform 1 0 295964 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3217
timestamp 1676037725
transform 1 0 297068 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3229
timestamp 1676037725
transform 1 0 298172 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3241
timestamp 1676037725
transform 1 0 299276 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3247
timestamp 1676037725
transform 1 0 299828 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3249
timestamp 1676037725
transform 1 0 300012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3261
timestamp 1676037725
transform 1 0 301116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3273
timestamp 1676037725
transform 1 0 302220 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3285
timestamp 1676037725
transform 1 0 303324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3297
timestamp 1676037725
transform 1 0 304428 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3303
timestamp 1676037725
transform 1 0 304980 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3305
timestamp 1676037725
transform 1 0 305164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3317
timestamp 1676037725
transform 1 0 306268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3329
timestamp 1676037725
transform 1 0 307372 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3332
timestamp 1676037725
transform 1 0 307648 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3345
timestamp 1676037725
transform 1 0 308844 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3357
timestamp 1676037725
transform 1 0 309948 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3361
timestamp 1676037725
transform 1 0 310316 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3377
timestamp 1676037725
transform 1 0 311788 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3393
timestamp 1676037725
transform 1 0 313260 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3399
timestamp 1676037725
transform 1 0 313812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3411
timestamp 1676037725
transform 1 0 314916 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3415
timestamp 1676037725
transform 1 0 315284 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3417
timestamp 1676037725
transform 1 0 315468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3429
timestamp 1676037725
transform 1 0 316572 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3441
timestamp 1676037725
transform 1 0 317676 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3453
timestamp 1676037725
transform 1 0 318780 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3465
timestamp 1676037725
transform 1 0 319884 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3471
timestamp 1676037725
transform 1 0 320436 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3473
timestamp 1676037725
transform 1 0 320620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3485
timestamp 1676037725
transform 1 0 321724 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3497
timestamp 1676037725
transform 1 0 322828 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3509
timestamp 1676037725
transform 1 0 323932 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3521
timestamp 1676037725
transform 1 0 325036 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3527
timestamp 1676037725
transform 1 0 325588 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3529
timestamp 1676037725
transform 1 0 325772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3541
timestamp 1676037725
transform 1 0 326876 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3553
timestamp 1676037725
transform 1 0 327980 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3565
timestamp 1676037725
transform 1 0 329084 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3577
timestamp 1676037725
transform 1 0 330188 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3583
timestamp 1676037725
transform 1 0 330740 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3585
timestamp 1676037725
transform 1 0 330924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3597
timestamp 1676037725
transform 1 0 332028 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3609
timestamp 1676037725
transform 1 0 333132 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3621
timestamp 1676037725
transform 1 0 334236 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3633
timestamp 1676037725
transform 1 0 335340 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3639
timestamp 1676037725
transform 1 0 335892 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3641
timestamp 1676037725
transform 1 0 336076 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3653
timestamp 1676037725
transform 1 0 337180 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3661
timestamp 1676037725
transform 1 0 337916 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3666
timestamp 1676037725
transform 1 0 338376 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3679
timestamp 1676037725
transform 1 0 339572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3691
timestamp 1676037725
transform 1 0 340676 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3695
timestamp 1676037725
transform 1 0 341044 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3697
timestamp 1676037725
transform 1 0 341228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3709
timestamp 1676037725
transform 1 0 342332 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3721
timestamp 1676037725
transform 1 0 343436 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3733
timestamp 1676037725
transform 1 0 344540 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3745
timestamp 1676037725
transform 1 0 345644 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3751
timestamp 1676037725
transform 1 0 346196 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3753
timestamp 1676037725
transform 1 0 346380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3765
timestamp 1676037725
transform 1 0 347484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3777
timestamp 1676037725
transform 1 0 348588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3789
timestamp 1676037725
transform 1 0 349692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3801
timestamp 1676037725
transform 1 0 350796 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3807
timestamp 1676037725
transform 1 0 351348 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3809
timestamp 1676037725
transform 1 0 351532 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3821
timestamp 1676037725
transform 1 0 352636 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3829
timestamp 1676037725
transform 1 0 353372 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3833
timestamp 1676037725
transform 1 0 353740 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3846
timestamp 1676037725
transform 1 0 354936 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3858
timestamp 1676037725
transform 1 0 356040 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3865
timestamp 1676037725
transform 1 0 356684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3877
timestamp 1676037725
transform 1 0 357788 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3889
timestamp 1676037725
transform 1 0 358892 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3901
timestamp 1676037725
transform 1 0 359996 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3913
timestamp 1676037725
transform 1 0 361100 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3919
timestamp 1676037725
transform 1 0 361652 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3921
timestamp 1676037725
transform 1 0 361836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3933
timestamp 1676037725
transform 1 0 362940 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3945
timestamp 1676037725
transform 1 0 364044 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3957
timestamp 1676037725
transform 1 0 365148 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3969
timestamp 1676037725
transform 1 0 366252 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3975
timestamp 1676037725
transform 1 0 366804 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3977
timestamp 1676037725
transform 1 0 366988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3989
timestamp 1676037725
transform 1 0 368092 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4001
timestamp 1676037725
transform 1 0 369196 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4013
timestamp 1676037725
transform 1 0 370300 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4025
timestamp 1676037725
transform 1 0 371404 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4031
timestamp 1676037725
transform 1 0 371956 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4033
timestamp 1676037725
transform 1 0 372140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4045
timestamp 1676037725
transform 1 0 373244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4057
timestamp 1676037725
transform 1 0 374348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4069
timestamp 1676037725
transform 1 0 375452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4081
timestamp 1676037725
transform 1 0 376556 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4087
timestamp 1676037725
transform 1 0 377108 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4089
timestamp 1676037725
transform 1 0 377292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4101
timestamp 1676037725
transform 1 0 378396 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4113
timestamp 1676037725
transform 1 0 379500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4125
timestamp 1676037725
transform 1 0 380604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4137
timestamp 1676037725
transform 1 0 381708 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4143
timestamp 1676037725
transform 1 0 382260 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4145
timestamp 1676037725
transform 1 0 382444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4157
timestamp 1676037725
transform 1 0 383548 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4169
timestamp 1676037725
transform 1 0 384652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4181
timestamp 1676037725
transform 1 0 385756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4193
timestamp 1676037725
transform 1 0 386860 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4199
timestamp 1676037725
transform 1 0 387412 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4201
timestamp 1676037725
transform 1 0 387596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4213
timestamp 1676037725
transform 1 0 388700 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4225
timestamp 1676037725
transform 1 0 389804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4237
timestamp 1676037725
transform 1 0 390908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4249
timestamp 1676037725
transform 1 0 392012 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4255
timestamp 1676037725
transform 1 0 392564 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4257
timestamp 1676037725
transform 1 0 392748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4269
timestamp 1676037725
transform 1 0 393852 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4281
timestamp 1676037725
transform 1 0 394956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4293
timestamp 1676037725
transform 1 0 396060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4305
timestamp 1676037725
transform 1 0 397164 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4311
timestamp 1676037725
transform 1 0 397716 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4313
timestamp 1676037725
transform 1 0 397900 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4325
timestamp 1676037725
transform 1 0 399004 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4337
timestamp 1676037725
transform 1 0 400108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4349
timestamp 1676037725
transform 1 0 401212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4361
timestamp 1676037725
transform 1 0 402316 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4367
timestamp 1676037725
transform 1 0 402868 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4369
timestamp 1676037725
transform 1 0 403052 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4381
timestamp 1676037725
transform 1 0 404156 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4393
timestamp 1676037725
transform 1 0 405260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4405
timestamp 1676037725
transform 1 0 406364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4417
timestamp 1676037725
transform 1 0 407468 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4423
timestamp 1676037725
transform 1 0 408020 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4425
timestamp 1676037725
transform 1 0 408204 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4437
timestamp 1676037725
transform 1 0 409308 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4449
timestamp 1676037725
transform 1 0 410412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4461
timestamp 1676037725
transform 1 0 411516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4473
timestamp 1676037725
transform 1 0 412620 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4479
timestamp 1676037725
transform 1 0 413172 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4481
timestamp 1676037725
transform 1 0 413356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4493
timestamp 1676037725
transform 1 0 414460 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4505
timestamp 1676037725
transform 1 0 415564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4517
timestamp 1676037725
transform 1 0 416668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4529
timestamp 1676037725
transform 1 0 417772 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4535
timestamp 1676037725
transform 1 0 418324 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4537
timestamp 1676037725
transform 1 0 418508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4549
timestamp 1676037725
transform 1 0 419612 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4561
timestamp 1676037725
transform 1 0 420716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4573
timestamp 1676037725
transform 1 0 421820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4585
timestamp 1676037725
transform 1 0 422924 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4591
timestamp 1676037725
transform 1 0 423476 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4593
timestamp 1676037725
transform 1 0 423660 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4605
timestamp 1676037725
transform 1 0 424764 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4617
timestamp 1676037725
transform 1 0 425868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4629
timestamp 1676037725
transform 1 0 426972 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4641
timestamp 1676037725
transform 1 0 428076 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4647
timestamp 1676037725
transform 1 0 428628 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4649
timestamp 1676037725
transform 1 0 428812 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4661
timestamp 1676037725
transform 1 0 429916 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4673
timestamp 1676037725
transform 1 0 431020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4685
timestamp 1676037725
transform 1 0 432124 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4697
timestamp 1676037725
transform 1 0 433228 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4703
timestamp 1676037725
transform 1 0 433780 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4705
timestamp 1676037725
transform 1 0 433964 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4717
timestamp 1676037725
transform 1 0 435068 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4729
timestamp 1676037725
transform 1 0 436172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4741
timestamp 1676037725
transform 1 0 437276 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4753
timestamp 1676037725
transform 1 0 438380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4759
timestamp 1676037725
transform 1 0 438932 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4761
timestamp 1676037725
transform 1 0 439116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4773
timestamp 1676037725
transform 1 0 440220 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4785
timestamp 1676037725
transform 1 0 441324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4797
timestamp 1676037725
transform 1 0 442428 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4809
timestamp 1676037725
transform 1 0 443532 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4815
timestamp 1676037725
transform 1 0 444084 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4817
timestamp 1676037725
transform 1 0 444268 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4829
timestamp 1676037725
transform 1 0 445372 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4841
timestamp 1676037725
transform 1 0 446476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4853
timestamp 1676037725
transform 1 0 447580 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4865
timestamp 1676037725
transform 1 0 448684 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4871
timestamp 1676037725
transform 1 0 449236 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4873
timestamp 1676037725
transform 1 0 449420 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4885
timestamp 1676037725
transform 1 0 450524 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4897
timestamp 1676037725
transform 1 0 451628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4909
timestamp 1676037725
transform 1 0 452732 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4921
timestamp 1676037725
transform 1 0 453836 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4927
timestamp 1676037725
transform 1 0 454388 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4929
timestamp 1676037725
transform 1 0 454572 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4941
timestamp 1676037725
transform 1 0 455676 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4953
timestamp 1676037725
transform 1 0 456780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4965
timestamp 1676037725
transform 1 0 457884 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4977
timestamp 1676037725
transform 1 0 458988 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4983
timestamp 1676037725
transform 1 0 459540 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4985
timestamp 1676037725
transform 1 0 459724 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4997
timestamp 1676037725
transform 1 0 460828 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5009
timestamp 1676037725
transform 1 0 461932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5021
timestamp 1676037725
transform 1 0 463036 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5033
timestamp 1676037725
transform 1 0 464140 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5039
timestamp 1676037725
transform 1 0 464692 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5041
timestamp 1676037725
transform 1 0 464876 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5053
timestamp 1676037725
transform 1 0 465980 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5065
timestamp 1676037725
transform 1 0 467084 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5077
timestamp 1676037725
transform 1 0 468188 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5089
timestamp 1676037725
transform 1 0 469292 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5095
timestamp 1676037725
transform 1 0 469844 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5097
timestamp 1676037725
transform 1 0 470028 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5109
timestamp 1676037725
transform 1 0 471132 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5121
timestamp 1676037725
transform 1 0 472236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5133
timestamp 1676037725
transform 1 0 473340 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5145
timestamp 1676037725
transform 1 0 474444 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5151
timestamp 1676037725
transform 1 0 474996 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5153
timestamp 1676037725
transform 1 0 475180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5165
timestamp 1676037725
transform 1 0 476284 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5177
timestamp 1676037725
transform 1 0 477388 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5189
timestamp 1676037725
transform 1 0 478492 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5201
timestamp 1676037725
transform 1 0 479596 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5207
timestamp 1676037725
transform 1 0 480148 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5209
timestamp 1676037725
transform 1 0 480332 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5221
timestamp 1676037725
transform 1 0 481436 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5233
timestamp 1676037725
transform 1 0 482540 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5245
timestamp 1676037725
transform 1 0 483644 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5257
timestamp 1676037725
transform 1 0 484748 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5263
timestamp 1676037725
transform 1 0 485300 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5265
timestamp 1676037725
transform 1 0 485484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5277
timestamp 1676037725
transform 1 0 486588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5289
timestamp 1676037725
transform 1 0 487692 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5301
timestamp 1676037725
transform 1 0 488796 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5313
timestamp 1676037725
transform 1 0 489900 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5319
timestamp 1676037725
transform 1 0 490452 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5321
timestamp 1676037725
transform 1 0 490636 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5333
timestamp 1676037725
transform 1 0 491740 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5345
timestamp 1676037725
transform 1 0 492844 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5357
timestamp 1676037725
transform 1 0 493948 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5369
timestamp 1676037725
transform 1 0 495052 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5375
timestamp 1676037725
transform 1 0 495604 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5377
timestamp 1676037725
transform 1 0 495788 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5389
timestamp 1676037725
transform 1 0 496892 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5401
timestamp 1676037725
transform 1 0 497996 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5413
timestamp 1676037725
transform 1 0 499100 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5425
timestamp 1676037725
transform 1 0 500204 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5431
timestamp 1676037725
transform 1 0 500756 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5433
timestamp 1676037725
transform 1 0 500940 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5445
timestamp 1676037725
transform 1 0 502044 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5457
timestamp 1676037725
transform 1 0 503148 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5469
timestamp 1676037725
transform 1 0 504252 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5481
timestamp 1676037725
transform 1 0 505356 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5487
timestamp 1676037725
transform 1 0 505908 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5489
timestamp 1676037725
transform 1 0 506092 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5501
timestamp 1676037725
transform 1 0 507196 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5513
timestamp 1676037725
transform 1 0 508300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5525
timestamp 1676037725
transform 1 0 509404 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5537
timestamp 1676037725
transform 1 0 510508 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5543
timestamp 1676037725
transform 1 0 511060 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5545
timestamp 1676037725
transform 1 0 511244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5557
timestamp 1676037725
transform 1 0 512348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5569
timestamp 1676037725
transform 1 0 513452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5581
timestamp 1676037725
transform 1 0 514556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5593
timestamp 1676037725
transform 1 0 515660 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5599
timestamp 1676037725
transform 1 0 516212 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5601
timestamp 1676037725
transform 1 0 516396 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5613
timestamp 1676037725
transform 1 0 517500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5625
timestamp 1676037725
transform 1 0 518604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5637
timestamp 1676037725
transform 1 0 519708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5649
timestamp 1676037725
transform 1 0 520812 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5655
timestamp 1676037725
transform 1 0 521364 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5657
timestamp 1676037725
transform 1 0 521548 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5669
timestamp 1676037725
transform 1 0 522652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5681
timestamp 1676037725
transform 1 0 523756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5693
timestamp 1676037725
transform 1 0 524860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5705
timestamp 1676037725
transform 1 0 525964 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5711
timestamp 1676037725
transform 1 0 526516 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5713
timestamp 1676037725
transform 1 0 526700 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5725
timestamp 1676037725
transform 1 0 527804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5737
timestamp 1676037725
transform 1 0 528908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5749
timestamp 1676037725
transform 1 0 530012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5761
timestamp 1676037725
transform 1 0 531116 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5767
timestamp 1676037725
transform 1 0 531668 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5769
timestamp 1676037725
transform 1 0 531852 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5781
timestamp 1676037725
transform 1 0 532956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5793
timestamp 1676037725
transform 1 0 534060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5805
timestamp 1676037725
transform 1 0 535164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5817
timestamp 1676037725
transform 1 0 536268 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5823
timestamp 1676037725
transform 1 0 536820 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5825
timestamp 1676037725
transform 1 0 537004 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5837
timestamp 1676037725
transform 1 0 538108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5849
timestamp 1676037725
transform 1 0 539212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5861
timestamp 1676037725
transform 1 0 540316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5873
timestamp 1676037725
transform 1 0 541420 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5879
timestamp 1676037725
transform 1 0 541972 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5881
timestamp 1676037725
transform 1 0 542156 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5893
timestamp 1676037725
transform 1 0 543260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5905
timestamp 1676037725
transform 1 0 544364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5917
timestamp 1676037725
transform 1 0 545468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5929
timestamp 1676037725
transform 1 0 546572 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5935
timestamp 1676037725
transform 1 0 547124 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5937
timestamp 1676037725
transform 1 0 547308 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5949
timestamp 1676037725
transform 1 0 548412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5961
timestamp 1676037725
transform 1 0 549516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5973
timestamp 1676037725
transform 1 0 550620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5985
timestamp 1676037725
transform 1 0 551724 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5991
timestamp 1676037725
transform 1 0 552276 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5993
timestamp 1676037725
transform 1 0 552460 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6005
timestamp 1676037725
transform 1 0 553564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6017
timestamp 1676037725
transform 1 0 554668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6029
timestamp 1676037725
transform 1 0 555772 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6041
timestamp 1676037725
transform 1 0 556876 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6047
timestamp 1676037725
transform 1 0 557428 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6049
timestamp 1676037725
transform 1 0 557612 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6061
timestamp 1676037725
transform 1 0 558716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6073
timestamp 1676037725
transform 1 0 559820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6085
timestamp 1676037725
transform 1 0 560924 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6097
timestamp 1676037725
transform 1 0 562028 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6103
timestamp 1676037725
transform 1 0 562580 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6105
timestamp 1676037725
transform 1 0 562764 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6117
timestamp 1676037725
transform 1 0 563868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6129
timestamp 1676037725
transform 1 0 564972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6141
timestamp 1676037725
transform 1 0 566076 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6153
timestamp 1676037725
transform 1 0 567180 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6159
timestamp 1676037725
transform 1 0 567732 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6161
timestamp 1676037725
transform 1 0 567916 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6173
timestamp 1676037725
transform 1 0 569020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6185
timestamp 1676037725
transform 1 0 570124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6197
timestamp 1676037725
transform 1 0 571228 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6209
timestamp 1676037725
transform 1 0 572332 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6215
timestamp 1676037725
transform 1 0 572884 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6217
timestamp 1676037725
transform 1 0 573068 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6229
timestamp 1676037725
transform 1 0 574172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6241
timestamp 1676037725
transform 1 0 575276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6253
timestamp 1676037725
transform 1 0 576380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6265
timestamp 1676037725
transform 1 0 577484 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6271
timestamp 1676037725
transform 1 0 578036 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6273
timestamp 1676037725
transform 1 0 578220 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6285
timestamp 1676037725
transform 1 0 579324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6297
timestamp 1676037725
transform 1 0 580428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6309
timestamp 1676037725
transform 1 0 581532 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6321
timestamp 1676037725
transform 1 0 582636 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6327
timestamp 1676037725
transform 1 0 583188 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6329
timestamp 1676037725
transform 1 0 583372 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6341
timestamp 1676037725
transform 1 0 584476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6353
timestamp 1676037725
transform 1 0 585580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6365
timestamp 1676037725
transform 1 0 586684 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6377
timestamp 1676037725
transform 1 0 587788 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6383
timestamp 1676037725
transform 1 0 588340 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6385
timestamp 1676037725
transform 1 0 588524 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6397
timestamp 1676037725
transform 1 0 589628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6409
timestamp 1676037725
transform 1 0 590732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6421
timestamp 1676037725
transform 1 0 591836 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6433
timestamp 1676037725
transform 1 0 592940 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6439
timestamp 1676037725
transform 1 0 593492 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6441
timestamp 1676037725
transform 1 0 593676 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6453
timestamp 1676037725
transform 1 0 594780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6465
timestamp 1676037725
transform 1 0 595884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6477
timestamp 1676037725
transform 1 0 596988 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6489
timestamp 1676037725
transform 1 0 598092 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6495
timestamp 1676037725
transform 1 0 598644 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6497
timestamp 1676037725
transform 1 0 598828 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6509
timestamp 1676037725
transform 1 0 599932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6521
timestamp 1676037725
transform 1 0 601036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6533
timestamp 1676037725
transform 1 0 602140 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6545
timestamp 1676037725
transform 1 0 603244 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6551
timestamp 1676037725
transform 1 0 603796 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6553
timestamp 1676037725
transform 1 0 603980 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6565
timestamp 1676037725
transform 1 0 605084 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6577
timestamp 1676037725
transform 1 0 606188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6589
timestamp 1676037725
transform 1 0 607292 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6601
timestamp 1676037725
transform 1 0 608396 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6607
timestamp 1676037725
transform 1 0 608948 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6609
timestamp 1676037725
transform 1 0 609132 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6621
timestamp 1676037725
transform 1 0 610236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6633
timestamp 1676037725
transform 1 0 611340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6645
timestamp 1676037725
transform 1 0 612444 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6657
timestamp 1676037725
transform 1 0 613548 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6663
timestamp 1676037725
transform 1 0 614100 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6665
timestamp 1676037725
transform 1 0 614284 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6677
timestamp 1676037725
transform 1 0 615388 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6689
timestamp 1676037725
transform 1 0 616492 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6701
timestamp 1676037725
transform 1 0 617596 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6713
timestamp 1676037725
transform 1 0 618700 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6719
timestamp 1676037725
transform 1 0 619252 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6721
timestamp 1676037725
transform 1 0 619436 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6733
timestamp 1676037725
transform 1 0 620540 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6745
timestamp 1676037725
transform 1 0 621644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6757
timestamp 1676037725
transform 1 0 622748 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6769
timestamp 1676037725
transform 1 0 623852 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6775
timestamp 1676037725
transform 1 0 624404 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6777
timestamp 1676037725
transform 1 0 624588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6789
timestamp 1676037725
transform 1 0 625692 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6801
timestamp 1676037725
transform 1 0 626796 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6813
timestamp 1676037725
transform 1 0 627900 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6825
timestamp 1676037725
transform 1 0 629004 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6831
timestamp 1676037725
transform 1 0 629556 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6833
timestamp 1676037725
transform 1 0 629740 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6845
timestamp 1676037725
transform 1 0 630844 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6857
timestamp 1676037725
transform 1 0 631948 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6869
timestamp 1676037725
transform 1 0 633052 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6881
timestamp 1676037725
transform 1 0 634156 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6887
timestamp 1676037725
transform 1 0 634708 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6889
timestamp 1676037725
transform 1 0 634892 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6901
timestamp 1676037725
transform 1 0 635996 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6913
timestamp 1676037725
transform 1 0 637100 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6925
timestamp 1676037725
transform 1 0 638204 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6937
timestamp 1676037725
transform 1 0 639308 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6943
timestamp 1676037725
transform 1 0 639860 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6945
timestamp 1676037725
transform 1 0 640044 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6957
timestamp 1676037725
transform 1 0 641148 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6969
timestamp 1676037725
transform 1 0 642252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6981
timestamp 1676037725
transform 1 0 643356 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6993
timestamp 1676037725
transform 1 0 644460 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6999
timestamp 1676037725
transform 1 0 645012 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7001
timestamp 1676037725
transform 1 0 645196 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7013
timestamp 1676037725
transform 1 0 646300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7025
timestamp 1676037725
transform 1 0 647404 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7037
timestamp 1676037725
transform 1 0 648508 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1676037725
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1676037725
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1676037725
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_371
timestamp 1676037725
transform 1 0 35236 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_383
timestamp 1676037725
transform 1 0 36340 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_395
timestamp 1676037725
transform 1 0 37444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_407
timestamp 1676037725
transform 1 0 38548 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1676037725
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1676037725
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1676037725
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1676037725
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1676037725
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1676037725
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1676037725
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1676037725
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1676037725
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1676037725
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1676037725
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1676037725
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1676037725
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1676037725
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1676037725
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1676037725
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1676037725
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1676037725
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1676037725
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_669
timestamp 1676037725
transform 1 0 62652 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_675
timestamp 1676037725
transform 1 0 63204 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_678
timestamp 1676037725
transform 1 0 63480 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_692
timestamp 1676037725
transform 1 0 64768 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1676037725
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1676037725
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_725
timestamp 1676037725
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_737
timestamp 1676037725
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1676037725
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1676037725
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_757
timestamp 1676037725
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_769
timestamp 1676037725
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_781
timestamp 1676037725
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_793
timestamp 1676037725
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1676037725
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1676037725
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_813
timestamp 1676037725
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_825
timestamp 1676037725
transform 1 0 77004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_837
timestamp 1676037725
transform 1 0 78108 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_849
timestamp 1676037725
transform 1 0 79212 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_857
timestamp 1676037725
transform 1 0 79948 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_865
timestamp 1676037725
transform 1 0 80684 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_869
timestamp 1676037725
transform 1 0 81052 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_882
timestamp 1676037725
transform 1 0 82248 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_894
timestamp 1676037725
transform 1 0 83352 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_906
timestamp 1676037725
transform 1 0 84456 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_918
timestamp 1676037725
transform 1 0 85560 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_925
timestamp 1676037725
transform 1 0 86204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_937
timestamp 1676037725
transform 1 0 87308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_949
timestamp 1676037725
transform 1 0 88412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_961
timestamp 1676037725
transform 1 0 89516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_973
timestamp 1676037725
transform 1 0 90620 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_979
timestamp 1676037725
transform 1 0 91172 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_981
timestamp 1676037725
transform 1 0 91356 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_993
timestamp 1676037725
transform 1 0 92460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1005
timestamp 1676037725
transform 1 0 93564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1017
timestamp 1676037725
transform 1 0 94668 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1029
timestamp 1676037725
transform 1 0 95772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1035
timestamp 1676037725
transform 1 0 96324 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1037
timestamp 1676037725
transform 1 0 96508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1049
timestamp 1676037725
transform 1 0 97612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1061
timestamp 1676037725
transform 1 0 98716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1073
timestamp 1676037725
transform 1 0 99820 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1085
timestamp 1676037725
transform 1 0 100924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1091
timestamp 1676037725
transform 1 0 101476 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1093
timestamp 1676037725
transform 1 0 101660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1105
timestamp 1676037725
transform 1 0 102764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1117
timestamp 1676037725
transform 1 0 103868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1129
timestamp 1676037725
transform 1 0 104972 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1141
timestamp 1676037725
transform 1 0 106076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1147
timestamp 1676037725
transform 1 0 106628 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1149
timestamp 1676037725
transform 1 0 106812 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1153
timestamp 1676037725
transform 1 0 107180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1165
timestamp 1676037725
transform 1 0 108284 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1169
timestamp 1676037725
transform 1 0 108652 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1182
timestamp 1676037725
transform 1 0 109848 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1194
timestamp 1676037725
transform 1 0 110952 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1202
timestamp 1676037725
transform 1 0 111688 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1205
timestamp 1676037725
transform 1 0 111964 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1217
timestamp 1676037725
transform 1 0 113068 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1229
timestamp 1676037725
transform 1 0 114172 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1241
timestamp 1676037725
transform 1 0 115276 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1258
timestamp 1676037725
transform 1 0 116840 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1261
timestamp 1676037725
transform 1 0 117116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1265
timestamp 1676037725
transform 1 0 117484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1269
timestamp 1676037725
transform 1 0 117852 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1272
timestamp 1676037725
transform 1 0 118128 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1280
timestamp 1676037725
transform 1 0 118864 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1283
timestamp 1676037725
transform 1 0 119140 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1296
timestamp 1676037725
transform 1 0 120336 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1309
timestamp 1676037725
transform 1 0 121532 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1315
timestamp 1676037725
transform 1 0 122084 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1317
timestamp 1676037725
transform 1 0 122268 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1325
timestamp 1676037725
transform 1 0 123004 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1338
timestamp 1676037725
transform 1 0 124200 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1351
timestamp 1676037725
transform 1 0 125396 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1357
timestamp 1676037725
transform 1 0 125948 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_1369
timestamp 1676037725
transform 1 0 127052 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1373
timestamp 1676037725
transform 1 0 127420 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1385
timestamp 1676037725
transform 1 0 128524 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1397
timestamp 1676037725
transform 1 0 129628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1409
timestamp 1676037725
transform 1 0 130732 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1421
timestamp 1676037725
transform 1 0 131836 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1427
timestamp 1676037725
transform 1 0 132388 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1429
timestamp 1676037725
transform 1 0 132572 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1441
timestamp 1676037725
transform 1 0 133676 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1453
timestamp 1676037725
transform 1 0 134780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1465
timestamp 1676037725
transform 1 0 135884 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1477
timestamp 1676037725
transform 1 0 136988 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1483
timestamp 1676037725
transform 1 0 137540 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1485
timestamp 1676037725
transform 1 0 137724 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1497
timestamp 1676037725
transform 1 0 138828 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1509
timestamp 1676037725
transform 1 0 139932 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1521
timestamp 1676037725
transform 1 0 141036 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1533
timestamp 1676037725
transform 1 0 142140 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1539
timestamp 1676037725
transform 1 0 142692 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1541
timestamp 1676037725
transform 1 0 142876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1553
timestamp 1676037725
transform 1 0 143980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1565
timestamp 1676037725
transform 1 0 145084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1577
timestamp 1676037725
transform 1 0 146188 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1589
timestamp 1676037725
transform 1 0 147292 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1595
timestamp 1676037725
transform 1 0 147844 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1597
timestamp 1676037725
transform 1 0 148028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1609
timestamp 1676037725
transform 1 0 149132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1621
timestamp 1676037725
transform 1 0 150236 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1627
timestamp 1676037725
transform 1 0 150788 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1630
timestamp 1676037725
transform 1 0 151064 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1642
timestamp 1676037725
transform 1 0 152168 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1650
timestamp 1676037725
transform 1 0 152904 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1653
timestamp 1676037725
transform 1 0 153180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1665
timestamp 1676037725
transform 1 0 154284 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1669
timestamp 1676037725
transform 1 0 154652 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1683
timestamp 1676037725
transform 1 0 155940 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1696
timestamp 1676037725
transform 1 0 157136 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1709
timestamp 1676037725
transform 1 0 158332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1721
timestamp 1676037725
transform 1 0 159436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1733
timestamp 1676037725
transform 1 0 160540 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1745
timestamp 1676037725
transform 1 0 161644 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1757
timestamp 1676037725
transform 1 0 162748 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1763
timestamp 1676037725
transform 1 0 163300 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1765
timestamp 1676037725
transform 1 0 163484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1777
timestamp 1676037725
transform 1 0 164588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1789
timestamp 1676037725
transform 1 0 165692 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1793
timestamp 1676037725
transform 1 0 166060 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1796
timestamp 1676037725
transform 1 0 166336 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1808
timestamp 1676037725
transform 1 0 167440 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1821
timestamp 1676037725
transform 1 0 168636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1833
timestamp 1676037725
transform 1 0 169740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1836
timestamp 1676037725
transform 1 0 170016 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_1844
timestamp 1676037725
transform 1 0 170752 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1849
timestamp 1676037725
transform 1 0 171212 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1862
timestamp 1676037725
transform 1 0 172408 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1874
timestamp 1676037725
transform 1 0 173512 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1877
timestamp 1676037725
transform 1 0 173788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1889
timestamp 1676037725
transform 1 0 174892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1901
timestamp 1676037725
transform 1 0 175996 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1913
timestamp 1676037725
transform 1 0 177100 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1925
timestamp 1676037725
transform 1 0 178204 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1931
timestamp 1676037725
transform 1 0 178756 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1933
timestamp 1676037725
transform 1 0 178940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1945
timestamp 1676037725
transform 1 0 180044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1957
timestamp 1676037725
transform 1 0 181148 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1969
timestamp 1676037725
transform 1 0 182252 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1981
timestamp 1676037725
transform 1 0 183356 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1987
timestamp 1676037725
transform 1 0 183908 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1989
timestamp 1676037725
transform 1 0 184092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2001
timestamp 1676037725
transform 1 0 185196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2013
timestamp 1676037725
transform 1 0 186300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2025
timestamp 1676037725
transform 1 0 187404 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2037
timestamp 1676037725
transform 1 0 188508 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2043
timestamp 1676037725
transform 1 0 189060 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2045
timestamp 1676037725
transform 1 0 189244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2057
timestamp 1676037725
transform 1 0 190348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2069
timestamp 1676037725
transform 1 0 191452 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2081
timestamp 1676037725
transform 1 0 192556 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2093
timestamp 1676037725
transform 1 0 193660 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2099
timestamp 1676037725
transform 1 0 194212 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2101
timestamp 1676037725
transform 1 0 194396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2113
timestamp 1676037725
transform 1 0 195500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2125
timestamp 1676037725
transform 1 0 196604 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2137
timestamp 1676037725
transform 1 0 197708 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2149
timestamp 1676037725
transform 1 0 198812 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2155
timestamp 1676037725
transform 1 0 199364 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2157
timestamp 1676037725
transform 1 0 199548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2169
timestamp 1676037725
transform 1 0 200652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2181
timestamp 1676037725
transform 1 0 201756 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2193
timestamp 1676037725
transform 1 0 202860 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2205
timestamp 1676037725
transform 1 0 203964 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2211
timestamp 1676037725
transform 1 0 204516 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2213
timestamp 1676037725
transform 1 0 204700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2225
timestamp 1676037725
transform 1 0 205804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2237
timestamp 1676037725
transform 1 0 206908 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2249
timestamp 1676037725
transform 1 0 208012 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2261
timestamp 1676037725
transform 1 0 209116 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2267
timestamp 1676037725
transform 1 0 209668 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2269
timestamp 1676037725
transform 1 0 209852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2281
timestamp 1676037725
transform 1 0 210956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2293
timestamp 1676037725
transform 1 0 212060 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2305
timestamp 1676037725
transform 1 0 213164 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2317
timestamp 1676037725
transform 1 0 214268 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2323
timestamp 1676037725
transform 1 0 214820 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_2325
timestamp 1676037725
transform 1 0 215004 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_2331
timestamp 1676037725
transform 1 0 215556 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2344
timestamp 1676037725
transform 1 0 216752 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_2366
timestamp 1676037725
transform 1 0 218776 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_2372
timestamp 1676037725
transform 1 0 219328 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2381
timestamp 1676037725
transform 1 0 220156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2393
timestamp 1676037725
transform 1 0 221260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2405
timestamp 1676037725
transform 1 0 222364 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2417
timestamp 1676037725
transform 1 0 223468 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2429
timestamp 1676037725
transform 1 0 224572 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2435
timestamp 1676037725
transform 1 0 225124 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2437
timestamp 1676037725
transform 1 0 225308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2449
timestamp 1676037725
transform 1 0 226412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2461
timestamp 1676037725
transform 1 0 227516 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2473
timestamp 1676037725
transform 1 0 228620 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2485
timestamp 1676037725
transform 1 0 229724 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2491
timestamp 1676037725
transform 1 0 230276 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2493
timestamp 1676037725
transform 1 0 230460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2505
timestamp 1676037725
transform 1 0 231564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2517
timestamp 1676037725
transform 1 0 232668 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2529
timestamp 1676037725
transform 1 0 233772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2541
timestamp 1676037725
transform 1 0 234876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2547
timestamp 1676037725
transform 1 0 235428 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2549
timestamp 1676037725
transform 1 0 235612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2561
timestamp 1676037725
transform 1 0 236716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2573
timestamp 1676037725
transform 1 0 237820 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2585
timestamp 1676037725
transform 1 0 238924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2597
timestamp 1676037725
transform 1 0 240028 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2603
timestamp 1676037725
transform 1 0 240580 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2605
timestamp 1676037725
transform 1 0 240764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2617
timestamp 1676037725
transform 1 0 241868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2629
timestamp 1676037725
transform 1 0 242972 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2641
timestamp 1676037725
transform 1 0 244076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2653
timestamp 1676037725
transform 1 0 245180 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2659
timestamp 1676037725
transform 1 0 245732 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_2661
timestamp 1676037725
transform 1 0 245916 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_2665
timestamp 1676037725
transform 1 0 246284 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2678
timestamp 1676037725
transform 1 0 247480 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2690
timestamp 1676037725
transform 1 0 248584 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2702
timestamp 1676037725
transform 1 0 249688 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_2714
timestamp 1676037725
transform 1 0 250792 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2717
timestamp 1676037725
transform 1 0 251068 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2729
timestamp 1676037725
transform 1 0 252172 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2741
timestamp 1676037725
transform 1 0 253276 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2753
timestamp 1676037725
transform 1 0 254380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2765
timestamp 1676037725
transform 1 0 255484 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2771
timestamp 1676037725
transform 1 0 256036 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2773
timestamp 1676037725
transform 1 0 256220 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2785
timestamp 1676037725
transform 1 0 257324 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2797
timestamp 1676037725
transform 1 0 258428 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2809
timestamp 1676037725
transform 1 0 259532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2821
timestamp 1676037725
transform 1 0 260636 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2827
timestamp 1676037725
transform 1 0 261188 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2829
timestamp 1676037725
transform 1 0 261372 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2844
timestamp 1676037725
transform 1 0 262752 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2856
timestamp 1676037725
transform 1 0 263856 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2868
timestamp 1676037725
transform 1 0 264960 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_2880
timestamp 1676037725
transform 1 0 266064 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2885
timestamp 1676037725
transform 1 0 266524 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2897
timestamp 1676037725
transform 1 0 267628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2909
timestamp 1676037725
transform 1 0 268732 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2921
timestamp 1676037725
transform 1 0 269836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2933
timestamp 1676037725
transform 1 0 270940 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2939
timestamp 1676037725
transform 1 0 271492 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2941
timestamp 1676037725
transform 1 0 271676 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2953
timestamp 1676037725
transform 1 0 272780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2965
timestamp 1676037725
transform 1 0 273884 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2977
timestamp 1676037725
transform 1 0 274988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2989
timestamp 1676037725
transform 1 0 276092 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2995
timestamp 1676037725
transform 1 0 276644 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2997
timestamp 1676037725
transform 1 0 276828 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3009
timestamp 1676037725
transform 1 0 277932 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3021
timestamp 1676037725
transform 1 0 279036 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3033
timestamp 1676037725
transform 1 0 280140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3045
timestamp 1676037725
transform 1 0 281244 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3051
timestamp 1676037725
transform 1 0 281796 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3053
timestamp 1676037725
transform 1 0 281980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3065
timestamp 1676037725
transform 1 0 283084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3077
timestamp 1676037725
transform 1 0 284188 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3089
timestamp 1676037725
transform 1 0 285292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3101
timestamp 1676037725
transform 1 0 286396 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3107
timestamp 1676037725
transform 1 0 286948 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3109
timestamp 1676037725
transform 1 0 287132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3121
timestamp 1676037725
transform 1 0 288236 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3133
timestamp 1676037725
transform 1 0 289340 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3145
timestamp 1676037725
transform 1 0 290444 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3157
timestamp 1676037725
transform 1 0 291548 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3163
timestamp 1676037725
transform 1 0 292100 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3165
timestamp 1676037725
transform 1 0 292284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3177
timestamp 1676037725
transform 1 0 293388 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3189
timestamp 1676037725
transform 1 0 294492 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3201
timestamp 1676037725
transform 1 0 295596 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3213
timestamp 1676037725
transform 1 0 296700 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3219
timestamp 1676037725
transform 1 0 297252 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3221
timestamp 1676037725
transform 1 0 297436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3233
timestamp 1676037725
transform 1 0 298540 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3245
timestamp 1676037725
transform 1 0 299644 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3257
timestamp 1676037725
transform 1 0 300748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3269
timestamp 1676037725
transform 1 0 301852 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3275
timestamp 1676037725
transform 1 0 302404 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3277
timestamp 1676037725
transform 1 0 302588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3289
timestamp 1676037725
transform 1 0 303692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3301
timestamp 1676037725
transform 1 0 304796 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3313
timestamp 1676037725
transform 1 0 305900 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3325
timestamp 1676037725
transform 1 0 307004 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3331
timestamp 1676037725
transform 1 0 307556 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3333
timestamp 1676037725
transform 1 0 307740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3345
timestamp 1676037725
transform 1 0 308844 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3357
timestamp 1676037725
transform 1 0 309948 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3369
timestamp 1676037725
transform 1 0 311052 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3381
timestamp 1676037725
transform 1 0 312156 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3387
timestamp 1676037725
transform 1 0 312708 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3389
timestamp 1676037725
transform 1 0 312892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3401
timestamp 1676037725
transform 1 0 313996 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3413
timestamp 1676037725
transform 1 0 315100 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3425
timestamp 1676037725
transform 1 0 316204 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3437
timestamp 1676037725
transform 1 0 317308 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3443
timestamp 1676037725
transform 1 0 317860 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3445
timestamp 1676037725
transform 1 0 318044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3457
timestamp 1676037725
transform 1 0 319148 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3469
timestamp 1676037725
transform 1 0 320252 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3481
timestamp 1676037725
transform 1 0 321356 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3493
timestamp 1676037725
transform 1 0 322460 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3499
timestamp 1676037725
transform 1 0 323012 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3501
timestamp 1676037725
transform 1 0 323196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3513
timestamp 1676037725
transform 1 0 324300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3525
timestamp 1676037725
transform 1 0 325404 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3537
timestamp 1676037725
transform 1 0 326508 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3549
timestamp 1676037725
transform 1 0 327612 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3555
timestamp 1676037725
transform 1 0 328164 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3557
timestamp 1676037725
transform 1 0 328348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3569
timestamp 1676037725
transform 1 0 329452 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3581
timestamp 1676037725
transform 1 0 330556 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3593
timestamp 1676037725
transform 1 0 331660 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3605
timestamp 1676037725
transform 1 0 332764 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3611
timestamp 1676037725
transform 1 0 333316 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3613
timestamp 1676037725
transform 1 0 333500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3625
timestamp 1676037725
transform 1 0 334604 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3637
timestamp 1676037725
transform 1 0 335708 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3649
timestamp 1676037725
transform 1 0 336812 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3661
timestamp 1676037725
transform 1 0 337916 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3667
timestamp 1676037725
transform 1 0 338468 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3669
timestamp 1676037725
transform 1 0 338652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3681
timestamp 1676037725
transform 1 0 339756 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3693
timestamp 1676037725
transform 1 0 340860 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3705
timestamp 1676037725
transform 1 0 341964 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3717
timestamp 1676037725
transform 1 0 343068 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3723
timestamp 1676037725
transform 1 0 343620 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3725
timestamp 1676037725
transform 1 0 343804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3737
timestamp 1676037725
transform 1 0 344908 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3749
timestamp 1676037725
transform 1 0 346012 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3761
timestamp 1676037725
transform 1 0 347116 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3773
timestamp 1676037725
transform 1 0 348220 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3779
timestamp 1676037725
transform 1 0 348772 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3781
timestamp 1676037725
transform 1 0 348956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3793
timestamp 1676037725
transform 1 0 350060 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3805
timestamp 1676037725
transform 1 0 351164 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3817
timestamp 1676037725
transform 1 0 352268 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3829
timestamp 1676037725
transform 1 0 353372 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3835
timestamp 1676037725
transform 1 0 353924 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3837
timestamp 1676037725
transform 1 0 354108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3849
timestamp 1676037725
transform 1 0 355212 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3861
timestamp 1676037725
transform 1 0 356316 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3873
timestamp 1676037725
transform 1 0 357420 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3885
timestamp 1676037725
transform 1 0 358524 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3891
timestamp 1676037725
transform 1 0 359076 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3893
timestamp 1676037725
transform 1 0 359260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3905
timestamp 1676037725
transform 1 0 360364 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3917
timestamp 1676037725
transform 1 0 361468 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3929
timestamp 1676037725
transform 1 0 362572 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3941
timestamp 1676037725
transform 1 0 363676 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3947
timestamp 1676037725
transform 1 0 364228 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3949
timestamp 1676037725
transform 1 0 364412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3961
timestamp 1676037725
transform 1 0 365516 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3973
timestamp 1676037725
transform 1 0 366620 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3985
timestamp 1676037725
transform 1 0 367724 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3997
timestamp 1676037725
transform 1 0 368828 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4003
timestamp 1676037725
transform 1 0 369380 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4005
timestamp 1676037725
transform 1 0 369564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4017
timestamp 1676037725
transform 1 0 370668 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4029
timestamp 1676037725
transform 1 0 371772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4041
timestamp 1676037725
transform 1 0 372876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4053
timestamp 1676037725
transform 1 0 373980 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4059
timestamp 1676037725
transform 1 0 374532 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4061
timestamp 1676037725
transform 1 0 374716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4073
timestamp 1676037725
transform 1 0 375820 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4085
timestamp 1676037725
transform 1 0 376924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4097
timestamp 1676037725
transform 1 0 378028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4109
timestamp 1676037725
transform 1 0 379132 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4115
timestamp 1676037725
transform 1 0 379684 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4117
timestamp 1676037725
transform 1 0 379868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4129
timestamp 1676037725
transform 1 0 380972 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4141
timestamp 1676037725
transform 1 0 382076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4153
timestamp 1676037725
transform 1 0 383180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4165
timestamp 1676037725
transform 1 0 384284 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4171
timestamp 1676037725
transform 1 0 384836 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4173
timestamp 1676037725
transform 1 0 385020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4185
timestamp 1676037725
transform 1 0 386124 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4197
timestamp 1676037725
transform 1 0 387228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4209
timestamp 1676037725
transform 1 0 388332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4221
timestamp 1676037725
transform 1 0 389436 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4227
timestamp 1676037725
transform 1 0 389988 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4229
timestamp 1676037725
transform 1 0 390172 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4241
timestamp 1676037725
transform 1 0 391276 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4253
timestamp 1676037725
transform 1 0 392380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4265
timestamp 1676037725
transform 1 0 393484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4277
timestamp 1676037725
transform 1 0 394588 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4283
timestamp 1676037725
transform 1 0 395140 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4285
timestamp 1676037725
transform 1 0 395324 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4297
timestamp 1676037725
transform 1 0 396428 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4309
timestamp 1676037725
transform 1 0 397532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4321
timestamp 1676037725
transform 1 0 398636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4333
timestamp 1676037725
transform 1 0 399740 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4339
timestamp 1676037725
transform 1 0 400292 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4341
timestamp 1676037725
transform 1 0 400476 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4353
timestamp 1676037725
transform 1 0 401580 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4365
timestamp 1676037725
transform 1 0 402684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4377
timestamp 1676037725
transform 1 0 403788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4389
timestamp 1676037725
transform 1 0 404892 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4395
timestamp 1676037725
transform 1 0 405444 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4397
timestamp 1676037725
transform 1 0 405628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4409
timestamp 1676037725
transform 1 0 406732 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4421
timestamp 1676037725
transform 1 0 407836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4433
timestamp 1676037725
transform 1 0 408940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4445
timestamp 1676037725
transform 1 0 410044 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4451
timestamp 1676037725
transform 1 0 410596 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4453
timestamp 1676037725
transform 1 0 410780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4465
timestamp 1676037725
transform 1 0 411884 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4477
timestamp 1676037725
transform 1 0 412988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4489
timestamp 1676037725
transform 1 0 414092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4501
timestamp 1676037725
transform 1 0 415196 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4507
timestamp 1676037725
transform 1 0 415748 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4509
timestamp 1676037725
transform 1 0 415932 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4521
timestamp 1676037725
transform 1 0 417036 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4533
timestamp 1676037725
transform 1 0 418140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4545
timestamp 1676037725
transform 1 0 419244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4557
timestamp 1676037725
transform 1 0 420348 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4563
timestamp 1676037725
transform 1 0 420900 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4565
timestamp 1676037725
transform 1 0 421084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4577
timestamp 1676037725
transform 1 0 422188 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4589
timestamp 1676037725
transform 1 0 423292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4601
timestamp 1676037725
transform 1 0 424396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4613
timestamp 1676037725
transform 1 0 425500 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4619
timestamp 1676037725
transform 1 0 426052 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4621
timestamp 1676037725
transform 1 0 426236 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4633
timestamp 1676037725
transform 1 0 427340 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4645
timestamp 1676037725
transform 1 0 428444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4657
timestamp 1676037725
transform 1 0 429548 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4669
timestamp 1676037725
transform 1 0 430652 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4675
timestamp 1676037725
transform 1 0 431204 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4677
timestamp 1676037725
transform 1 0 431388 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4689
timestamp 1676037725
transform 1 0 432492 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4701
timestamp 1676037725
transform 1 0 433596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4713
timestamp 1676037725
transform 1 0 434700 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4725
timestamp 1676037725
transform 1 0 435804 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4731
timestamp 1676037725
transform 1 0 436356 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4733
timestamp 1676037725
transform 1 0 436540 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4745
timestamp 1676037725
transform 1 0 437644 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4757
timestamp 1676037725
transform 1 0 438748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4769
timestamp 1676037725
transform 1 0 439852 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4781
timestamp 1676037725
transform 1 0 440956 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4787
timestamp 1676037725
transform 1 0 441508 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4789
timestamp 1676037725
transform 1 0 441692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4801
timestamp 1676037725
transform 1 0 442796 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4813
timestamp 1676037725
transform 1 0 443900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4825
timestamp 1676037725
transform 1 0 445004 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4837
timestamp 1676037725
transform 1 0 446108 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4843
timestamp 1676037725
transform 1 0 446660 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4845
timestamp 1676037725
transform 1 0 446844 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4857
timestamp 1676037725
transform 1 0 447948 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4869
timestamp 1676037725
transform 1 0 449052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4881
timestamp 1676037725
transform 1 0 450156 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4893
timestamp 1676037725
transform 1 0 451260 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4899
timestamp 1676037725
transform 1 0 451812 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4901
timestamp 1676037725
transform 1 0 451996 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4913
timestamp 1676037725
transform 1 0 453100 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4925
timestamp 1676037725
transform 1 0 454204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4937
timestamp 1676037725
transform 1 0 455308 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4949
timestamp 1676037725
transform 1 0 456412 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4955
timestamp 1676037725
transform 1 0 456964 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4957
timestamp 1676037725
transform 1 0 457148 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4969
timestamp 1676037725
transform 1 0 458252 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4981
timestamp 1676037725
transform 1 0 459356 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4993
timestamp 1676037725
transform 1 0 460460 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5005
timestamp 1676037725
transform 1 0 461564 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5011
timestamp 1676037725
transform 1 0 462116 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5013
timestamp 1676037725
transform 1 0 462300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5025
timestamp 1676037725
transform 1 0 463404 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5037
timestamp 1676037725
transform 1 0 464508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5049
timestamp 1676037725
transform 1 0 465612 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5061
timestamp 1676037725
transform 1 0 466716 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5067
timestamp 1676037725
transform 1 0 467268 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5069
timestamp 1676037725
transform 1 0 467452 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5081
timestamp 1676037725
transform 1 0 468556 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5093
timestamp 1676037725
transform 1 0 469660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5105
timestamp 1676037725
transform 1 0 470764 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5117
timestamp 1676037725
transform 1 0 471868 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5123
timestamp 1676037725
transform 1 0 472420 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5125
timestamp 1676037725
transform 1 0 472604 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5137
timestamp 1676037725
transform 1 0 473708 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5149
timestamp 1676037725
transform 1 0 474812 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5161
timestamp 1676037725
transform 1 0 475916 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5173
timestamp 1676037725
transform 1 0 477020 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5179
timestamp 1676037725
transform 1 0 477572 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5181
timestamp 1676037725
transform 1 0 477756 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5193
timestamp 1676037725
transform 1 0 478860 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5205
timestamp 1676037725
transform 1 0 479964 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5217
timestamp 1676037725
transform 1 0 481068 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5229
timestamp 1676037725
transform 1 0 482172 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5235
timestamp 1676037725
transform 1 0 482724 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5237
timestamp 1676037725
transform 1 0 482908 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5249
timestamp 1676037725
transform 1 0 484012 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5261
timestamp 1676037725
transform 1 0 485116 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5273
timestamp 1676037725
transform 1 0 486220 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5285
timestamp 1676037725
transform 1 0 487324 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5291
timestamp 1676037725
transform 1 0 487876 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5293
timestamp 1676037725
transform 1 0 488060 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5305
timestamp 1676037725
transform 1 0 489164 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5317
timestamp 1676037725
transform 1 0 490268 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5329
timestamp 1676037725
transform 1 0 491372 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5341
timestamp 1676037725
transform 1 0 492476 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5347
timestamp 1676037725
transform 1 0 493028 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5349
timestamp 1676037725
transform 1 0 493212 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5361
timestamp 1676037725
transform 1 0 494316 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5373
timestamp 1676037725
transform 1 0 495420 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5385
timestamp 1676037725
transform 1 0 496524 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5397
timestamp 1676037725
transform 1 0 497628 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5403
timestamp 1676037725
transform 1 0 498180 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5405
timestamp 1676037725
transform 1 0 498364 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5417
timestamp 1676037725
transform 1 0 499468 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5429
timestamp 1676037725
transform 1 0 500572 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5441
timestamp 1676037725
transform 1 0 501676 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5453
timestamp 1676037725
transform 1 0 502780 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5459
timestamp 1676037725
transform 1 0 503332 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5461
timestamp 1676037725
transform 1 0 503516 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5473
timestamp 1676037725
transform 1 0 504620 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5485
timestamp 1676037725
transform 1 0 505724 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5497
timestamp 1676037725
transform 1 0 506828 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5509
timestamp 1676037725
transform 1 0 507932 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5515
timestamp 1676037725
transform 1 0 508484 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5517
timestamp 1676037725
transform 1 0 508668 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5529
timestamp 1676037725
transform 1 0 509772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5541
timestamp 1676037725
transform 1 0 510876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5553
timestamp 1676037725
transform 1 0 511980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5565
timestamp 1676037725
transform 1 0 513084 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5571
timestamp 1676037725
transform 1 0 513636 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5573
timestamp 1676037725
transform 1 0 513820 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5585
timestamp 1676037725
transform 1 0 514924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5597
timestamp 1676037725
transform 1 0 516028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5609
timestamp 1676037725
transform 1 0 517132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5621
timestamp 1676037725
transform 1 0 518236 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5627
timestamp 1676037725
transform 1 0 518788 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5629
timestamp 1676037725
transform 1 0 518972 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5641
timestamp 1676037725
transform 1 0 520076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5653
timestamp 1676037725
transform 1 0 521180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5665
timestamp 1676037725
transform 1 0 522284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5677
timestamp 1676037725
transform 1 0 523388 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5683
timestamp 1676037725
transform 1 0 523940 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5685
timestamp 1676037725
transform 1 0 524124 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5697
timestamp 1676037725
transform 1 0 525228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5709
timestamp 1676037725
transform 1 0 526332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5721
timestamp 1676037725
transform 1 0 527436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5733
timestamp 1676037725
transform 1 0 528540 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5739
timestamp 1676037725
transform 1 0 529092 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5741
timestamp 1676037725
transform 1 0 529276 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5753
timestamp 1676037725
transform 1 0 530380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5765
timestamp 1676037725
transform 1 0 531484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5777
timestamp 1676037725
transform 1 0 532588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5789
timestamp 1676037725
transform 1 0 533692 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5795
timestamp 1676037725
transform 1 0 534244 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5797
timestamp 1676037725
transform 1 0 534428 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5809
timestamp 1676037725
transform 1 0 535532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5821
timestamp 1676037725
transform 1 0 536636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5833
timestamp 1676037725
transform 1 0 537740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5845
timestamp 1676037725
transform 1 0 538844 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5851
timestamp 1676037725
transform 1 0 539396 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5853
timestamp 1676037725
transform 1 0 539580 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5865
timestamp 1676037725
transform 1 0 540684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5877
timestamp 1676037725
transform 1 0 541788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5889
timestamp 1676037725
transform 1 0 542892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5901
timestamp 1676037725
transform 1 0 543996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5907
timestamp 1676037725
transform 1 0 544548 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5909
timestamp 1676037725
transform 1 0 544732 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5921
timestamp 1676037725
transform 1 0 545836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5933
timestamp 1676037725
transform 1 0 546940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5945
timestamp 1676037725
transform 1 0 548044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5957
timestamp 1676037725
transform 1 0 549148 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5963
timestamp 1676037725
transform 1 0 549700 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5965
timestamp 1676037725
transform 1 0 549884 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5977
timestamp 1676037725
transform 1 0 550988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5989
timestamp 1676037725
transform 1 0 552092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6001
timestamp 1676037725
transform 1 0 553196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6013
timestamp 1676037725
transform 1 0 554300 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6019
timestamp 1676037725
transform 1 0 554852 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6021
timestamp 1676037725
transform 1 0 555036 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6033
timestamp 1676037725
transform 1 0 556140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6045
timestamp 1676037725
transform 1 0 557244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6057
timestamp 1676037725
transform 1 0 558348 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6069
timestamp 1676037725
transform 1 0 559452 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6075
timestamp 1676037725
transform 1 0 560004 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6077
timestamp 1676037725
transform 1 0 560188 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6089
timestamp 1676037725
transform 1 0 561292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6101
timestamp 1676037725
transform 1 0 562396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6113
timestamp 1676037725
transform 1 0 563500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6125
timestamp 1676037725
transform 1 0 564604 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6131
timestamp 1676037725
transform 1 0 565156 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6133
timestamp 1676037725
transform 1 0 565340 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6145
timestamp 1676037725
transform 1 0 566444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6157
timestamp 1676037725
transform 1 0 567548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6169
timestamp 1676037725
transform 1 0 568652 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6181
timestamp 1676037725
transform 1 0 569756 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6187
timestamp 1676037725
transform 1 0 570308 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6189
timestamp 1676037725
transform 1 0 570492 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6201
timestamp 1676037725
transform 1 0 571596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6213
timestamp 1676037725
transform 1 0 572700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6225
timestamp 1676037725
transform 1 0 573804 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6237
timestamp 1676037725
transform 1 0 574908 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6243
timestamp 1676037725
transform 1 0 575460 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6245
timestamp 1676037725
transform 1 0 575644 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6257
timestamp 1676037725
transform 1 0 576748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6269
timestamp 1676037725
transform 1 0 577852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6281
timestamp 1676037725
transform 1 0 578956 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6293
timestamp 1676037725
transform 1 0 580060 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6299
timestamp 1676037725
transform 1 0 580612 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6301
timestamp 1676037725
transform 1 0 580796 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6313
timestamp 1676037725
transform 1 0 581900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6325
timestamp 1676037725
transform 1 0 583004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6337
timestamp 1676037725
transform 1 0 584108 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6349
timestamp 1676037725
transform 1 0 585212 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6355
timestamp 1676037725
transform 1 0 585764 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6357
timestamp 1676037725
transform 1 0 585948 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6369
timestamp 1676037725
transform 1 0 587052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6381
timestamp 1676037725
transform 1 0 588156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6393
timestamp 1676037725
transform 1 0 589260 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6405
timestamp 1676037725
transform 1 0 590364 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6411
timestamp 1676037725
transform 1 0 590916 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6413
timestamp 1676037725
transform 1 0 591100 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6425
timestamp 1676037725
transform 1 0 592204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6437
timestamp 1676037725
transform 1 0 593308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6449
timestamp 1676037725
transform 1 0 594412 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6461
timestamp 1676037725
transform 1 0 595516 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6467
timestamp 1676037725
transform 1 0 596068 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6469
timestamp 1676037725
transform 1 0 596252 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6481
timestamp 1676037725
transform 1 0 597356 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6493
timestamp 1676037725
transform 1 0 598460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6505
timestamp 1676037725
transform 1 0 599564 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6517
timestamp 1676037725
transform 1 0 600668 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6523
timestamp 1676037725
transform 1 0 601220 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6525
timestamp 1676037725
transform 1 0 601404 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6537
timestamp 1676037725
transform 1 0 602508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6549
timestamp 1676037725
transform 1 0 603612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6561
timestamp 1676037725
transform 1 0 604716 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6573
timestamp 1676037725
transform 1 0 605820 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6579
timestamp 1676037725
transform 1 0 606372 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6581
timestamp 1676037725
transform 1 0 606556 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6593
timestamp 1676037725
transform 1 0 607660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6605
timestamp 1676037725
transform 1 0 608764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6617
timestamp 1676037725
transform 1 0 609868 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6629
timestamp 1676037725
transform 1 0 610972 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6635
timestamp 1676037725
transform 1 0 611524 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6637
timestamp 1676037725
transform 1 0 611708 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6649
timestamp 1676037725
transform 1 0 612812 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6661
timestamp 1676037725
transform 1 0 613916 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6673
timestamp 1676037725
transform 1 0 615020 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6685
timestamp 1676037725
transform 1 0 616124 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6691
timestamp 1676037725
transform 1 0 616676 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6693
timestamp 1676037725
transform 1 0 616860 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6705
timestamp 1676037725
transform 1 0 617964 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6717
timestamp 1676037725
transform 1 0 619068 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6729
timestamp 1676037725
transform 1 0 620172 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6741
timestamp 1676037725
transform 1 0 621276 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6747
timestamp 1676037725
transform 1 0 621828 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6749
timestamp 1676037725
transform 1 0 622012 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6761
timestamp 1676037725
transform 1 0 623116 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6773
timestamp 1676037725
transform 1 0 624220 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6785
timestamp 1676037725
transform 1 0 625324 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6797
timestamp 1676037725
transform 1 0 626428 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6803
timestamp 1676037725
transform 1 0 626980 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6805
timestamp 1676037725
transform 1 0 627164 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6817
timestamp 1676037725
transform 1 0 628268 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6829
timestamp 1676037725
transform 1 0 629372 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6841
timestamp 1676037725
transform 1 0 630476 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6853
timestamp 1676037725
transform 1 0 631580 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6859
timestamp 1676037725
transform 1 0 632132 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6861
timestamp 1676037725
transform 1 0 632316 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6873
timestamp 1676037725
transform 1 0 633420 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6885
timestamp 1676037725
transform 1 0 634524 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6897
timestamp 1676037725
transform 1 0 635628 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6909
timestamp 1676037725
transform 1 0 636732 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6915
timestamp 1676037725
transform 1 0 637284 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6917
timestamp 1676037725
transform 1 0 637468 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6929
timestamp 1676037725
transform 1 0 638572 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6941
timestamp 1676037725
transform 1 0 639676 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6953
timestamp 1676037725
transform 1 0 640780 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6965
timestamp 1676037725
transform 1 0 641884 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6971
timestamp 1676037725
transform 1 0 642436 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6973
timestamp 1676037725
transform 1 0 642620 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6985
timestamp 1676037725
transform 1 0 643724 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6997
timestamp 1676037725
transform 1 0 644828 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7009
timestamp 1676037725
transform 1 0 645932 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_7021
timestamp 1676037725
transform 1 0 647036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7027
timestamp 1676037725
transform 1 0 647588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_7029
timestamp 1676037725
transform 1 0 647772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7037
timestamp 1676037725
transform 1 0 648508 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_29
timestamp 1676037725
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_41
timestamp 1676037725
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1676037725
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_85
timestamp 1676037725
transform 1 0 8924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_97
timestamp 1676037725
transform 1 0 10028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1676037725
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_141
timestamp 1676037725
transform 1 0 14076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_153
timestamp 1676037725
transform 1 0 15180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1676037725
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_197
timestamp 1676037725
transform 1 0 19228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_209
timestamp 1676037725
transform 1 0 20332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp 1676037725
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_253
timestamp 1676037725
transform 1 0 24380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_265
timestamp 1676037725
transform 1 0 25484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1676037725
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_309
timestamp 1676037725
transform 1 0 29532 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_321
timestamp 1676037725
transform 1 0 30636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp 1676037725
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_345
timestamp 1676037725
transform 1 0 32844 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_355
timestamp 1676037725
transform 1 0 33764 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_363
timestamp 1676037725
transform 1 0 34500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_365
timestamp 1676037725
transform 1 0 34684 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_377
timestamp 1676037725
transform 1 0 35788 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_385
timestamp 1676037725
transform 1 0 36524 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_390
timestamp 1676037725
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_401
timestamp 1676037725
transform 1 0 37996 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_413
timestamp 1676037725
transform 1 0 39100 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_419
timestamp 1676037725
transform 1 0 39652 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_421
timestamp 1676037725
transform 1 0 39836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_433
timestamp 1676037725
transform 1 0 40940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_445
timestamp 1676037725
transform 1 0 42044 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_473
timestamp 1676037725
transform 1 0 44620 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_477
timestamp 1676037725
transform 1 0 44988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_489
timestamp 1676037725
transform 1 0 46092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_501
timestamp 1676037725
transform 1 0 47196 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1676037725
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_529
timestamp 1676037725
transform 1 0 49772 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_533
timestamp 1676037725
transform 1 0 50140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_545
timestamp 1676037725
transform 1 0 51244 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_557
timestamp 1676037725
transform 1 0 52348 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1676037725
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1676037725
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_585
timestamp 1676037725
transform 1 0 54924 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_589
timestamp 1676037725
transform 1 0 55292 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_601
timestamp 1676037725
transform 1 0 56396 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_604
timestamp 1676037725
transform 1 0 56672 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_614
timestamp 1676037725
transform 1 0 57592 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_617
timestamp 1676037725
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_625
timestamp 1676037725
transform 1 0 58604 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_629
timestamp 1676037725
transform 1 0 58972 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_639
timestamp 1676037725
transform 1 0 59892 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_643
timestamp 1676037725
transform 1 0 60260 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_645
timestamp 1676037725
transform 1 0 60444 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_649
timestamp 1676037725
transform 1 0 60812 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_652
timestamp 1676037725
transform 1 0 61088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_662
timestamp 1676037725
transform 1 0 62008 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_670
timestamp 1676037725
transform 1 0 62744 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_673
timestamp 1676037725
transform 1 0 63020 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_677
timestamp 1676037725
transform 1 0 63388 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_684
timestamp 1676037725
transform 1 0 64032 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_698
timestamp 1676037725
transform 1 0 65320 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_701
timestamp 1676037725
transform 1 0 65596 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_706
timestamp 1676037725
transform 1 0 66056 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_716
timestamp 1676037725
transform 1 0 66976 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_729
timestamp 1676037725
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_741
timestamp 1676037725
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_753
timestamp 1676037725
transform 1 0 70380 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_757
timestamp 1676037725
transform 1 0 70748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_769
timestamp 1676037725
transform 1 0 71852 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_772
timestamp 1676037725
transform 1 0 72128 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_782
timestamp 1676037725
transform 1 0 73048 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_785
timestamp 1676037725
transform 1 0 73324 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_795
timestamp 1676037725
transform 1 0 74244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_805
timestamp 1676037725
transform 1 0 75164 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_811
timestamp 1676037725
transform 1 0 75716 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_813
timestamp 1676037725
transform 1 0 75900 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_817
timestamp 1676037725
transform 1 0 76268 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_827
timestamp 1676037725
transform 1 0 77188 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_835
timestamp 1676037725
transform 1 0 77924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_838
timestamp 1676037725
transform 1 0 78200 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_841
timestamp 1676037725
transform 1 0 78476 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_852
timestamp 1676037725
transform 1 0 79488 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_856
timestamp 1676037725
transform 1 0 79856 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_866
timestamp 1676037725
transform 1 0 80776 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_869
timestamp 1676037725
transform 1 0 81052 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_881
timestamp 1676037725
transform 1 0 82156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_893
timestamp 1676037725
transform 1 0 83260 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_897
timestamp 1676037725
transform 1 0 83628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_909
timestamp 1676037725
transform 1 0 84732 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_921
timestamp 1676037725
transform 1 0 85836 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_925
timestamp 1676037725
transform 1 0 86204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_937
timestamp 1676037725
transform 1 0 87308 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_949
timestamp 1676037725
transform 1 0 88412 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_953
timestamp 1676037725
transform 1 0 88780 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_965
timestamp 1676037725
transform 1 0 89884 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_977
timestamp 1676037725
transform 1 0 90988 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_981
timestamp 1676037725
transform 1 0 91356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_993
timestamp 1676037725
transform 1 0 92460 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1005
timestamp 1676037725
transform 1 0 93564 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1009
timestamp 1676037725
transform 1 0 93932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1021
timestamp 1676037725
transform 1 0 95036 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1033
timestamp 1676037725
transform 1 0 96140 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1037
timestamp 1676037725
transform 1 0 96508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1049
timestamp 1676037725
transform 1 0 97612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1061
timestamp 1676037725
transform 1 0 98716 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1065
timestamp 1676037725
transform 1 0 99084 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1077
timestamp 1676037725
transform 1 0 100188 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1089
timestamp 1676037725
transform 1 0 101292 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1093
timestamp 1676037725
transform 1 0 101660 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1105
timestamp 1676037725
transform 1 0 102764 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1117
timestamp 1676037725
transform 1 0 103868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1121
timestamp 1676037725
transform 1 0 104236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1127
timestamp 1676037725
transform 1 0 104788 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1140
timestamp 1676037725
transform 1 0 105984 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1149
timestamp 1676037725
transform 1 0 106812 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1162
timestamp 1676037725
transform 1 0 108008 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1174
timestamp 1676037725
transform 1 0 109112 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1177
timestamp 1676037725
transform 1 0 109388 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1187
timestamp 1676037725
transform 1 0 110308 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1200
timestamp 1676037725
transform 1 0 111504 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1205
timestamp 1676037725
transform 1 0 111964 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1217
timestamp 1676037725
transform 1 0 113068 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1229
timestamp 1676037725
transform 1 0 114172 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1233
timestamp 1676037725
transform 1 0 114540 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1245
timestamp 1676037725
transform 1 0 115644 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1257
timestamp 1676037725
transform 1 0 116748 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1261
timestamp 1676037725
transform 1 0 117116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1270
timestamp 1676037725
transform 1 0 117944 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1276
timestamp 1676037725
transform 1 0 118496 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1286
timestamp 1676037725
transform 1 0 119416 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1289
timestamp 1676037725
transform 1 0 119692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1301
timestamp 1676037725
transform 1 0 120796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1314
timestamp 1676037725
transform 1 0 121992 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1317
timestamp 1676037725
transform 1 0 122268 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1329
timestamp 1676037725
transform 1 0 123372 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1342
timestamp 1676037725
transform 1 0 124568 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1345
timestamp 1676037725
transform 1 0 124844 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1349
timestamp 1676037725
transform 1 0 125212 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1352
timestamp 1676037725
transform 1 0 125488 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1365
timestamp 1676037725
transform 1 0 126684 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1371
timestamp 1676037725
transform 1 0 127236 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1373
timestamp 1676037725
transform 1 0 127420 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1385
timestamp 1676037725
transform 1 0 128524 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1397
timestamp 1676037725
transform 1 0 129628 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1401
timestamp 1676037725
transform 1 0 129996 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1413
timestamp 1676037725
transform 1 0 131100 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1425
timestamp 1676037725
transform 1 0 132204 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1429
timestamp 1676037725
transform 1 0 132572 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1441
timestamp 1676037725
transform 1 0 133676 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1453
timestamp 1676037725
transform 1 0 134780 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1457
timestamp 1676037725
transform 1 0 135148 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1469
timestamp 1676037725
transform 1 0 136252 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1481
timestamp 1676037725
transform 1 0 137356 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1485
timestamp 1676037725
transform 1 0 137724 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1497
timestamp 1676037725
transform 1 0 138828 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1509
timestamp 1676037725
transform 1 0 139932 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1513
timestamp 1676037725
transform 1 0 140300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1525
timestamp 1676037725
transform 1 0 141404 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1537
timestamp 1676037725
transform 1 0 142508 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1541
timestamp 1676037725
transform 1 0 142876 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1553
timestamp 1676037725
transform 1 0 143980 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1565
timestamp 1676037725
transform 1 0 145084 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1569
timestamp 1676037725
transform 1 0 145452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1581
timestamp 1676037725
transform 1 0 146556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1593
timestamp 1676037725
transform 1 0 147660 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1597
timestamp 1676037725
transform 1 0 148028 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1609
timestamp 1676037725
transform 1 0 149132 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1621
timestamp 1676037725
transform 1 0 150236 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1625
timestamp 1676037725
transform 1 0 150604 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1629
timestamp 1676037725
transform 1 0 150972 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1639
timestamp 1676037725
transform 1 0 151892 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1647
timestamp 1676037725
transform 1 0 152628 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1650
timestamp 1676037725
transform 1 0 152904 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1653
timestamp 1676037725
transform 1 0 153180 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1664
timestamp 1676037725
transform 1 0 154192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1668
timestamp 1676037725
transform 1 0 154560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1678
timestamp 1676037725
transform 1 0 155480 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1681
timestamp 1676037725
transform 1 0 155756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1693
timestamp 1676037725
transform 1 0 156860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1705
timestamp 1676037725
transform 1 0 157964 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1709
timestamp 1676037725
transform 1 0 158332 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1721
timestamp 1676037725
transform 1 0 159436 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1733
timestamp 1676037725
transform 1 0 160540 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1737
timestamp 1676037725
transform 1 0 160908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1749
timestamp 1676037725
transform 1 0 162012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1761
timestamp 1676037725
transform 1 0 163116 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1765
timestamp 1676037725
transform 1 0 163484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1777
timestamp 1676037725
transform 1 0 164588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1789
timestamp 1676037725
transform 1 0 165692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1793
timestamp 1676037725
transform 1 0 166060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1805
timestamp 1676037725
transform 1 0 167164 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1813
timestamp 1676037725
transform 1 0 167900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1818
timestamp 1676037725
transform 1 0 168360 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1821
timestamp 1676037725
transform 1 0 168636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1832
timestamp 1676037725
transform 1 0 169648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1845
timestamp 1676037725
transform 1 0 170844 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1849
timestamp 1676037725
transform 1 0 171212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1861
timestamp 1676037725
transform 1 0 172316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1873
timestamp 1676037725
transform 1 0 173420 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1877
timestamp 1676037725
transform 1 0 173788 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1889
timestamp 1676037725
transform 1 0 174892 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1901
timestamp 1676037725
transform 1 0 175996 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1905
timestamp 1676037725
transform 1 0 176364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1917
timestamp 1676037725
transform 1 0 177468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1929
timestamp 1676037725
transform 1 0 178572 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1933
timestamp 1676037725
transform 1 0 178940 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1945
timestamp 1676037725
transform 1 0 180044 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1957
timestamp 1676037725
transform 1 0 181148 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1961
timestamp 1676037725
transform 1 0 181516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1973
timestamp 1676037725
transform 1 0 182620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1985
timestamp 1676037725
transform 1 0 183724 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1989
timestamp 1676037725
transform 1 0 184092 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2001
timestamp 1676037725
transform 1 0 185196 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2013
timestamp 1676037725
transform 1 0 186300 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2017
timestamp 1676037725
transform 1 0 186668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2029
timestamp 1676037725
transform 1 0 187772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2041
timestamp 1676037725
transform 1 0 188876 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2045
timestamp 1676037725
transform 1 0 189244 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2057
timestamp 1676037725
transform 1 0 190348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2069
timestamp 1676037725
transform 1 0 191452 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2073
timestamp 1676037725
transform 1 0 191820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2085
timestamp 1676037725
transform 1 0 192924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2097
timestamp 1676037725
transform 1 0 194028 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2101
timestamp 1676037725
transform 1 0 194396 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2113
timestamp 1676037725
transform 1 0 195500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2125
timestamp 1676037725
transform 1 0 196604 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_2129
timestamp 1676037725
transform 1 0 196972 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_2137
timestamp 1676037725
transform 1 0 197708 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_2141
timestamp 1676037725
transform 1 0 198076 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_2154
timestamp 1676037725
transform 1 0 199272 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2157
timestamp 1676037725
transform 1 0 199548 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_2165
timestamp 1676037725
transform 1 0 200284 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2178
timestamp 1676037725
transform 1 0 201480 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2185
timestamp 1676037725
transform 1 0 202124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2197
timestamp 1676037725
transform 1 0 203228 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2209
timestamp 1676037725
transform 1 0 204332 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2213
timestamp 1676037725
transform 1 0 204700 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2225
timestamp 1676037725
transform 1 0 205804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2237
timestamp 1676037725
transform 1 0 206908 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2241
timestamp 1676037725
transform 1 0 207276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2253
timestamp 1676037725
transform 1 0 208380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2265
timestamp 1676037725
transform 1 0 209484 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2269
timestamp 1676037725
transform 1 0 209852 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2281
timestamp 1676037725
transform 1 0 210956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2293
timestamp 1676037725
transform 1 0 212060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_2297
timestamp 1676037725
transform 1 0 212428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_2305
timestamp 1676037725
transform 1 0 213164 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_2309
timestamp 1676037725
transform 1 0 213532 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_2322
timestamp 1676037725
transform 1 0 214728 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_2325
timestamp 1676037725
transform 1 0 215004 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2333
timestamp 1676037725
transform 1 0 215740 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_2350
timestamp 1676037725
transform 1 0 217304 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_2353
timestamp 1676037725
transform 1 0 217580 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_2357
timestamp 1676037725
transform 1 0 217948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2377
timestamp 1676037725
transform 1 0 219788 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_2381
timestamp 1676037725
transform 1 0 220156 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2385
timestamp 1676037725
transform 1 0 220524 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_2397
timestamp 1676037725
transform 1 0 221628 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2405
timestamp 1676037725
transform 1 0 222364 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2409
timestamp 1676037725
transform 1 0 222732 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2421
timestamp 1676037725
transform 1 0 223836 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2433
timestamp 1676037725
transform 1 0 224940 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2437
timestamp 1676037725
transform 1 0 225308 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2449
timestamp 1676037725
transform 1 0 226412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2461
timestamp 1676037725
transform 1 0 227516 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2465
timestamp 1676037725
transform 1 0 227884 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2477
timestamp 1676037725
transform 1 0 228988 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2489
timestamp 1676037725
transform 1 0 230092 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2493
timestamp 1676037725
transform 1 0 230460 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2505
timestamp 1676037725
transform 1 0 231564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2517
timestamp 1676037725
transform 1 0 232668 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2521
timestamp 1676037725
transform 1 0 233036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2533
timestamp 1676037725
transform 1 0 234140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2545
timestamp 1676037725
transform 1 0 235244 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2549
timestamp 1676037725
transform 1 0 235612 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2561
timestamp 1676037725
transform 1 0 236716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2573
timestamp 1676037725
transform 1 0 237820 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2577
timestamp 1676037725
transform 1 0 238188 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2589
timestamp 1676037725
transform 1 0 239292 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2601
timestamp 1676037725
transform 1 0 240396 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2605
timestamp 1676037725
transform 1 0 240764 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2617
timestamp 1676037725
transform 1 0 241868 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2629
timestamp 1676037725
transform 1 0 242972 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_2633
timestamp 1676037725
transform 1 0 243340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_2641
timestamp 1676037725
transform 1 0 244076 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_2645
timestamp 1676037725
transform 1 0 244444 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_2658
timestamp 1676037725
transform 1 0 245640 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2661
timestamp 1676037725
transform 1 0 245916 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2673
timestamp 1676037725
transform 1 0 247020 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2685
timestamp 1676037725
transform 1 0 248124 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2689
timestamp 1676037725
transform 1 0 248492 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2701
timestamp 1676037725
transform 1 0 249596 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2713
timestamp 1676037725
transform 1 0 250700 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2717
timestamp 1676037725
transform 1 0 251068 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2729
timestamp 1676037725
transform 1 0 252172 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2741
timestamp 1676037725
transform 1 0 253276 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2745
timestamp 1676037725
transform 1 0 253644 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2757
timestamp 1676037725
transform 1 0 254748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2769
timestamp 1676037725
transform 1 0 255852 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2773
timestamp 1676037725
transform 1 0 256220 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2785
timestamp 1676037725
transform 1 0 257324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2797
timestamp 1676037725
transform 1 0 258428 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_2801
timestamp 1676037725
transform 1 0 258796 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_2809
timestamp 1676037725
transform 1 0 259532 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_2813
timestamp 1676037725
transform 1 0 259900 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_2826
timestamp 1676037725
transform 1 0 261096 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2829
timestamp 1676037725
transform 1 0 261372 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2841
timestamp 1676037725
transform 1 0 262476 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2853
timestamp 1676037725
transform 1 0 263580 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2857
timestamp 1676037725
transform 1 0 263948 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2869
timestamp 1676037725
transform 1 0 265052 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2881
timestamp 1676037725
transform 1 0 266156 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2885
timestamp 1676037725
transform 1 0 266524 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2897
timestamp 1676037725
transform 1 0 267628 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2909
timestamp 1676037725
transform 1 0 268732 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2913
timestamp 1676037725
transform 1 0 269100 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2925
timestamp 1676037725
transform 1 0 270204 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2937
timestamp 1676037725
transform 1 0 271308 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2941
timestamp 1676037725
transform 1 0 271676 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2953
timestamp 1676037725
transform 1 0 272780 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2965
timestamp 1676037725
transform 1 0 273884 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2969
timestamp 1676037725
transform 1 0 274252 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2981
timestamp 1676037725
transform 1 0 275356 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2993
timestamp 1676037725
transform 1 0 276460 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2997
timestamp 1676037725
transform 1 0 276828 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3009
timestamp 1676037725
transform 1 0 277932 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3021
timestamp 1676037725
transform 1 0 279036 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3025
timestamp 1676037725
transform 1 0 279404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3037
timestamp 1676037725
transform 1 0 280508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3049
timestamp 1676037725
transform 1 0 281612 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3053
timestamp 1676037725
transform 1 0 281980 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3065
timestamp 1676037725
transform 1 0 283084 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3077
timestamp 1676037725
transform 1 0 284188 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3081
timestamp 1676037725
transform 1 0 284556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3093
timestamp 1676037725
transform 1 0 285660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3105
timestamp 1676037725
transform 1 0 286764 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3109
timestamp 1676037725
transform 1 0 287132 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3121
timestamp 1676037725
transform 1 0 288236 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3133
timestamp 1676037725
transform 1 0 289340 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3137
timestamp 1676037725
transform 1 0 289708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3149
timestamp 1676037725
transform 1 0 290812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3161
timestamp 1676037725
transform 1 0 291916 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3165
timestamp 1676037725
transform 1 0 292284 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3177
timestamp 1676037725
transform 1 0 293388 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3189
timestamp 1676037725
transform 1 0 294492 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3193
timestamp 1676037725
transform 1 0 294860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3205
timestamp 1676037725
transform 1 0 295964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3217
timestamp 1676037725
transform 1 0 297068 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3221
timestamp 1676037725
transform 1 0 297436 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3233
timestamp 1676037725
transform 1 0 298540 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3245
timestamp 1676037725
transform 1 0 299644 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3249
timestamp 1676037725
transform 1 0 300012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3261
timestamp 1676037725
transform 1 0 301116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3273
timestamp 1676037725
transform 1 0 302220 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3277
timestamp 1676037725
transform 1 0 302588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3289
timestamp 1676037725
transform 1 0 303692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3301
timestamp 1676037725
transform 1 0 304796 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3305
timestamp 1676037725
transform 1 0 305164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3317
timestamp 1676037725
transform 1 0 306268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3329
timestamp 1676037725
transform 1 0 307372 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3333
timestamp 1676037725
transform 1 0 307740 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3345
timestamp 1676037725
transform 1 0 308844 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3357
timestamp 1676037725
transform 1 0 309948 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3361
timestamp 1676037725
transform 1 0 310316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3373
timestamp 1676037725
transform 1 0 311420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3385
timestamp 1676037725
transform 1 0 312524 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3389
timestamp 1676037725
transform 1 0 312892 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3401
timestamp 1676037725
transform 1 0 313996 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3413
timestamp 1676037725
transform 1 0 315100 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3417
timestamp 1676037725
transform 1 0 315468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3429
timestamp 1676037725
transform 1 0 316572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3441
timestamp 1676037725
transform 1 0 317676 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3445
timestamp 1676037725
transform 1 0 318044 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3457
timestamp 1676037725
transform 1 0 319148 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3469
timestamp 1676037725
transform 1 0 320252 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3473
timestamp 1676037725
transform 1 0 320620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3485
timestamp 1676037725
transform 1 0 321724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3497
timestamp 1676037725
transform 1 0 322828 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3501
timestamp 1676037725
transform 1 0 323196 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3513
timestamp 1676037725
transform 1 0 324300 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3525
timestamp 1676037725
transform 1 0 325404 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3529
timestamp 1676037725
transform 1 0 325772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3541
timestamp 1676037725
transform 1 0 326876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3553
timestamp 1676037725
transform 1 0 327980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3557
timestamp 1676037725
transform 1 0 328348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3569
timestamp 1676037725
transform 1 0 329452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3581
timestamp 1676037725
transform 1 0 330556 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3585
timestamp 1676037725
transform 1 0 330924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3597
timestamp 1676037725
transform 1 0 332028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3609
timestamp 1676037725
transform 1 0 333132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3613
timestamp 1676037725
transform 1 0 333500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3625
timestamp 1676037725
transform 1 0 334604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3637
timestamp 1676037725
transform 1 0 335708 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3641
timestamp 1676037725
transform 1 0 336076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3653
timestamp 1676037725
transform 1 0 337180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3665
timestamp 1676037725
transform 1 0 338284 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3669
timestamp 1676037725
transform 1 0 338652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3681
timestamp 1676037725
transform 1 0 339756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3693
timestamp 1676037725
transform 1 0 340860 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3697
timestamp 1676037725
transform 1 0 341228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3709
timestamp 1676037725
transform 1 0 342332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3721
timestamp 1676037725
transform 1 0 343436 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3725
timestamp 1676037725
transform 1 0 343804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3737
timestamp 1676037725
transform 1 0 344908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3749
timestamp 1676037725
transform 1 0 346012 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3753
timestamp 1676037725
transform 1 0 346380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3765
timestamp 1676037725
transform 1 0 347484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3777
timestamp 1676037725
transform 1 0 348588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3781
timestamp 1676037725
transform 1 0 348956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3793
timestamp 1676037725
transform 1 0 350060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3805
timestamp 1676037725
transform 1 0 351164 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3809
timestamp 1676037725
transform 1 0 351532 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3821
timestamp 1676037725
transform 1 0 352636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3833
timestamp 1676037725
transform 1 0 353740 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3837
timestamp 1676037725
transform 1 0 354108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3849
timestamp 1676037725
transform 1 0 355212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3861
timestamp 1676037725
transform 1 0 356316 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3865
timestamp 1676037725
transform 1 0 356684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3877
timestamp 1676037725
transform 1 0 357788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3889
timestamp 1676037725
transform 1 0 358892 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3893
timestamp 1676037725
transform 1 0 359260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3905
timestamp 1676037725
transform 1 0 360364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3917
timestamp 1676037725
transform 1 0 361468 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3921
timestamp 1676037725
transform 1 0 361836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3933
timestamp 1676037725
transform 1 0 362940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3945
timestamp 1676037725
transform 1 0 364044 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3949
timestamp 1676037725
transform 1 0 364412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3961
timestamp 1676037725
transform 1 0 365516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3973
timestamp 1676037725
transform 1 0 366620 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3977
timestamp 1676037725
transform 1 0 366988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3989
timestamp 1676037725
transform 1 0 368092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4001
timestamp 1676037725
transform 1 0 369196 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4005
timestamp 1676037725
transform 1 0 369564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4017
timestamp 1676037725
transform 1 0 370668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4029
timestamp 1676037725
transform 1 0 371772 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4033
timestamp 1676037725
transform 1 0 372140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4045
timestamp 1676037725
transform 1 0 373244 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4057
timestamp 1676037725
transform 1 0 374348 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4061
timestamp 1676037725
transform 1 0 374716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4073
timestamp 1676037725
transform 1 0 375820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4085
timestamp 1676037725
transform 1 0 376924 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4089
timestamp 1676037725
transform 1 0 377292 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4101
timestamp 1676037725
transform 1 0 378396 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4113
timestamp 1676037725
transform 1 0 379500 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4117
timestamp 1676037725
transform 1 0 379868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4129
timestamp 1676037725
transform 1 0 380972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4141
timestamp 1676037725
transform 1 0 382076 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4145
timestamp 1676037725
transform 1 0 382444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4157
timestamp 1676037725
transform 1 0 383548 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4169
timestamp 1676037725
transform 1 0 384652 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4173
timestamp 1676037725
transform 1 0 385020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4185
timestamp 1676037725
transform 1 0 386124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4197
timestamp 1676037725
transform 1 0 387228 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4201
timestamp 1676037725
transform 1 0 387596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4213
timestamp 1676037725
transform 1 0 388700 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4225
timestamp 1676037725
transform 1 0 389804 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4229
timestamp 1676037725
transform 1 0 390172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4241
timestamp 1676037725
transform 1 0 391276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4253
timestamp 1676037725
transform 1 0 392380 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4257
timestamp 1676037725
transform 1 0 392748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4269
timestamp 1676037725
transform 1 0 393852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4281
timestamp 1676037725
transform 1 0 394956 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4285
timestamp 1676037725
transform 1 0 395324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4297
timestamp 1676037725
transform 1 0 396428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4309
timestamp 1676037725
transform 1 0 397532 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4313
timestamp 1676037725
transform 1 0 397900 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4325
timestamp 1676037725
transform 1 0 399004 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4337
timestamp 1676037725
transform 1 0 400108 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4341
timestamp 1676037725
transform 1 0 400476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4353
timestamp 1676037725
transform 1 0 401580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4365
timestamp 1676037725
transform 1 0 402684 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4369
timestamp 1676037725
transform 1 0 403052 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4381
timestamp 1676037725
transform 1 0 404156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4393
timestamp 1676037725
transform 1 0 405260 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4397
timestamp 1676037725
transform 1 0 405628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4409
timestamp 1676037725
transform 1 0 406732 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4421
timestamp 1676037725
transform 1 0 407836 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4425
timestamp 1676037725
transform 1 0 408204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4437
timestamp 1676037725
transform 1 0 409308 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4449
timestamp 1676037725
transform 1 0 410412 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4453
timestamp 1676037725
transform 1 0 410780 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4465
timestamp 1676037725
transform 1 0 411884 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4477
timestamp 1676037725
transform 1 0 412988 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4481
timestamp 1676037725
transform 1 0 413356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4493
timestamp 1676037725
transform 1 0 414460 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4505
timestamp 1676037725
transform 1 0 415564 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4509
timestamp 1676037725
transform 1 0 415932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4521
timestamp 1676037725
transform 1 0 417036 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4533
timestamp 1676037725
transform 1 0 418140 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4537
timestamp 1676037725
transform 1 0 418508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4549
timestamp 1676037725
transform 1 0 419612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4561
timestamp 1676037725
transform 1 0 420716 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4565
timestamp 1676037725
transform 1 0 421084 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4577
timestamp 1676037725
transform 1 0 422188 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4589
timestamp 1676037725
transform 1 0 423292 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4593
timestamp 1676037725
transform 1 0 423660 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4605
timestamp 1676037725
transform 1 0 424764 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4617
timestamp 1676037725
transform 1 0 425868 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4621
timestamp 1676037725
transform 1 0 426236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4633
timestamp 1676037725
transform 1 0 427340 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4645
timestamp 1676037725
transform 1 0 428444 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4649
timestamp 1676037725
transform 1 0 428812 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4661
timestamp 1676037725
transform 1 0 429916 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4673
timestamp 1676037725
transform 1 0 431020 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4677
timestamp 1676037725
transform 1 0 431388 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4689
timestamp 1676037725
transform 1 0 432492 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4701
timestamp 1676037725
transform 1 0 433596 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4705
timestamp 1676037725
transform 1 0 433964 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4717
timestamp 1676037725
transform 1 0 435068 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4729
timestamp 1676037725
transform 1 0 436172 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4733
timestamp 1676037725
transform 1 0 436540 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4745
timestamp 1676037725
transform 1 0 437644 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4757
timestamp 1676037725
transform 1 0 438748 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4761
timestamp 1676037725
transform 1 0 439116 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4773
timestamp 1676037725
transform 1 0 440220 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4785
timestamp 1676037725
transform 1 0 441324 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4789
timestamp 1676037725
transform 1 0 441692 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4801
timestamp 1676037725
transform 1 0 442796 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4813
timestamp 1676037725
transform 1 0 443900 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4817
timestamp 1676037725
transform 1 0 444268 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4829
timestamp 1676037725
transform 1 0 445372 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4841
timestamp 1676037725
transform 1 0 446476 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4845
timestamp 1676037725
transform 1 0 446844 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4857
timestamp 1676037725
transform 1 0 447948 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4869
timestamp 1676037725
transform 1 0 449052 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4873
timestamp 1676037725
transform 1 0 449420 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4885
timestamp 1676037725
transform 1 0 450524 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4897
timestamp 1676037725
transform 1 0 451628 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4901
timestamp 1676037725
transform 1 0 451996 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4913
timestamp 1676037725
transform 1 0 453100 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4925
timestamp 1676037725
transform 1 0 454204 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4929
timestamp 1676037725
transform 1 0 454572 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4941
timestamp 1676037725
transform 1 0 455676 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4953
timestamp 1676037725
transform 1 0 456780 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4957
timestamp 1676037725
transform 1 0 457148 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4969
timestamp 1676037725
transform 1 0 458252 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4981
timestamp 1676037725
transform 1 0 459356 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4985
timestamp 1676037725
transform 1 0 459724 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4997
timestamp 1676037725
transform 1 0 460828 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5009
timestamp 1676037725
transform 1 0 461932 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5013
timestamp 1676037725
transform 1 0 462300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5025
timestamp 1676037725
transform 1 0 463404 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5037
timestamp 1676037725
transform 1 0 464508 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5041
timestamp 1676037725
transform 1 0 464876 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5053
timestamp 1676037725
transform 1 0 465980 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5065
timestamp 1676037725
transform 1 0 467084 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5069
timestamp 1676037725
transform 1 0 467452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5081
timestamp 1676037725
transform 1 0 468556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5093
timestamp 1676037725
transform 1 0 469660 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5097
timestamp 1676037725
transform 1 0 470028 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5109
timestamp 1676037725
transform 1 0 471132 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5121
timestamp 1676037725
transform 1 0 472236 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5125
timestamp 1676037725
transform 1 0 472604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5137
timestamp 1676037725
transform 1 0 473708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5149
timestamp 1676037725
transform 1 0 474812 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5153
timestamp 1676037725
transform 1 0 475180 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5165
timestamp 1676037725
transform 1 0 476284 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5177
timestamp 1676037725
transform 1 0 477388 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5181
timestamp 1676037725
transform 1 0 477756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5193
timestamp 1676037725
transform 1 0 478860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5205
timestamp 1676037725
transform 1 0 479964 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5209
timestamp 1676037725
transform 1 0 480332 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5221
timestamp 1676037725
transform 1 0 481436 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5233
timestamp 1676037725
transform 1 0 482540 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5237
timestamp 1676037725
transform 1 0 482908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5249
timestamp 1676037725
transform 1 0 484012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5261
timestamp 1676037725
transform 1 0 485116 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5265
timestamp 1676037725
transform 1 0 485484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5277
timestamp 1676037725
transform 1 0 486588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5289
timestamp 1676037725
transform 1 0 487692 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5293
timestamp 1676037725
transform 1 0 488060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5305
timestamp 1676037725
transform 1 0 489164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5317
timestamp 1676037725
transform 1 0 490268 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5321
timestamp 1676037725
transform 1 0 490636 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5333
timestamp 1676037725
transform 1 0 491740 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5345
timestamp 1676037725
transform 1 0 492844 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5349
timestamp 1676037725
transform 1 0 493212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5361
timestamp 1676037725
transform 1 0 494316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5373
timestamp 1676037725
transform 1 0 495420 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5377
timestamp 1676037725
transform 1 0 495788 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5389
timestamp 1676037725
transform 1 0 496892 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5401
timestamp 1676037725
transform 1 0 497996 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5405
timestamp 1676037725
transform 1 0 498364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5417
timestamp 1676037725
transform 1 0 499468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5429
timestamp 1676037725
transform 1 0 500572 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5433
timestamp 1676037725
transform 1 0 500940 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5445
timestamp 1676037725
transform 1 0 502044 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5457
timestamp 1676037725
transform 1 0 503148 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5461
timestamp 1676037725
transform 1 0 503516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5473
timestamp 1676037725
transform 1 0 504620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5485
timestamp 1676037725
transform 1 0 505724 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5489
timestamp 1676037725
transform 1 0 506092 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5501
timestamp 1676037725
transform 1 0 507196 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5513
timestamp 1676037725
transform 1 0 508300 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5517
timestamp 1676037725
transform 1 0 508668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5529
timestamp 1676037725
transform 1 0 509772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5541
timestamp 1676037725
transform 1 0 510876 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5545
timestamp 1676037725
transform 1 0 511244 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5557
timestamp 1676037725
transform 1 0 512348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5569
timestamp 1676037725
transform 1 0 513452 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5573
timestamp 1676037725
transform 1 0 513820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5585
timestamp 1676037725
transform 1 0 514924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5597
timestamp 1676037725
transform 1 0 516028 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5601
timestamp 1676037725
transform 1 0 516396 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5613
timestamp 1676037725
transform 1 0 517500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5625
timestamp 1676037725
transform 1 0 518604 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5629
timestamp 1676037725
transform 1 0 518972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5641
timestamp 1676037725
transform 1 0 520076 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5653
timestamp 1676037725
transform 1 0 521180 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5657
timestamp 1676037725
transform 1 0 521548 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5669
timestamp 1676037725
transform 1 0 522652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5681
timestamp 1676037725
transform 1 0 523756 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5685
timestamp 1676037725
transform 1 0 524124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5697
timestamp 1676037725
transform 1 0 525228 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5709
timestamp 1676037725
transform 1 0 526332 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5713
timestamp 1676037725
transform 1 0 526700 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5725
timestamp 1676037725
transform 1 0 527804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5737
timestamp 1676037725
transform 1 0 528908 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5741
timestamp 1676037725
transform 1 0 529276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5753
timestamp 1676037725
transform 1 0 530380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5765
timestamp 1676037725
transform 1 0 531484 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5769
timestamp 1676037725
transform 1 0 531852 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5781
timestamp 1676037725
transform 1 0 532956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5793
timestamp 1676037725
transform 1 0 534060 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5797
timestamp 1676037725
transform 1 0 534428 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5809
timestamp 1676037725
transform 1 0 535532 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5821
timestamp 1676037725
transform 1 0 536636 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5825
timestamp 1676037725
transform 1 0 537004 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5837
timestamp 1676037725
transform 1 0 538108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5849
timestamp 1676037725
transform 1 0 539212 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5853
timestamp 1676037725
transform 1 0 539580 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5865
timestamp 1676037725
transform 1 0 540684 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5877
timestamp 1676037725
transform 1 0 541788 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5881
timestamp 1676037725
transform 1 0 542156 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5893
timestamp 1676037725
transform 1 0 543260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5905
timestamp 1676037725
transform 1 0 544364 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5909
timestamp 1676037725
transform 1 0 544732 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5921
timestamp 1676037725
transform 1 0 545836 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5933
timestamp 1676037725
transform 1 0 546940 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5937
timestamp 1676037725
transform 1 0 547308 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5949
timestamp 1676037725
transform 1 0 548412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5961
timestamp 1676037725
transform 1 0 549516 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5965
timestamp 1676037725
transform 1 0 549884 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5977
timestamp 1676037725
transform 1 0 550988 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5989
timestamp 1676037725
transform 1 0 552092 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5993
timestamp 1676037725
transform 1 0 552460 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6005
timestamp 1676037725
transform 1 0 553564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6017
timestamp 1676037725
transform 1 0 554668 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6021
timestamp 1676037725
transform 1 0 555036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6033
timestamp 1676037725
transform 1 0 556140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6045
timestamp 1676037725
transform 1 0 557244 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6049
timestamp 1676037725
transform 1 0 557612 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6061
timestamp 1676037725
transform 1 0 558716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6073
timestamp 1676037725
transform 1 0 559820 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6077
timestamp 1676037725
transform 1 0 560188 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6089
timestamp 1676037725
transform 1 0 561292 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6101
timestamp 1676037725
transform 1 0 562396 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6105
timestamp 1676037725
transform 1 0 562764 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6117
timestamp 1676037725
transform 1 0 563868 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6129
timestamp 1676037725
transform 1 0 564972 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6133
timestamp 1676037725
transform 1 0 565340 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6145
timestamp 1676037725
transform 1 0 566444 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6157
timestamp 1676037725
transform 1 0 567548 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6161
timestamp 1676037725
transform 1 0 567916 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6173
timestamp 1676037725
transform 1 0 569020 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6185
timestamp 1676037725
transform 1 0 570124 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6189
timestamp 1676037725
transform 1 0 570492 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6201
timestamp 1676037725
transform 1 0 571596 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6213
timestamp 1676037725
transform 1 0 572700 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6217
timestamp 1676037725
transform 1 0 573068 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6229
timestamp 1676037725
transform 1 0 574172 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6241
timestamp 1676037725
transform 1 0 575276 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6245
timestamp 1676037725
transform 1 0 575644 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6257
timestamp 1676037725
transform 1 0 576748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6269
timestamp 1676037725
transform 1 0 577852 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6273
timestamp 1676037725
transform 1 0 578220 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6285
timestamp 1676037725
transform 1 0 579324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6297
timestamp 1676037725
transform 1 0 580428 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6301
timestamp 1676037725
transform 1 0 580796 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6313
timestamp 1676037725
transform 1 0 581900 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6325
timestamp 1676037725
transform 1 0 583004 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6329
timestamp 1676037725
transform 1 0 583372 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6341
timestamp 1676037725
transform 1 0 584476 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6353
timestamp 1676037725
transform 1 0 585580 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6357
timestamp 1676037725
transform 1 0 585948 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6369
timestamp 1676037725
transform 1 0 587052 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6381
timestamp 1676037725
transform 1 0 588156 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6385
timestamp 1676037725
transform 1 0 588524 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6397
timestamp 1676037725
transform 1 0 589628 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6409
timestamp 1676037725
transform 1 0 590732 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6413
timestamp 1676037725
transform 1 0 591100 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6425
timestamp 1676037725
transform 1 0 592204 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6437
timestamp 1676037725
transform 1 0 593308 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6441
timestamp 1676037725
transform 1 0 593676 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6453
timestamp 1676037725
transform 1 0 594780 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6465
timestamp 1676037725
transform 1 0 595884 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6469
timestamp 1676037725
transform 1 0 596252 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6481
timestamp 1676037725
transform 1 0 597356 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6493
timestamp 1676037725
transform 1 0 598460 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6497
timestamp 1676037725
transform 1 0 598828 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6509
timestamp 1676037725
transform 1 0 599932 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6521
timestamp 1676037725
transform 1 0 601036 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6525
timestamp 1676037725
transform 1 0 601404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6537
timestamp 1676037725
transform 1 0 602508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6549
timestamp 1676037725
transform 1 0 603612 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6553
timestamp 1676037725
transform 1 0 603980 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6565
timestamp 1676037725
transform 1 0 605084 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6577
timestamp 1676037725
transform 1 0 606188 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6581
timestamp 1676037725
transform 1 0 606556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6593
timestamp 1676037725
transform 1 0 607660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6605
timestamp 1676037725
transform 1 0 608764 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6609
timestamp 1676037725
transform 1 0 609132 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6621
timestamp 1676037725
transform 1 0 610236 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6633
timestamp 1676037725
transform 1 0 611340 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6637
timestamp 1676037725
transform 1 0 611708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6649
timestamp 1676037725
transform 1 0 612812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6661
timestamp 1676037725
transform 1 0 613916 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6665
timestamp 1676037725
transform 1 0 614284 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6677
timestamp 1676037725
transform 1 0 615388 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6689
timestamp 1676037725
transform 1 0 616492 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6693
timestamp 1676037725
transform 1 0 616860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6705
timestamp 1676037725
transform 1 0 617964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6717
timestamp 1676037725
transform 1 0 619068 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6721
timestamp 1676037725
transform 1 0 619436 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6733
timestamp 1676037725
transform 1 0 620540 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6745
timestamp 1676037725
transform 1 0 621644 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6749
timestamp 1676037725
transform 1 0 622012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6761
timestamp 1676037725
transform 1 0 623116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6773
timestamp 1676037725
transform 1 0 624220 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6777
timestamp 1676037725
transform 1 0 624588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6789
timestamp 1676037725
transform 1 0 625692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6801
timestamp 1676037725
transform 1 0 626796 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6805
timestamp 1676037725
transform 1 0 627164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6817
timestamp 1676037725
transform 1 0 628268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6829
timestamp 1676037725
transform 1 0 629372 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6833
timestamp 1676037725
transform 1 0 629740 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6845
timestamp 1676037725
transform 1 0 630844 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6857
timestamp 1676037725
transform 1 0 631948 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6861
timestamp 1676037725
transform 1 0 632316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6873
timestamp 1676037725
transform 1 0 633420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6885
timestamp 1676037725
transform 1 0 634524 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6889
timestamp 1676037725
transform 1 0 634892 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6901
timestamp 1676037725
transform 1 0 635996 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6913
timestamp 1676037725
transform 1 0 637100 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6917
timestamp 1676037725
transform 1 0 637468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6929
timestamp 1676037725
transform 1 0 638572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6941
timestamp 1676037725
transform 1 0 639676 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6945
timestamp 1676037725
transform 1 0 640044 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6957
timestamp 1676037725
transform 1 0 641148 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6969
timestamp 1676037725
transform 1 0 642252 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6973
timestamp 1676037725
transform 1 0 642620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6985
timestamp 1676037725
transform 1 0 643724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6997
timestamp 1676037725
transform 1 0 644828 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7001
timestamp 1676037725
transform 1 0 645196 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7013
timestamp 1676037725
transform 1 0 646300 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_7025
timestamp 1676037725
transform 1 0 647404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_7029
timestamp 1676037725
transform 1 0 647772 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7037
timestamp 1676037725
transform 1 0 648508 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 648876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 648876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 648876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 648876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 648876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 648876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 648876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 648876 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 648876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 648876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1676037725
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1676037725
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1676037725
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1676037725
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1676037725
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1676037725
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1676037725
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1676037725
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1676037725
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1676037725
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1676037725
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1676037725
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1676037725
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1676037725
transform 1 0 83536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1676037725
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1676037725
transform 1 0 88688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1676037725
transform 1 0 91264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1676037725
transform 1 0 93840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1676037725
transform 1 0 96416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1676037725
transform 1 0 98992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1676037725
transform 1 0 101568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1676037725
transform 1 0 104144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1676037725
transform 1 0 106720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1676037725
transform 1 0 109296 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1676037725
transform 1 0 111872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1676037725
transform 1 0 114448 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1676037725
transform 1 0 117024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1676037725
transform 1 0 119600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1676037725
transform 1 0 122176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1676037725
transform 1 0 124752 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1676037725
transform 1 0 127328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1676037725
transform 1 0 129904 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1676037725
transform 1 0 132480 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1676037725
transform 1 0 135056 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1676037725
transform 1 0 137632 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 140208 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 142784 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 145360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 147936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 150512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 153088 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 155664 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 158240 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 160816 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 163392 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 165968 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 168544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 171120 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 173696 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 176272 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 178848 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 181424 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 184000 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 186576 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 189152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 191728 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 194304 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 196880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 199456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 202032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 204608 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 207184 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 209760 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 212336 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 214912 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 217488 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 220064 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 222640 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 225216 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 227792 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 230368 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 232944 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 235520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 238096 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 240672 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 243248 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 245824 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 248400 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 250976 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 253552 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 256128 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 258704 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 261280 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 263856 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 266432 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 269008 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 271584 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 274160 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 276736 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 279312 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 281888 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 284464 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 287040 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 289616 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 292192 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 294768 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 297344 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 299920 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 302496 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 305072 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 307648 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 310224 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 312800 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 315376 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 317952 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 320528 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 323104 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 325680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 328256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 330832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 333408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 335984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 338560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 341136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 343712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 346288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 348864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 351440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 354016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 356592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 359168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 361744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 364320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 366896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 369472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 372048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 374624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 377200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 379776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 382352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 384928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 387504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 390080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 392656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 395232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 397808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 400384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 402960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 405536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 408112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 410688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 413264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 415840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 418416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 420992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 423568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 426144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 428720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 431296 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 433872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 436448 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 439024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 441600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 444176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 446752 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 449328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 451904 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 454480 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 457056 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 459632 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 462208 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 464784 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 467360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 469936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 472512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 475088 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 477664 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 480240 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 482816 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 485392 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 487968 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 490544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 493120 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 495696 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 498272 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 500848 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 503424 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 506000 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 508576 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 511152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 513728 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 516304 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 518880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 521456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 524032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 526608 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 529184 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 531760 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 534336 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 536912 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 539488 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 542064 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 544640 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 547216 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 549792 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 552368 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 554944 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 557520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 560096 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 562672 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 565248 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 567824 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 570400 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 572976 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 575552 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 578128 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 580704 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 583280 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 585856 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 588432 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 591008 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 593584 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 596160 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 598736 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 601312 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 603888 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 606464 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 609040 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 611616 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 614192 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 616768 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 619344 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 621920 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 624496 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 627072 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 629648 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 632224 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 634800 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 637376 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 639952 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 642528 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 645104 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 647680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 88688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 93840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 98992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 104144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 109296 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 114448 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 119600 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 124752 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 129904 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 135056 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 140208 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 145360 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 150512 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 155664 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 160816 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 165968 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 171120 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 176272 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 181424 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 186576 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 191728 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 196880 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 202032 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 207184 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 212336 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 217488 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 222640 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 227792 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 232944 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 238096 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 243248 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 248400 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 253552 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 258704 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 263856 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 269008 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 274160 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 279312 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 284464 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 289616 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 294768 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 299920 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 305072 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 310224 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 315376 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 320528 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 325680 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 330832 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 335984 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 341136 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 346288 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 351440 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 356592 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 361744 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 366896 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 372048 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 377200 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 382352 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 387504 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 392656 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 397808 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 402960 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 408112 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 413264 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 418416 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 423568 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 428720 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 433872 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 439024 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 444176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 449328 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 454480 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 459632 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 464784 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 469936 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 475088 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 480240 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 485392 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 490544 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 495696 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 500848 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 506000 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 511152 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 516304 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 521456 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 526608 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 531760 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 536912 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 542064 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 547216 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 552368 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 557520 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 562672 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 567824 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 572976 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 578128 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 583280 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 588432 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 593584 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 598736 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 603888 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 609040 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 614192 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 619344 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 624496 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 629648 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 634800 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 639952 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 645104 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 91264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 96416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 101568 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 106720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 111872 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 117024 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 122176 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 127328 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 132480 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 137632 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 142784 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 147936 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 153088 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 158240 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 163392 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 168544 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 173696 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 178848 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 184000 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 189152 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 194304 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 199456 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 204608 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 209760 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 214912 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 220064 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 225216 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 230368 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 235520 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 240672 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 245824 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 250976 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 256128 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 261280 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 266432 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 271584 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 276736 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 281888 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 287040 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 292192 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 297344 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 302496 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 307648 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 312800 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 317952 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 323104 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 328256 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 333408 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 338560 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 343712 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 348864 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 354016 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 359168 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 364320 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 369472 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 374624 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 379776 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 384928 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 390080 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 395232 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 400384 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 405536 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 410688 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 415840 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 420992 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 426144 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 431296 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 436448 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 441600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 446752 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 451904 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 457056 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 462208 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 467360 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 472512 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 477664 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 482816 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 487968 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 493120 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 498272 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 503424 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 508576 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 513728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 518880 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 524032 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 529184 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 534336 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 539488 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 544640 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 549792 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 554944 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 560096 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 565248 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 570400 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 575552 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 580704 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 585856 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 591008 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 596160 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 601312 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 606464 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 611616 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 616768 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 621920 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 627072 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 632224 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 637376 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 642528 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 647680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 88688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 93840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 98992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 104144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 109296 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 114448 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 119600 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 124752 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 129904 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 135056 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 140208 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 145360 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 150512 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 155664 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 160816 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 165968 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 171120 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 176272 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 181424 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 186576 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 191728 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 196880 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 202032 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 207184 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 212336 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 217488 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 222640 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 227792 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 232944 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 238096 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 243248 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 248400 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 253552 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 258704 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 263856 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 269008 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 274160 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 279312 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 284464 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 289616 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 294768 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 299920 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 305072 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 310224 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 315376 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 320528 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 325680 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 330832 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 335984 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 341136 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 346288 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 351440 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 356592 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 361744 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 366896 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 372048 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 377200 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 382352 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 387504 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 392656 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 397808 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 402960 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 408112 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 413264 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 418416 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 423568 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 428720 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 433872 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 439024 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 444176 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 449328 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 454480 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 459632 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 464784 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 469936 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 475088 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 480240 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 485392 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 490544 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 495696 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 500848 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 506000 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 511152 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 516304 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 521456 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 526608 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 531760 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 536912 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 542064 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 547216 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 552368 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 557520 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 562672 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 567824 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 572976 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1676037725
transform 1 0 578128 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1676037725
transform 1 0 583280 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1676037725
transform 1 0 588432 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1676037725
transform 1 0 593584 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1676037725
transform 1 0 598736 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1676037725
transform 1 0 603888 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1676037725
transform 1 0 609040 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1676037725
transform 1 0 614192 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1676037725
transform 1 0 619344 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1676037725
transform 1 0 624496 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1676037725
transform 1 0 629648 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1676037725
transform 1 0 634800 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1676037725
transform 1 0 639952 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1676037725
transform 1 0 645104 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1676037725
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1676037725
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1676037725
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1676037725
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1676037725
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1676037725
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1676037725
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1676037725
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1676037725
transform 1 0 91264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1676037725
transform 1 0 96416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1676037725
transform 1 0 101568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1676037725
transform 1 0 106720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1676037725
transform 1 0 111872 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1676037725
transform 1 0 117024 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1676037725
transform 1 0 122176 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1676037725
transform 1 0 127328 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1676037725
transform 1 0 132480 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1676037725
transform 1 0 137632 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1676037725
transform 1 0 142784 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1676037725
transform 1 0 147936 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1676037725
transform 1 0 153088 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1676037725
transform 1 0 158240 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1676037725
transform 1 0 163392 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1676037725
transform 1 0 168544 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1676037725
transform 1 0 173696 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1676037725
transform 1 0 178848 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1676037725
transform 1 0 184000 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1676037725
transform 1 0 189152 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1676037725
transform 1 0 194304 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1676037725
transform 1 0 199456 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1676037725
transform 1 0 204608 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1676037725
transform 1 0 209760 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1676037725
transform 1 0 214912 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1676037725
transform 1 0 220064 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1676037725
transform 1 0 225216 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1676037725
transform 1 0 230368 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1676037725
transform 1 0 235520 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1676037725
transform 1 0 240672 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1676037725
transform 1 0 245824 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1676037725
transform 1 0 250976 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1676037725
transform 1 0 256128 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1676037725
transform 1 0 261280 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1676037725
transform 1 0 266432 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1676037725
transform 1 0 271584 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1676037725
transform 1 0 276736 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1676037725
transform 1 0 281888 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1676037725
transform 1 0 287040 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1676037725
transform 1 0 292192 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1676037725
transform 1 0 297344 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1676037725
transform 1 0 302496 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1676037725
transform 1 0 307648 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1676037725
transform 1 0 312800 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1676037725
transform 1 0 317952 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1676037725
transform 1 0 323104 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1676037725
transform 1 0 328256 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1676037725
transform 1 0 333408 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1676037725
transform 1 0 338560 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1676037725
transform 1 0 343712 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1676037725
transform 1 0 348864 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1676037725
transform 1 0 354016 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1676037725
transform 1 0 359168 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1676037725
transform 1 0 364320 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1676037725
transform 1 0 369472 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1676037725
transform 1 0 374624 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1676037725
transform 1 0 379776 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1676037725
transform 1 0 384928 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1676037725
transform 1 0 390080 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1676037725
transform 1 0 395232 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1676037725
transform 1 0 400384 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1676037725
transform 1 0 405536 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1676037725
transform 1 0 410688 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1676037725
transform 1 0 415840 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1676037725
transform 1 0 420992 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1676037725
transform 1 0 426144 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1676037725
transform 1 0 431296 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1676037725
transform 1 0 436448 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1676037725
transform 1 0 441600 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1676037725
transform 1 0 446752 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1676037725
transform 1 0 451904 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1676037725
transform 1 0 457056 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1676037725
transform 1 0 462208 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1676037725
transform 1 0 467360 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1676037725
transform 1 0 472512 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1676037725
transform 1 0 477664 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1676037725
transform 1 0 482816 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1676037725
transform 1 0 487968 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1676037725
transform 1 0 493120 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1676037725
transform 1 0 498272 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1676037725
transform 1 0 503424 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1676037725
transform 1 0 508576 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1676037725
transform 1 0 513728 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1676037725
transform 1 0 518880 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1676037725
transform 1 0 524032 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1676037725
transform 1 0 529184 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1676037725
transform 1 0 534336 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1676037725
transform 1 0 539488 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1676037725
transform 1 0 544640 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1676037725
transform 1 0 549792 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1676037725
transform 1 0 554944 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1676037725
transform 1 0 560096 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1676037725
transform 1 0 565248 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1676037725
transform 1 0 570400 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1676037725
transform 1 0 575552 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1676037725
transform 1 0 580704 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1676037725
transform 1 0 585856 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1676037725
transform 1 0 591008 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1676037725
transform 1 0 596160 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1676037725
transform 1 0 601312 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1676037725
transform 1 0 606464 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1676037725
transform 1 0 611616 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1676037725
transform 1 0 616768 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1676037725
transform 1 0 621920 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1676037725
transform 1 0 627072 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1676037725
transform 1 0 632224 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1676037725
transform 1 0 637376 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1676037725
transform 1 0 642528 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1676037725
transform 1 0 647680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1676037725
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1676037725
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1676037725
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1676037725
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1676037725
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1676037725
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1676037725
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1676037725
transform 1 0 88688 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1676037725
transform 1 0 93840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1676037725
transform 1 0 98992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1676037725
transform 1 0 104144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1676037725
transform 1 0 109296 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1676037725
transform 1 0 114448 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1676037725
transform 1 0 119600 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1676037725
transform 1 0 124752 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1676037725
transform 1 0 129904 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1676037725
transform 1 0 135056 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1676037725
transform 1 0 140208 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1676037725
transform 1 0 145360 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1676037725
transform 1 0 150512 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1676037725
transform 1 0 155664 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1676037725
transform 1 0 160816 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1676037725
transform 1 0 165968 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1676037725
transform 1 0 171120 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1676037725
transform 1 0 176272 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1676037725
transform 1 0 181424 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1676037725
transform 1 0 186576 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1676037725
transform 1 0 191728 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1676037725
transform 1 0 196880 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1676037725
transform 1 0 202032 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1676037725
transform 1 0 207184 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1676037725
transform 1 0 212336 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1676037725
transform 1 0 217488 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1676037725
transform 1 0 222640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1676037725
transform 1 0 227792 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1676037725
transform 1 0 232944 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1676037725
transform 1 0 238096 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1676037725
transform 1 0 243248 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1676037725
transform 1 0 248400 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1676037725
transform 1 0 253552 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1676037725
transform 1 0 258704 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1676037725
transform 1 0 263856 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1676037725
transform 1 0 269008 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1676037725
transform 1 0 274160 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1676037725
transform 1 0 279312 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1676037725
transform 1 0 284464 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1676037725
transform 1 0 289616 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1676037725
transform 1 0 294768 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1676037725
transform 1 0 299920 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1676037725
transform 1 0 305072 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1676037725
transform 1 0 310224 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1676037725
transform 1 0 315376 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1676037725
transform 1 0 320528 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1676037725
transform 1 0 325680 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1676037725
transform 1 0 330832 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1676037725
transform 1 0 335984 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1676037725
transform 1 0 341136 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1676037725
transform 1 0 346288 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1676037725
transform 1 0 351440 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1676037725
transform 1 0 356592 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1676037725
transform 1 0 361744 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1676037725
transform 1 0 366896 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1676037725
transform 1 0 372048 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1676037725
transform 1 0 377200 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1676037725
transform 1 0 382352 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1676037725
transform 1 0 387504 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1676037725
transform 1 0 392656 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1676037725
transform 1 0 397808 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1676037725
transform 1 0 402960 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1676037725
transform 1 0 408112 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1676037725
transform 1 0 413264 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1676037725
transform 1 0 418416 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1676037725
transform 1 0 423568 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1676037725
transform 1 0 428720 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1676037725
transform 1 0 433872 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1676037725
transform 1 0 439024 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1676037725
transform 1 0 444176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1676037725
transform 1 0 449328 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1676037725
transform 1 0 454480 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1676037725
transform 1 0 459632 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1676037725
transform 1 0 464784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1676037725
transform 1 0 469936 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1676037725
transform 1 0 475088 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1676037725
transform 1 0 480240 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1676037725
transform 1 0 485392 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1676037725
transform 1 0 490544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1676037725
transform 1 0 495696 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1676037725
transform 1 0 500848 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1676037725
transform 1 0 506000 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1676037725
transform 1 0 511152 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1676037725
transform 1 0 516304 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1676037725
transform 1 0 521456 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1676037725
transform 1 0 526608 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1676037725
transform 1 0 531760 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1676037725
transform 1 0 536912 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1676037725
transform 1 0 542064 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1676037725
transform 1 0 547216 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1676037725
transform 1 0 552368 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1676037725
transform 1 0 557520 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1676037725
transform 1 0 562672 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1676037725
transform 1 0 567824 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1676037725
transform 1 0 572976 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1676037725
transform 1 0 578128 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1676037725
transform 1 0 583280 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1676037725
transform 1 0 588432 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1676037725
transform 1 0 593584 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1676037725
transform 1 0 598736 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1676037725
transform 1 0 603888 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1676037725
transform 1 0 609040 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1676037725
transform 1 0 614192 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1676037725
transform 1 0 619344 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1676037725
transform 1 0 624496 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1676037725
transform 1 0 629648 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1676037725
transform 1 0 634800 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1676037725
transform 1 0 639952 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1676037725
transform 1 0 645104 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1676037725
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1676037725
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1676037725
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1676037725
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1676037725
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1676037725
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1676037725
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1676037725
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1676037725
transform 1 0 91264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1676037725
transform 1 0 96416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1676037725
transform 1 0 101568 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1676037725
transform 1 0 106720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1676037725
transform 1 0 111872 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1676037725
transform 1 0 117024 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1676037725
transform 1 0 122176 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1676037725
transform 1 0 127328 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1676037725
transform 1 0 132480 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1676037725
transform 1 0 137632 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1676037725
transform 1 0 142784 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1676037725
transform 1 0 147936 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1676037725
transform 1 0 153088 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1676037725
transform 1 0 158240 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1676037725
transform 1 0 163392 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1676037725
transform 1 0 168544 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1676037725
transform 1 0 173696 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1676037725
transform 1 0 178848 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1676037725
transform 1 0 184000 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1676037725
transform 1 0 189152 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1676037725
transform 1 0 194304 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1676037725
transform 1 0 199456 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1676037725
transform 1 0 204608 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1676037725
transform 1 0 209760 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1676037725
transform 1 0 214912 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1676037725
transform 1 0 220064 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1676037725
transform 1 0 225216 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1676037725
transform 1 0 230368 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1676037725
transform 1 0 235520 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1676037725
transform 1 0 240672 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1676037725
transform 1 0 245824 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1676037725
transform 1 0 250976 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1676037725
transform 1 0 256128 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1676037725
transform 1 0 261280 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1676037725
transform 1 0 266432 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1676037725
transform 1 0 271584 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1676037725
transform 1 0 276736 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1676037725
transform 1 0 281888 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1676037725
transform 1 0 287040 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1676037725
transform 1 0 292192 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1676037725
transform 1 0 297344 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1676037725
transform 1 0 302496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1676037725
transform 1 0 307648 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1676037725
transform 1 0 312800 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1676037725
transform 1 0 317952 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1676037725
transform 1 0 323104 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1676037725
transform 1 0 328256 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1676037725
transform 1 0 333408 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1676037725
transform 1 0 338560 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1676037725
transform 1 0 343712 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1676037725
transform 1 0 348864 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1676037725
transform 1 0 354016 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1676037725
transform 1 0 359168 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1676037725
transform 1 0 364320 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1676037725
transform 1 0 369472 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1676037725
transform 1 0 374624 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1676037725
transform 1 0 379776 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1676037725
transform 1 0 384928 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1676037725
transform 1 0 390080 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1676037725
transform 1 0 395232 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1676037725
transform 1 0 400384 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1676037725
transform 1 0 405536 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1676037725
transform 1 0 410688 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1676037725
transform 1 0 415840 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1676037725
transform 1 0 420992 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1676037725
transform 1 0 426144 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1676037725
transform 1 0 431296 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1676037725
transform 1 0 436448 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1676037725
transform 1 0 441600 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1676037725
transform 1 0 446752 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1676037725
transform 1 0 451904 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1676037725
transform 1 0 457056 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1676037725
transform 1 0 462208 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1676037725
transform 1 0 467360 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1676037725
transform 1 0 472512 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1676037725
transform 1 0 477664 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1676037725
transform 1 0 482816 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1676037725
transform 1 0 487968 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1676037725
transform 1 0 493120 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1676037725
transform 1 0 498272 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1676037725
transform 1 0 503424 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1676037725
transform 1 0 508576 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1676037725
transform 1 0 513728 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1676037725
transform 1 0 518880 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1676037725
transform 1 0 524032 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1676037725
transform 1 0 529184 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1676037725
transform 1 0 534336 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1676037725
transform 1 0 539488 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1676037725
transform 1 0 544640 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1676037725
transform 1 0 549792 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1676037725
transform 1 0 554944 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1676037725
transform 1 0 560096 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1676037725
transform 1 0 565248 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1676037725
transform 1 0 570400 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1676037725
transform 1 0 575552 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1676037725
transform 1 0 580704 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1676037725
transform 1 0 585856 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1676037725
transform 1 0 591008 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1676037725
transform 1 0 596160 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1676037725
transform 1 0 601312 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1676037725
transform 1 0 606464 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1676037725
transform 1 0 611616 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1676037725
transform 1 0 616768 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1676037725
transform 1 0 621920 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1676037725
transform 1 0 627072 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1676037725
transform 1 0 632224 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1676037725
transform 1 0 637376 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1676037725
transform 1 0 642528 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1676037725
transform 1 0 647680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1676037725
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1676037725
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1676037725
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1676037725
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1676037725
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1676037725
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1676037725
transform 1 0 83536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1676037725
transform 1 0 88688 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1676037725
transform 1 0 93840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1676037725
transform 1 0 98992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1676037725
transform 1 0 104144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1676037725
transform 1 0 109296 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1676037725
transform 1 0 114448 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1676037725
transform 1 0 119600 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1676037725
transform 1 0 124752 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1676037725
transform 1 0 129904 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1676037725
transform 1 0 135056 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1676037725
transform 1 0 140208 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1676037725
transform 1 0 145360 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1676037725
transform 1 0 150512 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1676037725
transform 1 0 155664 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1676037725
transform 1 0 160816 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1676037725
transform 1 0 165968 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1676037725
transform 1 0 171120 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1676037725
transform 1 0 176272 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1676037725
transform 1 0 181424 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1676037725
transform 1 0 186576 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1676037725
transform 1 0 191728 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1676037725
transform 1 0 196880 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1676037725
transform 1 0 202032 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1676037725
transform 1 0 207184 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1676037725
transform 1 0 212336 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1676037725
transform 1 0 217488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1676037725
transform 1 0 222640 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1676037725
transform 1 0 227792 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1676037725
transform 1 0 232944 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1676037725
transform 1 0 238096 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1676037725
transform 1 0 243248 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1676037725
transform 1 0 248400 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1676037725
transform 1 0 253552 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1676037725
transform 1 0 258704 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1676037725
transform 1 0 263856 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1676037725
transform 1 0 269008 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1676037725
transform 1 0 274160 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1676037725
transform 1 0 279312 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1676037725
transform 1 0 284464 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1676037725
transform 1 0 289616 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1676037725
transform 1 0 294768 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1676037725
transform 1 0 299920 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1676037725
transform 1 0 305072 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1676037725
transform 1 0 310224 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1676037725
transform 1 0 315376 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1676037725
transform 1 0 320528 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1676037725
transform 1 0 325680 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1676037725
transform 1 0 330832 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1676037725
transform 1 0 335984 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1676037725
transform 1 0 341136 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1676037725
transform 1 0 346288 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1676037725
transform 1 0 351440 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1676037725
transform 1 0 356592 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1676037725
transform 1 0 361744 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1676037725
transform 1 0 366896 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1676037725
transform 1 0 372048 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1676037725
transform 1 0 377200 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1676037725
transform 1 0 382352 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1676037725
transform 1 0 387504 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1676037725
transform 1 0 392656 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1676037725
transform 1 0 397808 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1676037725
transform 1 0 402960 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1676037725
transform 1 0 408112 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1676037725
transform 1 0 413264 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1676037725
transform 1 0 418416 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1676037725
transform 1 0 423568 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1676037725
transform 1 0 428720 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1676037725
transform 1 0 433872 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1676037725
transform 1 0 439024 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1676037725
transform 1 0 444176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1676037725
transform 1 0 449328 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1676037725
transform 1 0 454480 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1676037725
transform 1 0 459632 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1676037725
transform 1 0 464784 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1676037725
transform 1 0 469936 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1676037725
transform 1 0 475088 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1676037725
transform 1 0 480240 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1676037725
transform 1 0 485392 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1676037725
transform 1 0 490544 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1676037725
transform 1 0 495696 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1676037725
transform 1 0 500848 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1676037725
transform 1 0 506000 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1676037725
transform 1 0 511152 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1676037725
transform 1 0 516304 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1676037725
transform 1 0 521456 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1676037725
transform 1 0 526608 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1676037725
transform 1 0 531760 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1676037725
transform 1 0 536912 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1676037725
transform 1 0 542064 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1676037725
transform 1 0 547216 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1676037725
transform 1 0 552368 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1676037725
transform 1 0 557520 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1676037725
transform 1 0 562672 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1676037725
transform 1 0 567824 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1676037725
transform 1 0 572976 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1676037725
transform 1 0 578128 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1676037725
transform 1 0 583280 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1676037725
transform 1 0 588432 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1676037725
transform 1 0 593584 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1676037725
transform 1 0 598736 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1676037725
transform 1 0 603888 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1676037725
transform 1 0 609040 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1676037725
transform 1 0 614192 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1676037725
transform 1 0 619344 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1676037725
transform 1 0 624496 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1676037725
transform 1 0 629648 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1676037725
transform 1 0 634800 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1676037725
transform 1 0 639952 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1676037725
transform 1 0 645104 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1676037725
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1676037725
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1676037725
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1676037725
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1676037725
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1676037725
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1676037725
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1676037725
transform 1 0 86112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1676037725
transform 1 0 91264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1676037725
transform 1 0 96416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1676037725
transform 1 0 101568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1676037725
transform 1 0 106720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1676037725
transform 1 0 111872 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1676037725
transform 1 0 117024 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1676037725
transform 1 0 122176 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1676037725
transform 1 0 127328 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1676037725
transform 1 0 132480 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1676037725
transform 1 0 137632 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1676037725
transform 1 0 142784 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1676037725
transform 1 0 147936 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1676037725
transform 1 0 153088 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1676037725
transform 1 0 158240 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1676037725
transform 1 0 163392 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1676037725
transform 1 0 168544 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1676037725
transform 1 0 173696 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1676037725
transform 1 0 178848 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1676037725
transform 1 0 184000 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1676037725
transform 1 0 189152 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1676037725
transform 1 0 194304 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1676037725
transform 1 0 199456 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1676037725
transform 1 0 204608 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1676037725
transform 1 0 209760 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1676037725
transform 1 0 214912 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1676037725
transform 1 0 220064 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1676037725
transform 1 0 225216 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1676037725
transform 1 0 230368 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1676037725
transform 1 0 235520 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1676037725
transform 1 0 240672 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1676037725
transform 1 0 245824 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1676037725
transform 1 0 250976 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1676037725
transform 1 0 256128 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1676037725
transform 1 0 261280 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1676037725
transform 1 0 266432 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1676037725
transform 1 0 271584 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1676037725
transform 1 0 276736 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1676037725
transform 1 0 281888 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1676037725
transform 1 0 287040 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1676037725
transform 1 0 292192 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1676037725
transform 1 0 297344 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1676037725
transform 1 0 302496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1676037725
transform 1 0 307648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1676037725
transform 1 0 312800 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1676037725
transform 1 0 317952 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1676037725
transform 1 0 323104 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1676037725
transform 1 0 328256 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1676037725
transform 1 0 333408 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1676037725
transform 1 0 338560 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1676037725
transform 1 0 343712 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1676037725
transform 1 0 348864 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1676037725
transform 1 0 354016 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1676037725
transform 1 0 359168 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1676037725
transform 1 0 364320 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1676037725
transform 1 0 369472 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1676037725
transform 1 0 374624 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1676037725
transform 1 0 379776 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1676037725
transform 1 0 384928 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1676037725
transform 1 0 390080 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1676037725
transform 1 0 395232 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1676037725
transform 1 0 400384 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1676037725
transform 1 0 405536 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1676037725
transform 1 0 410688 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1676037725
transform 1 0 415840 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1676037725
transform 1 0 420992 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1676037725
transform 1 0 426144 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1676037725
transform 1 0 431296 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1676037725
transform 1 0 436448 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1676037725
transform 1 0 441600 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1676037725
transform 1 0 446752 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1676037725
transform 1 0 451904 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1676037725
transform 1 0 457056 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1676037725
transform 1 0 462208 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1676037725
transform 1 0 467360 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1676037725
transform 1 0 472512 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1676037725
transform 1 0 477664 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1676037725
transform 1 0 482816 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1676037725
transform 1 0 487968 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1676037725
transform 1 0 493120 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1676037725
transform 1 0 498272 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1676037725
transform 1 0 503424 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1676037725
transform 1 0 508576 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1676037725
transform 1 0 513728 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1676037725
transform 1 0 518880 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1676037725
transform 1 0 524032 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1676037725
transform 1 0 529184 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1676037725
transform 1 0 534336 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1676037725
transform 1 0 539488 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1676037725
transform 1 0 544640 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1676037725
transform 1 0 549792 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1676037725
transform 1 0 554944 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1676037725
transform 1 0 560096 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1676037725
transform 1 0 565248 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1676037725
transform 1 0 570400 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1676037725
transform 1 0 575552 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1676037725
transform 1 0 580704 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1676037725
transform 1 0 585856 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1676037725
transform 1 0 591008 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1676037725
transform 1 0 596160 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1676037725
transform 1 0 601312 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1676037725
transform 1 0 606464 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1676037725
transform 1 0 611616 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1676037725
transform 1 0 616768 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1676037725
transform 1 0 621920 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1676037725
transform 1 0 627072 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1676037725
transform 1 0 632224 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1676037725
transform 1 0 637376 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1676037725
transform 1 0 642528 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1676037725
transform 1 0 647680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1676037725
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1676037725
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1676037725
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1676037725
transform 1 0 19136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1676037725
transform 1 0 24288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1676037725
transform 1 0 29440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1676037725
transform 1 0 34592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1676037725
transform 1 0 39744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1676037725
transform 1 0 44896 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1676037725
transform 1 0 50048 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1676037725
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1676037725
transform 1 0 55200 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1676037725
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1676037725
transform 1 0 60352 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1676037725
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1676037725
transform 1 0 65504 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1676037725
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1676037725
transform 1 0 70656 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1676037725
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1676037725
transform 1 0 75808 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1676037725
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1676037725
transform 1 0 80960 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1676037725
transform 1 0 83536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1676037725
transform 1 0 86112 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1676037725
transform 1 0 88688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1676037725
transform 1 0 91264 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1676037725
transform 1 0 93840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1676037725
transform 1 0 96416 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1676037725
transform 1 0 98992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1676037725
transform 1 0 101568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1676037725
transform 1 0 104144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1676037725
transform 1 0 106720 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1676037725
transform 1 0 109296 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1676037725
transform 1 0 111872 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1676037725
transform 1 0 114448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1676037725
transform 1 0 117024 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1676037725
transform 1 0 119600 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1676037725
transform 1 0 122176 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1676037725
transform 1 0 124752 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1676037725
transform 1 0 127328 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1676037725
transform 1 0 129904 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1676037725
transform 1 0 132480 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1676037725
transform 1 0 135056 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1676037725
transform 1 0 137632 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1676037725
transform 1 0 140208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1676037725
transform 1 0 142784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1676037725
transform 1 0 145360 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1676037725
transform 1 0 147936 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1676037725
transform 1 0 150512 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1676037725
transform 1 0 153088 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1676037725
transform 1 0 155664 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1676037725
transform 1 0 158240 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1676037725
transform 1 0 160816 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1676037725
transform 1 0 163392 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1676037725
transform 1 0 165968 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1676037725
transform 1 0 168544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1676037725
transform 1 0 171120 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1676037725
transform 1 0 173696 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1676037725
transform 1 0 176272 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1676037725
transform 1 0 178848 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1676037725
transform 1 0 181424 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1676037725
transform 1 0 184000 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1676037725
transform 1 0 186576 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1676037725
transform 1 0 189152 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1676037725
transform 1 0 191728 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1676037725
transform 1 0 194304 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1676037725
transform 1 0 196880 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1676037725
transform 1 0 199456 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1676037725
transform 1 0 202032 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1676037725
transform 1 0 204608 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1676037725
transform 1 0 207184 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1676037725
transform 1 0 209760 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1676037725
transform 1 0 212336 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1676037725
transform 1 0 214912 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1676037725
transform 1 0 217488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1676037725
transform 1 0 220064 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1676037725
transform 1 0 222640 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1676037725
transform 1 0 225216 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1676037725
transform 1 0 227792 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1676037725
transform 1 0 230368 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1676037725
transform 1 0 232944 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1676037725
transform 1 0 235520 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1676037725
transform 1 0 238096 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1676037725
transform 1 0 240672 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1676037725
transform 1 0 243248 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1676037725
transform 1 0 245824 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1676037725
transform 1 0 248400 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1676037725
transform 1 0 250976 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1676037725
transform 1 0 253552 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1676037725
transform 1 0 256128 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1676037725
transform 1 0 258704 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1676037725
transform 1 0 261280 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1676037725
transform 1 0 263856 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1676037725
transform 1 0 266432 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1676037725
transform 1 0 269008 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1676037725
transform 1 0 271584 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1676037725
transform 1 0 274160 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1676037725
transform 1 0 276736 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1676037725
transform 1 0 279312 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1676037725
transform 1 0 281888 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1676037725
transform 1 0 284464 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1676037725
transform 1 0 287040 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1676037725
transform 1 0 289616 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1676037725
transform 1 0 292192 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1676037725
transform 1 0 294768 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1676037725
transform 1 0 297344 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1676037725
transform 1 0 299920 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1676037725
transform 1 0 302496 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1676037725
transform 1 0 305072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1676037725
transform 1 0 307648 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1676037725
transform 1 0 310224 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1676037725
transform 1 0 312800 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1676037725
transform 1 0 315376 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1676037725
transform 1 0 317952 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1676037725
transform 1 0 320528 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1676037725
transform 1 0 323104 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1676037725
transform 1 0 325680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1676037725
transform 1 0 328256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1676037725
transform 1 0 330832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1676037725
transform 1 0 333408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1676037725
transform 1 0 335984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1676037725
transform 1 0 338560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1676037725
transform 1 0 341136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1676037725
transform 1 0 343712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1676037725
transform 1 0 346288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1676037725
transform 1 0 348864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1676037725
transform 1 0 351440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1676037725
transform 1 0 354016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1676037725
transform 1 0 356592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1676037725
transform 1 0 359168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1676037725
transform 1 0 361744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1676037725
transform 1 0 364320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1676037725
transform 1 0 366896 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1676037725
transform 1 0 369472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1676037725
transform 1 0 372048 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1676037725
transform 1 0 374624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1676037725
transform 1 0 377200 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1676037725
transform 1 0 379776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1676037725
transform 1 0 382352 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1676037725
transform 1 0 384928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1676037725
transform 1 0 387504 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1676037725
transform 1 0 390080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1676037725
transform 1 0 392656 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1676037725
transform 1 0 395232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1676037725
transform 1 0 397808 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1676037725
transform 1 0 400384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1676037725
transform 1 0 402960 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1676037725
transform 1 0 405536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1676037725
transform 1 0 408112 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1676037725
transform 1 0 410688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1676037725
transform 1 0 413264 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1676037725
transform 1 0 415840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1676037725
transform 1 0 418416 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1676037725
transform 1 0 420992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1676037725
transform 1 0 423568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1439
timestamp 1676037725
transform 1 0 426144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1440
timestamp 1676037725
transform 1 0 428720 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1441
timestamp 1676037725
transform 1 0 431296 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1442
timestamp 1676037725
transform 1 0 433872 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1443
timestamp 1676037725
transform 1 0 436448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1444
timestamp 1676037725
transform 1 0 439024 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1445
timestamp 1676037725
transform 1 0 441600 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1446
timestamp 1676037725
transform 1 0 444176 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1447
timestamp 1676037725
transform 1 0 446752 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1448
timestamp 1676037725
transform 1 0 449328 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1449
timestamp 1676037725
transform 1 0 451904 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1450
timestamp 1676037725
transform 1 0 454480 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1451
timestamp 1676037725
transform 1 0 457056 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1452
timestamp 1676037725
transform 1 0 459632 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1453
timestamp 1676037725
transform 1 0 462208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1454
timestamp 1676037725
transform 1 0 464784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1455
timestamp 1676037725
transform 1 0 467360 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1456
timestamp 1676037725
transform 1 0 469936 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1457
timestamp 1676037725
transform 1 0 472512 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1458
timestamp 1676037725
transform 1 0 475088 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1459
timestamp 1676037725
transform 1 0 477664 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1460
timestamp 1676037725
transform 1 0 480240 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1461
timestamp 1676037725
transform 1 0 482816 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1462
timestamp 1676037725
transform 1 0 485392 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1463
timestamp 1676037725
transform 1 0 487968 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1464
timestamp 1676037725
transform 1 0 490544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1465
timestamp 1676037725
transform 1 0 493120 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1466
timestamp 1676037725
transform 1 0 495696 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1467
timestamp 1676037725
transform 1 0 498272 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1468
timestamp 1676037725
transform 1 0 500848 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1469
timestamp 1676037725
transform 1 0 503424 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1470
timestamp 1676037725
transform 1 0 506000 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1471
timestamp 1676037725
transform 1 0 508576 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1472
timestamp 1676037725
transform 1 0 511152 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1473
timestamp 1676037725
transform 1 0 513728 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1474
timestamp 1676037725
transform 1 0 516304 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1475
timestamp 1676037725
transform 1 0 518880 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1476
timestamp 1676037725
transform 1 0 521456 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1477
timestamp 1676037725
transform 1 0 524032 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1478
timestamp 1676037725
transform 1 0 526608 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1479
timestamp 1676037725
transform 1 0 529184 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1480
timestamp 1676037725
transform 1 0 531760 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1481
timestamp 1676037725
transform 1 0 534336 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1482
timestamp 1676037725
transform 1 0 536912 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1483
timestamp 1676037725
transform 1 0 539488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1484
timestamp 1676037725
transform 1 0 542064 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1485
timestamp 1676037725
transform 1 0 544640 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1486
timestamp 1676037725
transform 1 0 547216 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1487
timestamp 1676037725
transform 1 0 549792 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1488
timestamp 1676037725
transform 1 0 552368 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1489
timestamp 1676037725
transform 1 0 554944 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1490
timestamp 1676037725
transform 1 0 557520 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1491
timestamp 1676037725
transform 1 0 560096 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1492
timestamp 1676037725
transform 1 0 562672 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1493
timestamp 1676037725
transform 1 0 565248 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1494
timestamp 1676037725
transform 1 0 567824 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1495
timestamp 1676037725
transform 1 0 570400 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1496
timestamp 1676037725
transform 1 0 572976 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1497
timestamp 1676037725
transform 1 0 575552 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1498
timestamp 1676037725
transform 1 0 578128 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1499
timestamp 1676037725
transform 1 0 580704 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1500
timestamp 1676037725
transform 1 0 583280 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1501
timestamp 1676037725
transform 1 0 585856 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1502
timestamp 1676037725
transform 1 0 588432 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1503
timestamp 1676037725
transform 1 0 591008 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1504
timestamp 1676037725
transform 1 0 593584 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1505
timestamp 1676037725
transform 1 0 596160 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1506
timestamp 1676037725
transform 1 0 598736 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1507
timestamp 1676037725
transform 1 0 601312 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1508
timestamp 1676037725
transform 1 0 603888 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1509
timestamp 1676037725
transform 1 0 606464 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1510
timestamp 1676037725
transform 1 0 609040 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1511
timestamp 1676037725
transform 1 0 611616 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1512
timestamp 1676037725
transform 1 0 614192 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1513
timestamp 1676037725
transform 1 0 616768 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1514
timestamp 1676037725
transform 1 0 619344 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1515
timestamp 1676037725
transform 1 0 621920 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1516
timestamp 1676037725
transform 1 0 624496 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1517
timestamp 1676037725
transform 1 0 627072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1518
timestamp 1676037725
transform 1 0 629648 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1519
timestamp 1676037725
transform 1 0 632224 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1520
timestamp 1676037725
transform 1 0 634800 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1521
timestamp 1676037725
transform 1 0 637376 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1522
timestamp 1676037725
transform 1 0 639952 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1523
timestamp 1676037725
transform 1 0 642528 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1524
timestamp 1676037725
transform 1 0 645104 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1525
timestamp 1676037725
transform 1 0 647680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  u_rp\[0\].u_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[1\].u_buf
timestamp 1676037725
transform -1 0 17572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[2\].u_buf
timestamp 1676037725
transform -1 0 33028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[3\].u_buf
timestamp 1676037725
transform -1 0 48484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[4\].u_buf
timestamp 1676037725
transform -1 0 63940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[5\].u_buf
timestamp 1676037725
transform -1 0 79396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[6\].u_buf
timestamp 1676037725
transform -1 0 94852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[7\].u_buf
timestamp 1676037725
transform -1 0 110308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[8\].u_buf
timestamp 1676037725
transform -1 0 125764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[9\].u_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 141220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[10\].u_buf
timestamp 1676037725
transform -1 0 156676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[11\].u_buf
timestamp 1676037725
transform -1 0 172132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[12\].u_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 187588 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[13\].u_buf
timestamp 1676037725
transform -1 0 203044 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[14\].u_buf
timestamp 1676037725
transform -1 0 218500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[15\].u_buf
timestamp 1676037725
transform -1 0 233956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[16\].u_buf
timestamp 1676037725
transform -1 0 249412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[17\].u_buf
timestamp 1676037725
transform -1 0 264868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[18\].u_buf
timestamp 1676037725
transform -1 0 280324 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[19\].u_buf
timestamp 1676037725
transform -1 0 295780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[20\].u_buf
timestamp 1676037725
transform -1 0 311236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[21\].u_buf
timestamp 1676037725
transform -1 0 326692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[22\].u_buf
timestamp 1676037725
transform -1 0 342148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[23\].u_buf
timestamp 1676037725
transform -1 0 357604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[24\].u_buf
timestamp 1676037725
transform -1 0 373060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[25\].u_buf
timestamp 1676037725
transform -1 0 388516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[26\].u_buf
timestamp 1676037725
transform -1 0 403972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  u_rp\[27\].u_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 419428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  u_rp\[28\].u_buf
timestamp 1676037725
transform -1 0 434884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[29\].u_buf
timestamp 1676037725
transform -1 0 450340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[30\].u_buf
timestamp 1676037725
transform -1 0 465796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[31\].u_buf
timestamp 1676037725
transform -1 0 481252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[32\].u_buf
timestamp 1676037725
transform -1 0 496708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  u_rp\[33\].u_buf
timestamp 1676037725
transform -1 0 512164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  u_rp\[34\].u_buf
timestamp 1676037725
transform -1 0 527620 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[35\].u_buf
timestamp 1676037725
transform -1 0 543076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[36\].u_buf
timestamp 1676037725
transform -1 0 558532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[37\].u_buf
timestamp 1676037725
transform -1 0 573988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[38\].u_buf
timestamp 1676037725
transform -1 0 589444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  u_rp\[39\].u_buf
timestamp 1676037725
transform -1 0 604900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  u_rp\[40\].u_buf
timestamp 1676037725
transform -1 0 620356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[41\].u_buf
timestamp 1676037725
transform -1 0 635812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  wire1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 112700 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 125396 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  wire3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 219788 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  wire4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 313260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  wire5
timestamp 1676037725
transform -1 0 406824 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire6
timestamp 1676037725
transform -1 0 500664 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire7
timestamp 1676037725
transform -1 0 594412 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire8
timestamp 1676037725
transform -1 0 124200 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  wire9
timestamp 1676037725
transform -1 0 218776 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  wire10
timestamp 1676037725
transform -1 0 311788 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  wire11
timestamp 1676037725
transform -1 0 405352 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire12
timestamp 1676037725
transform -1 0 499376 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire13
timestamp 1676037725
transform -1 0 123372 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  wire14
timestamp 1676037725
transform -1 0 217304 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  wire15
timestamp 1676037725
transform -1 0 310960 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  wire16
timestamp 1676037725
transform -1 0 404340 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire17
timestamp 1676037725
transform -1 0 497628 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire18
timestamp 1676037725
transform -1 0 121992 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire19
timestamp 1676037725
transform -1 0 216016 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire20
timestamp 1676037725
transform -1 0 309488 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire21
timestamp 1676037725
transform -1 0 402960 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire22
timestamp 1676037725
transform -1 0 121532 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire23
timestamp 1676037725
transform -1 0 214820 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire24
timestamp 1676037725
transform -1 0 308752 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire25
timestamp 1676037725
transform -1 0 401120 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire26
timestamp 1676037725
transform -1 0 120336 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire27
timestamp 1676037725
transform -1 0 213624 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire28
timestamp 1676037725
transform -1 0 306636 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire29
timestamp 1676037725
transform -1 0 119416 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire30
timestamp 1676037725
transform -1 0 212244 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire31
timestamp 1676037725
transform -1 0 304704 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire32
timestamp 1676037725
transform -1 0 117944 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire33
timestamp 1676037725
transform -1 0 210864 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire34
timestamp 1676037725
transform -1 0 116840 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire35
timestamp 1676037725
transform -1 0 208472 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire36
timestamp 1676037725
transform -1 0 115184 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire37
timestamp 1676037725
transform 1 0 37444 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  wire38
timestamp 1676037725
transform 1 0 541880 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  wire39
timestamp 1676037725
transform 1 0 447948 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  wire40
timestamp 1676037725
transform 1 0 354108 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire41
timestamp 1676037725
transform 1 0 260268 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire42
timestamp 1676037725
transform 1 0 166336 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire43
timestamp 1676037725
transform 1 0 72496 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  wire44
timestamp 1676037725
transform 1 0 526884 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  wire45
timestamp 1676037725
transform 1 0 432584 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  wire46
timestamp 1676037725
transform 1 0 338744 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire47
timestamp 1676037725
transform 1 0 244812 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire48
timestamp 1676037725
transform 1 0 151064 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire49
timestamp 1676037725
transform 1 0 57040 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  wire50
timestamp 1676037725
transform 1 0 495972 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  wire51
timestamp 1676037725
transform 1 0 401672 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  wire52
timestamp 1676037725
transform 1 0 308016 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire53
timestamp 1676037725
transform 1 0 213900 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire54
timestamp 1676037725
transform 1 0 119968 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  wire55
timestamp 1676037725
transform 1 0 480516 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  wire56
timestamp 1676037725
transform 1 0 386216 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  wire57
timestamp 1676037725
transform 1 0 292652 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire58
timestamp 1676037725
transform 1 0 198444 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire59
timestamp 1676037725
transform 1 0 105156 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  wire60
timestamp 1676037725
transform 1 0 449604 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  wire61
timestamp 1676037725
transform 1 0 355304 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  wire62
timestamp 1676037725
transform 1 0 261924 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire63
timestamp 1676037725
transform 1 0 168820 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire64
timestamp 1676037725
transform 1 0 74612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  wire65
timestamp 1676037725
transform 1 0 434148 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  wire66
timestamp 1676037725
transform 1 0 339848 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  wire67
timestamp 1676037725
transform 1 0 246652 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire68
timestamp 1676037725
transform 1 0 153364 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire69
timestamp 1676037725
transform 1 0 59340 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  wire70
timestamp 1676037725
transform 1 0 403236 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  wire71
timestamp 1676037725
transform 1 0 309488 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  wire72
timestamp 1676037725
transform 1 0 215924 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire73
timestamp 1676037725
transform 1 0 122452 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  wire74
timestamp 1676037725
transform 1 0 387780 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  wire75
timestamp 1676037725
transform 1 0 294216 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  wire76
timestamp 1676037725
transform 1 0 200652 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire77
timestamp 1676037725
transform 1 0 107180 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  wire78
timestamp 1676037725
transform 1 0 356868 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  wire79
timestamp 1676037725
transform 1 0 263488 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  wire80
timestamp 1676037725
transform 1 0 170016 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire81
timestamp 1676037725
transform 1 0 76636 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  wire82
timestamp 1676037725
transform 1 0 341504 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  wire83
timestamp 1676037725
transform 1 0 248124 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  wire84
timestamp 1676037725
transform 1 0 154652 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire85
timestamp 1676037725
transform 1 0 61456 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire86
timestamp 1676037725
transform 1 0 310960 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire87
timestamp 1676037725
transform 1 0 217764 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire88
timestamp 1676037725
transform 1 0 123740 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire89
timestamp 1676037725
transform 1 0 295320 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire90
timestamp 1676037725
transform 1 0 202308 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire91
timestamp 1676037725
transform 1 0 109020 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire92
timestamp 1676037725
transform 1 0 264592 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire93
timestamp 1676037725
transform 1 0 171580 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire94
timestamp 1676037725
transform 1 0 78660 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire95
timestamp 1676037725
transform 1 0 249228 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire96
timestamp 1676037725
transform 1 0 156308 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire97
timestamp 1676037725
transform 1 0 63480 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire98
timestamp 1676037725
transform 1 0 218500 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire99
timestamp 1676037725
transform 1 0 125856 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire100
timestamp 1676037725
transform 1 0 33212 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire101
timestamp 1676037725
transform 1 0 203228 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire102
timestamp 1676037725
transform 1 0 110676 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire103
timestamp 1676037725
transform 1 0 172592 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire104
timestamp 1676037725
transform 1 0 79948 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire105
timestamp 1676037725
transform 1 0 157228 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire106
timestamp 1676037725
transform 1 0 64768 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire107
timestamp 1676037725
transform 1 0 126868 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire108
timestamp 1676037725
transform 1 0 35236 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire109
timestamp 1676037725
transform 1 0 111688 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire110
timestamp 1676037725
transform 1 0 81420 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire111
timestamp 1676037725
transform 1 0 66424 0 -1 7616
box -38 -48 590 592
<< labels >>
flabel metal1 s 74 0 130 800 0 FreeSans 224 90 0 0 ch_in[0]
port 0 nsew signal input
flabel metal1 s 22786 9200 22842 10000 0 FreeSans 224 90 0 0 ch_in[10]
port 1 nsew signal input
flabel metal1 s 23058 9200 23114 10000 0 FreeSans 224 90 0 0 ch_in[11]
port 2 nsew signal input
flabel metal1 s 183674 0 183730 800 0 FreeSans 224 90 0 0 ch_in[12]
port 3 nsew signal input
flabel metal1 s 23602 9200 23658 10000 0 FreeSans 224 90 0 0 ch_in[13]
port 4 nsew signal input
flabel metal1 s 23874 9200 23930 10000 0 FreeSans 224 90 0 0 ch_in[14]
port 5 nsew signal input
flabel metal1 s 229574 0 229630 800 0 FreeSans 224 90 0 0 ch_in[15]
port 6 nsew signal input
flabel metal1 s 24418 9200 24474 10000 0 FreeSans 224 90 0 0 ch_in[16]
port 7 nsew signal input
flabel metal1 s 24690 9200 24746 10000 0 FreeSans 224 90 0 0 ch_in[17]
port 8 nsew signal input
flabel metal1 s 275474 0 275530 800 0 FreeSans 224 90 0 0 ch_in[18]
port 9 nsew signal input
flabel metal1 s 25234 9200 25290 10000 0 FreeSans 224 90 0 0 ch_in[19]
port 10 nsew signal input
flabel metal1 s 20338 9200 20394 10000 0 FreeSans 224 90 0 0 ch_in[1]
port 11 nsew signal input
flabel metal1 s 25506 9200 25562 10000 0 FreeSans 224 90 0 0 ch_in[20]
port 12 nsew signal input
flabel metal1 s 321374 0 321430 800 0 FreeSans 224 90 0 0 ch_in[21]
port 13 nsew signal input
flabel metal1 s 26050 9200 26106 10000 0 FreeSans 224 90 0 0 ch_in[22]
port 14 nsew signal input
flabel metal1 s 26322 9200 26378 10000 0 FreeSans 224 90 0 0 ch_in[23]
port 15 nsew signal input
flabel metal1 s 367274 0 367330 800 0 FreeSans 224 90 0 0 ch_in[24]
port 16 nsew signal input
flabel metal1 s 26866 9200 26922 10000 0 FreeSans 224 90 0 0 ch_in[25]
port 17 nsew signal input
flabel metal1 s 27138 9200 27194 10000 0 FreeSans 224 90 0 0 ch_in[26]
port 18 nsew signal input
flabel metal1 s 413174 0 413230 800 0 FreeSans 224 90 0 0 ch_in[27]
port 19 nsew signal input
flabel metal1 s 27682 9200 27738 10000 0 FreeSans 224 90 0 0 ch_in[28]
port 20 nsew signal input
flabel metal1 s 27954 9200 28010 10000 0 FreeSans 224 90 0 0 ch_in[29]
port 21 nsew signal input
flabel metal1 s 20610 9200 20666 10000 0 FreeSans 224 90 0 0 ch_in[2]
port 22 nsew signal input
flabel metal1 s 459074 0 459130 800 0 FreeSans 224 90 0 0 ch_in[30]
port 23 nsew signal input
flabel metal1 s 28498 9200 28554 10000 0 FreeSans 224 90 0 0 ch_in[31]
port 24 nsew signal input
flabel metal1 s 28770 9200 28826 10000 0 FreeSans 224 90 0 0 ch_in[32]
port 25 nsew signal input
flabel metal1 s 504974 0 505030 800 0 FreeSans 224 90 0 0 ch_in[33]
port 26 nsew signal input
flabel metal1 s 29314 9200 29370 10000 0 FreeSans 224 90 0 0 ch_in[34]
port 27 nsew signal input
flabel metal1 s 29586 9200 29642 10000 0 FreeSans 224 90 0 0 ch_in[35]
port 28 nsew signal input
flabel metal1 s 550874 0 550930 800 0 FreeSans 224 90 0 0 ch_in[36]
port 29 nsew signal input
flabel metal1 s 30130 9200 30186 10000 0 FreeSans 224 90 0 0 ch_in[37]
port 30 nsew signal input
flabel metal1 s 30402 9200 30458 10000 0 FreeSans 224 90 0 0 ch_in[38]
port 31 nsew signal input
flabel metal1 s 596774 0 596830 800 0 FreeSans 224 90 0 0 ch_in[39]
port 32 nsew signal input
flabel metal1 s 45974 0 46030 800 0 FreeSans 224 90 0 0 ch_in[3]
port 33 nsew signal input
flabel metal1 s 30946 9200 31002 10000 0 FreeSans 224 90 0 0 ch_in[40]
port 34 nsew signal input
flabel metal1 s 31218 9200 31274 10000 0 FreeSans 224 90 0 0 ch_in[41]
port 35 nsew signal input
flabel metal1 s 21154 9200 21210 10000 0 FreeSans 224 90 0 0 ch_in[4]
port 36 nsew signal input
flabel metal1 s 21426 9200 21482 10000 0 FreeSans 224 90 0 0 ch_in[5]
port 37 nsew signal input
flabel metal1 s 91874 0 91930 800 0 FreeSans 224 90 0 0 ch_in[6]
port 38 nsew signal input
flabel metal1 s 21970 9200 22026 10000 0 FreeSans 224 90 0 0 ch_in[7]
port 39 nsew signal input
flabel metal1 s 22242 9200 22298 10000 0 FreeSans 224 90 0 0 ch_in[8]
port 40 nsew signal input
flabel metal1 s 137774 0 137830 800 0 FreeSans 224 90 0 0 ch_in[9]
port 41 nsew signal input
flabel metal1 s 20066 9200 20122 10000 0 FreeSans 224 90 0 0 ch_out[0]
port 42 nsew signal tristate
flabel metal1 s 153074 0 153130 800 0 FreeSans 224 90 0 0 ch_out[10]
port 43 nsew signal tristate
flabel metal1 s 168374 0 168430 800 0 FreeSans 224 90 0 0 ch_out[11]
port 44 nsew signal tristate
flabel metal1 s 23330 9200 23386 10000 0 FreeSans 224 90 0 0 ch_out[12]
port 45 nsew signal tristate
flabel metal1 s 198974 0 199030 800 0 FreeSans 224 90 0 0 ch_out[13]
port 46 nsew signal tristate
flabel metal1 s 214274 0 214330 800 0 FreeSans 224 90 0 0 ch_out[14]
port 47 nsew signal tristate
flabel metal1 s 24146 9200 24202 10000 0 FreeSans 224 90 0 0 ch_out[15]
port 48 nsew signal tristate
flabel metal1 s 244874 0 244930 800 0 FreeSans 224 90 0 0 ch_out[16]
port 49 nsew signal tristate
flabel metal1 s 260174 0 260230 800 0 FreeSans 224 90 0 0 ch_out[17]
port 50 nsew signal tristate
flabel metal1 s 24962 9200 25018 10000 0 FreeSans 224 90 0 0 ch_out[18]
port 51 nsew signal tristate
flabel metal1 s 290774 0 290830 800 0 FreeSans 224 90 0 0 ch_out[19]
port 52 nsew signal tristate
flabel metal1 s 15374 0 15430 800 0 FreeSans 224 90 0 0 ch_out[1]
port 53 nsew signal tristate
flabel metal1 s 306074 0 306130 800 0 FreeSans 224 90 0 0 ch_out[20]
port 54 nsew signal tristate
flabel metal1 s 25778 9200 25834 10000 0 FreeSans 224 90 0 0 ch_out[21]
port 55 nsew signal tristate
flabel metal1 s 336674 0 336730 800 0 FreeSans 224 90 0 0 ch_out[22]
port 56 nsew signal tristate
flabel metal1 s 351974 0 352030 800 0 FreeSans 224 90 0 0 ch_out[23]
port 57 nsew signal tristate
flabel metal1 s 26594 9200 26650 10000 0 FreeSans 224 90 0 0 ch_out[24]
port 58 nsew signal tristate
flabel metal1 s 382574 0 382630 800 0 FreeSans 224 90 0 0 ch_out[25]
port 59 nsew signal tristate
flabel metal1 s 397874 0 397930 800 0 FreeSans 224 90 0 0 ch_out[26]
port 60 nsew signal tristate
flabel metal1 s 27410 9200 27466 10000 0 FreeSans 224 90 0 0 ch_out[27]
port 61 nsew signal tristate
flabel metal1 s 428474 0 428530 800 0 FreeSans 224 90 0 0 ch_out[28]
port 62 nsew signal tristate
flabel metal1 s 443774 0 443830 800 0 FreeSans 224 90 0 0 ch_out[29]
port 63 nsew signal tristate
flabel metal1 s 30674 0 30730 800 0 FreeSans 224 90 0 0 ch_out[2]
port 64 nsew signal tristate
flabel metal1 s 28226 9200 28282 10000 0 FreeSans 224 90 0 0 ch_out[30]
port 65 nsew signal tristate
flabel metal1 s 474374 0 474430 800 0 FreeSans 224 90 0 0 ch_out[31]
port 66 nsew signal tristate
flabel metal1 s 489674 0 489730 800 0 FreeSans 224 90 0 0 ch_out[32]
port 67 nsew signal tristate
flabel metal1 s 29042 9200 29098 10000 0 FreeSans 224 90 0 0 ch_out[33]
port 68 nsew signal tristate
flabel metal1 s 520274 0 520330 800 0 FreeSans 224 90 0 0 ch_out[34]
port 69 nsew signal tristate
flabel metal1 s 535574 0 535630 800 0 FreeSans 224 90 0 0 ch_out[35]
port 70 nsew signal tristate
flabel metal1 s 29858 9200 29914 10000 0 FreeSans 224 90 0 0 ch_out[36]
port 71 nsew signal tristate
flabel metal1 s 566174 0 566230 800 0 FreeSans 224 90 0 0 ch_out[37]
port 72 nsew signal tristate
flabel metal1 s 581474 0 581530 800 0 FreeSans 224 90 0 0 ch_out[38]
port 73 nsew signal tristate
flabel metal1 s 30674 9200 30730 10000 0 FreeSans 224 90 0 0 ch_out[39]
port 74 nsew signal tristate
flabel metal1 s 20882 9200 20938 10000 0 FreeSans 224 90 0 0 ch_out[3]
port 75 nsew signal tristate
flabel metal1 s 612074 0 612130 800 0 FreeSans 224 90 0 0 ch_out[40]
port 76 nsew signal tristate
flabel metal1 s 627374 0 627430 800 0 FreeSans 224 90 0 0 ch_out[41]
port 77 nsew signal tristate
flabel metal1 s 61274 0 61330 800 0 FreeSans 224 90 0 0 ch_out[4]
port 78 nsew signal tristate
flabel metal1 s 76574 0 76630 800 0 FreeSans 224 90 0 0 ch_out[5]
port 79 nsew signal tristate
flabel metal1 s 21698 9200 21754 10000 0 FreeSans 224 90 0 0 ch_out[6]
port 80 nsew signal tristate
flabel metal1 s 107174 0 107230 800 0 FreeSans 224 90 0 0 ch_out[7]
port 81 nsew signal tristate
flabel metal1 s 122474 0 122530 800 0 FreeSans 224 90 0 0 ch_out[8]
port 82 nsew signal tristate
flabel metal1 s 22514 9200 22570 10000 0 FreeSans 224 90 0 0 ch_out[9]
port 83 nsew signal tristate
flabel metal2 s -416 656 -96 9136 0 FreeSans 1792 90 0 0 vccd1
port 84 nsew power bidirectional
flabel metal3 s -416 656 650396 976 0 FreeSans 1920 0 0 0 vccd1
port 84 nsew power bidirectional
flabel metal3 s -416 8816 650396 9136 0 FreeSans 1920 0 0 0 vccd1
port 84 nsew power bidirectional
flabel metal2 s 650076 656 650396 9136 0 FreeSans 1792 90 0 0 vccd1
port 84 nsew power bidirectional
flabel metal2 s 81915 -4 82235 9796 0 FreeSans 1792 90 0 0 vccd1
port 84 nsew power bidirectional
flabel metal2 s 243858 -4 244178 9796 0 FreeSans 1792 90 0 0 vccd1
port 84 nsew power bidirectional
flabel metal2 s 405801 -4 406121 9796 0 FreeSans 1792 90 0 0 vccd1
port 84 nsew power bidirectional
flabel metal2 s 567744 -4 568064 9796 0 FreeSans 1792 90 0 0 vccd1
port 84 nsew power bidirectional
flabel metal3 s -1076 2695 651056 3015 0 FreeSans 1920 0 0 0 vccd1
port 84 nsew power bidirectional
flabel metal3 s -1076 4054 651056 4374 0 FreeSans 1920 0 0 0 vccd1
port 84 nsew power bidirectional
flabel metal3 s -1076 5413 651056 5733 0 FreeSans 1920 0 0 0 vccd1
port 84 nsew power bidirectional
flabel metal3 s -1076 6772 651056 7092 0 FreeSans 1920 0 0 0 vccd1
port 84 nsew power bidirectional
flabel metal2 s -1076 -4 -756 9796 0 FreeSans 1792 90 0 0 vssd1
port 85 nsew ground bidirectional
flabel metal3 s -1076 -4 651056 316 0 FreeSans 1920 0 0 0 vssd1
port 85 nsew ground bidirectional
flabel metal3 s -1076 9476 651056 9796 0 FreeSans 1920 0 0 0 vssd1
port 85 nsew ground bidirectional
flabel metal2 s 650736 -4 651056 9796 0 FreeSans 1792 90 0 0 vssd1
port 85 nsew ground bidirectional
flabel metal2 s 82575 -4 82895 9796 0 FreeSans 1792 90 0 0 vssd1
port 85 nsew ground bidirectional
flabel metal2 s 244518 -4 244838 9796 0 FreeSans 1792 90 0 0 vssd1
port 85 nsew ground bidirectional
flabel metal2 s 406461 -4 406781 9796 0 FreeSans 1792 90 0 0 vssd1
port 85 nsew ground bidirectional
flabel metal2 s 568404 -4 568724 9796 0 FreeSans 1792 90 0 0 vssd1
port 85 nsew ground bidirectional
flabel metal3 s -1076 3355 651056 3675 0 FreeSans 1920 0 0 0 vssd1
port 85 nsew ground bidirectional
flabel metal3 s -1076 4714 651056 5034 0 FreeSans 1920 0 0 0 vssd1
port 85 nsew ground bidirectional
flabel metal3 s -1076 6073 651056 6393 0 FreeSans 1920 0 0 0 vssd1
port 85 nsew ground bidirectional
flabel metal3 s -1076 7432 651056 7752 0 FreeSans 1920 0 0 0 vssd1
port 85 nsew ground bidirectional
rlabel metal1 324990 7072 324990 7072 0 vccd1
rlabel metal1 324990 7616 324990 7616 0 vssd1
rlabel metal2 1610 1802 1610 1802 0 ch_in[0]
rlabel metal2 65918 7752 65918 7752 0 ch_in[10]
rlabel metal2 81558 6426 81558 6426 0 ch_in[11]
rlabel metal2 186898 1802 186898 1802 0 ch_in[12]
rlabel metal1 111504 6290 111504 6290 0 ch_in[13]
rlabel metal2 35282 7990 35282 7990 0 ch_in[14]
rlabel metal2 233818 1564 233818 1564 0 ch_in[15]
rlabel metal2 64814 7140 64814 7140 0 ch_in[16]
rlabel metal1 79718 6766 79718 6766 0 ch_in[17]
rlabel metal2 279634 1802 279634 1802 0 ch_in[18]
rlabel metal2 110170 8228 110170 8228 0 ch_in[19]
rlabel metal2 18078 4692 18078 4692 0 ch_in[1]
rlabel metal2 32706 7922 32706 7922 0 ch_in[20]
rlabel metal2 326554 1564 326554 1564 0 ch_in[21]
rlabel metal1 63204 6766 63204 6766 0 ch_in[22]
rlabel metal2 78062 8092 78062 8092 0 ch_in[23]
rlabel metal2 372646 1802 372646 1802 0 ch_in[24]
rlabel metal1 108836 6766 108836 6766 0 ch_in[25]
rlabel metal2 27278 8806 27278 8806 0 ch_in[26]
rlabel metal1 418646 2414 418646 2414 0 ch_in[27]
rlabel metal2 60950 7582 60950 7582 0 ch_in[28]
rlabel metal2 76130 7718 76130 7718 0 ch_in[29]
rlabel via1 20646 8874 20646 8874 0 ch_in[2]
rlabel metal2 465290 1428 465290 1428 0 ch_in[30]
rlabel metal2 107318 8160 107318 8160 0 ch_in[31]
rlabel metal2 28934 7378 28934 7378 0 ch_in[32]
rlabel metal2 511934 1598 511934 1598 0 ch_in[33]
rlabel metal1 59110 7378 59110 7378 0 ch_in[34]
rlabel metal2 74106 8058 74106 8058 0 ch_in[35]
rlabel metal2 558026 1802 558026 1802 0 ch_in[36]
rlabel metal2 104650 8126 104650 8126 0 ch_in[37]
rlabel metal1 30590 9180 30590 9180 0 ch_in[38]
rlabel metal1 604532 2414 604532 2414 0 ch_in[39]
rlabel metal2 47978 1802 47978 1802 0 ch_in[3]
rlabel metal2 56626 7650 56626 7650 0 ch_in[40]
rlabel metal2 71990 7548 71990 7548 0 ch_in[41]
rlabel metal2 63894 2652 63894 2652 0 ch_in[4]
rlabel metal2 79350 2686 79350 2686 0 ch_in[5]
rlabel metal2 94346 1802 94346 1802 0 ch_in[6]
rlabel via1 22011 8942 22011 8942 0 ch_in[7]
rlabel metal2 36846 7990 36846 7990 0 ch_in[8]
rlabel metal2 141082 1564 141082 1564 0 ch_in[9]
rlabel metal2 17894 4590 17894 4590 0 ch_out[0]
rlabel metal1 154774 782 154774 782 0 ch_out[10]
rlabel metal1 169057 782 169057 782 0 ch_out[11]
rlabel metal2 23414 7378 23414 7378 0 ch_out[12]
rlabel metal1 199256 782 199256 782 0 ch_out[13]
rlabel metal1 216299 782 216299 782 0 ch_out[14]
rlabel metal2 116150 6290 116150 6290 0 ch_out[15]
rlabel metal2 249182 1530 249182 1530 0 ch_out[16]
rlabel metal1 262427 782 262427 782 0 ch_out[17]
rlabel metal1 117622 7480 117622 7480 0 ch_out[18]
rlabel metal1 292406 782 292406 782 0 ch_out[19]
rlabel metal1 15693 782 15693 782 0 ch_out[1]
rlabel metal2 309166 1156 309166 1156 0 ch_out[20]
rlabel metal1 107778 7412 107778 7412 0 ch_out[21]
rlabel metal1 338121 782 338121 782 0 ch_out[22]
rlabel metal2 357374 1530 357374 1530 0 ch_out[23]
rlabel metal2 26726 8024 26726 8024 0 ch_out[24]
rlabel metal2 386446 1156 386446 1156 0 ch_out[25]
rlabel metal1 400322 782 400322 782 0 ch_out[26]
rlabel metal1 103500 6256 103500 6256 0 ch_out[27]
rlabel metal2 432814 1530 432814 1530 0 ch_out[28]
rlabel metal1 446966 782 446966 782 0 ch_out[29]
rlabel metal1 31205 782 31205 782 0 ch_out[2]
rlabel metal2 28382 8653 28382 8653 0 ch_out[30]
rlabel metal2 481022 1530 481022 1530 0 ch_out[31]
rlabel metal2 496478 1156 496478 1156 0 ch_out[32]
rlabel metal2 29210 8585 29210 8585 0 ch_out[33]
rlabel metal1 523855 782 523855 782 0 ch_out[34]
rlabel metal2 542846 1156 542846 1156 0 ch_out[35]
rlabel metal1 81650 6732 81650 6732 0 ch_out[36]
rlabel metal2 573758 1156 573758 1156 0 ch_out[37]
rlabel metal2 589214 1530 589214 1530 0 ch_out[38]
rlabel metal2 30866 7905 30866 7905 0 ch_out[39]
rlabel metal1 20973 9214 20973 9214 0 ch_out[3]
rlabel metal2 618286 1156 618286 1156 0 ch_out[40]
rlabel metal1 630437 782 630437 782 0 ch_out[41]
rlabel metal1 61685 782 61685 782 0 ch_out[4]
rlabel metal1 76919 782 76919 782 0 ch_out[5]
rlabel metal1 21781 8942 21781 8942 0 ch_out[6]
rlabel metal1 107405 782 107405 782 0 ch_out[7]
rlabel metal1 122597 782 122597 782 0 ch_out[8]
rlabel metal2 23322 6732 23322 6732 0 ch_out[9]
rlabel metal2 114494 3468 114494 3468 0 net1
rlabel metal1 246606 6664 246606 6664 0 net10
rlabel metal2 33534 7616 33534 7616 0 net100
rlabel metal2 203918 4148 203918 4148 0 net101
rlabel metal1 180780 5100 180780 5100 0 net102
rlabel metal2 264822 2754 264822 2754 0 net103
rlabel metal2 80638 6528 80638 6528 0 net104
rlabel metal1 249182 2414 249182 2414 0 net105
rlabel metal1 114954 5644 114954 5644 0 net106
rlabel metal2 127558 4624 127558 4624 0 net107
rlabel metal2 35558 6732 35558 6732 0 net108
rlabel metal2 112378 4692 112378 4692 0 net109
rlabel metal2 311926 5032 311926 5032 0 net11
rlabel metal2 82478 4828 82478 4828 0 net110
rlabel metal2 156630 2652 156630 2652 0 net111
rlabel metal1 406088 4454 406088 4454 0 net12
rlabel metal1 511336 2618 511336 2618 0 net13
rlabel metal2 123234 7446 123234 7446 0 net14
rlabel metal2 217902 6494 217902 6494 0 net15
rlabel metal1 402362 3468 402362 3468 0 net16
rlabel metal1 404524 3502 404524 3502 0 net17
rlabel metal2 403374 2652 403374 2652 0 net18
rlabel metal2 214958 6137 214958 6137 0 net19
rlabel metal1 603888 2618 603888 2618 0 net2
rlabel metal2 216522 5678 216522 5678 0 net20
rlabel metal2 309994 4284 309994 4284 0 net21
rlabel metal1 401350 3026 401350 3026 0 net22
rlabel metal2 214130 6018 214130 6018 0 net23
rlabel metal1 214820 6290 214820 6290 0 net24
rlabel metal2 308890 3468 308890 3468 0 net25
rlabel metal1 311581 2346 311581 2346 0 net26
rlabel metal2 212934 6052 212934 6052 0 net27
rlabel metal2 213762 4760 213762 4760 0 net28
rlabel metal2 326370 2856 326370 2856 0 net29
rlabel metal1 132480 6732 132480 6732 0 net3
rlabel metal2 211554 5950 211554 5950 0 net30
rlabel metal2 212750 4250 212750 4250 0 net31
rlabel metal2 211370 3468 211370 3468 0 net32
rlabel metal2 117990 5576 117990 5576 0 net33
rlabel metal2 233634 3026 233634 3026 0 net34
rlabel metal2 117438 5032 117438 5032 0 net35
rlabel metal2 115690 4080 115690 4080 0 net36
rlabel metal2 37766 5168 37766 5168 0 net37
rlabel metal2 635306 3298 635306 3298 0 net38
rlabel metal2 448822 4250 448822 4250 0 net39
rlabel metal2 220478 6732 220478 6732 0 net4
rlabel metal2 354614 5440 354614 5440 0 net40
rlabel metal1 353924 6290 353924 6290 0 net41
rlabel metal1 260084 7378 260084 7378 0 net42
rlabel metal2 72818 7752 72818 7752 0 net43
rlabel metal2 619850 3604 619850 3604 0 net44
rlabel metal1 526930 4080 526930 4080 0 net45
rlabel metal1 432400 5202 432400 5202 0 net46
rlabel metal2 245502 6596 245502 6596 0 net47
rlabel metal1 154422 6936 154422 6936 0 net48
rlabel metal2 57362 7820 57362 7820 0 net49
rlabel metal2 404570 4794 404570 4794 0 net5
rlabel metal2 497214 3876 497214 3876 0 net50
rlabel metal2 402546 4080 402546 4080 0 net51
rlabel metal1 401442 5202 401442 5202 0 net52
rlabel metal2 214590 6868 214590 6868 0 net53
rlabel metal1 213716 7378 213716 7378 0 net54
rlabel metal2 573482 3570 573482 3570 0 net55
rlabel metal2 387090 4352 387090 4352 0 net56
rlabel metal1 385986 5202 385986 5202 0 net57
rlabel metal1 215050 6120 215050 6120 0 net58
rlabel metal2 105846 7548 105846 7548 0 net59
rlabel metal2 407330 4896 407330 4896 0 net6
rlabel metal2 450846 3604 450846 3604 0 net60
rlabel metal1 387918 4080 387918 4080 0 net61
rlabel metal2 262614 5984 262614 5984 0 net62
rlabel metal2 261786 6494 261786 6494 0 net63
rlabel metal2 74934 7786 74934 7786 0 net64
rlabel metal2 527574 2754 527574 2754 0 net65
rlabel metal1 434194 4046 434194 4046 0 net66
rlabel metal2 247342 5848 247342 5848 0 net67
rlabel metal1 154284 7310 154284 7310 0 net68
rlabel metal2 59662 7140 59662 7140 0 net69
rlabel metal2 500526 4012 500526 4012 0 net7
rlabel metal2 404478 3876 404478 3876 0 net70
rlabel metal2 402638 3808 402638 3808 0 net71
rlabel metal1 262798 4692 262798 4692 0 net72
rlabel metal1 200790 6324 200790 6324 0 net73
rlabel metal2 389022 3468 389022 3468 0 net74
rlabel metal2 387826 4012 387826 4012 0 net75
rlabel metal1 205620 5712 205620 5712 0 net76
rlabel metal2 107870 7616 107870 7616 0 net77
rlabel metal2 450294 2788 450294 2788 0 net78
rlabel metal2 264362 4828 264362 4828 0 net79
rlabel metal2 499882 2856 499882 2856 0 net8
rlabel metal2 262982 6256 262982 6256 0 net80
rlabel metal2 76958 7650 76958 7650 0 net81
rlabel metal1 404662 3400 404662 3400 0 net82
rlabel metal2 248998 4862 248998 4862 0 net83
rlabel metal2 167210 6171 167210 6171 0 net84
rlabel metal1 61778 7276 61778 7276 0 net85
rlabel metal1 403443 2414 403443 2414 0 net86
rlabel metal1 310960 4590 310960 4590 0 net87
rlabel metal2 154330 6256 154330 6256 0 net88
rlabel metal2 388010 3366 388010 3366 0 net89
rlabel metal1 209760 6392 209760 6392 0 net9
rlabel metal1 211186 4488 211186 4488 0 net90
rlabel metal1 117254 6664 117254 6664 0 net91
rlabel metal2 265282 3808 265282 3808 0 net92
rlabel metal1 261073 4794 261073 4794 0 net93
rlabel metal2 79350 6613 79350 6613 0 net94
rlabel metal2 249734 3706 249734 3706 0 net95
rlabel metal2 156998 5678 156998 5678 0 net96
rlabel metal2 155802 6528 155802 6528 0 net97
rlabel metal1 307648 2958 307648 2958 0 net98
rlabel metal1 209760 5032 209760 5032 0 net99
<< properties >>
string FIXED_BBOX 0 0 650000 10000
<< end >>
